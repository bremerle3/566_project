
module system_top ( HCLK_top, HRESETn_top, SYSRESETREQ_top_out, LOCKUP_top_out, 
        TXEV_top_out );
  input HCLK_top, HRESETn_top;
  output SYSRESETREQ_top_out, LOCKUP_top_out, TXEV_top_out;
  wire   HREADY_top, PID_hmastlock_top, \PID_htrans_top[1] , PID_hwrite_top,
         RAM_hready_resp_top, \RAM_hresp_top[0] , RAM_hsel_top,
         i_ssi_ssi_clk_top, i_ssi_ssi_rst_n_top, i_ssi_sclk_out_top,
         i_ssi_ss_0_n_top, i_ssi_ssi_mst_intr_n_top, i_ssi_ssi_oe_n_top,
         i_ssi_ssi_rxf_intr_n_top, i_ssi_ssi_rxo_intr_n_top,
         i_ssi_ssi_rxu_intr_n_top, i_ssi_ssi_sleep_top,
         i_ssi_ssi_txe_intr_n_top, i_ssi_ssi_intr_n_top, i_ssi_txd_top,
         \interconnect_ip_inst/n5991 , \interconnect_ip_inst/n6491 ,
         \interconnect_ip_inst/i_apb_hready_resp ,
         \interconnect_ip_inst/n4829 , \interconnect_ip_inst/i_ssi_fsm_sleep ,
         \interconnect_ip_inst/i_ssi_U_mstfsm_c_state[3] ,
         \interconnect_ip_inst/n4860 , \interconnect_ip_inst/n4861 ,
         \interconnect_ip_inst/n4862 , \interconnect_ip_inst/n4863 ,
         \interconnect_ip_inst/n4864 ,
         \interconnect_ip_inst/i_ahb_hresp_none_0_ ,
         \interconnect_ip_inst/i_ahb_U_dfltslv_N4 ,
         \interconnect_ip_inst/i_ahb_U_dfltslv_current_state ,
         \interconnect_ip_inst/n10765 , \interconnect_ip_inst/n11572 ,
         \CORTEXM0DS_INST/cm0_primask[0] , \CORTEXM0DS_INST/cm0_control[1] ,
         \CORTEXM0DS_INST/cm0_xpsr[24] , \CORTEXM0DS_INST/u_logic/N4816 ,
         \CORTEXM0DS_INST/u_logic/N4767 , \CORTEXM0DS_INST/u_logic/N4751 ,
         \CORTEXM0DS_INST/u_logic/N4674 , \CORTEXM0DS_INST/u_logic/N4518 ,
         \CORTEXM0DS_INST/u_logic/N4439 , \CORTEXM0DS_INST/u_logic/N4422 ,
         \CORTEXM0DS_INST/u_logic/N4421 , \CORTEXM0DS_INST/u_logic/N4396 ,
         \CORTEXM0DS_INST/u_logic/N4359 , \CORTEXM0DS_INST/u_logic/N4282 ,
         \CORTEXM0DS_INST/u_logic/N4227 , \CORTEXM0DS_INST/u_logic/N4170 ,
         \CORTEXM0DS_INST/u_logic/N4116 , \CORTEXM0DS_INST/u_logic/N4005 ,
         \CORTEXM0DS_INST/u_logic/N3967 , \CORTEXM0DS_INST/u_logic/N3966 ,
         \CORTEXM0DS_INST/u_logic/N3946 , \CORTEXM0DS_INST/u_logic/N3783 ,
         \CORTEXM0DS_INST/u_logic/N2678 , \CORTEXM0DS_INST/u_logic/N1447 ,
         \CORTEXM0DS_INST/u_logic/N586 , \CORTEXM0DS_INST/u_logic/E562z4 ,
         \CORTEXM0DS_INST/u_logic/Q462z4 , \CORTEXM0DS_INST/u_logic/A362z4 ,
         \CORTEXM0DS_INST/u_logic/Oq42z4 , \CORTEXM0DS_INST/u_logic/Xmywx4 ,
         \CORTEXM0DS_INST/u_logic/Ldhvx4 , \CORTEXM0DS_INST/u_logic/Sdhvx4 ,
         \CORTEXM0DS_INST/u_logic/Zdhvx4 , \CORTEXM0DS_INST/u_logic/Gehvx4 ,
         \CORTEXM0DS_INST/u_logic/Nehvx4 , \CORTEXM0DS_INST/u_logic/Uehvx4 ,
         \CORTEXM0DS_INST/u_logic/Bfhvx4 , \CORTEXM0DS_INST/u_logic/Ifhvx4 ,
         \CORTEXM0DS_INST/u_logic/Pfhvx4 , \CORTEXM0DS_INST/u_logic/Wfhvx4 ,
         \CORTEXM0DS_INST/u_logic/Dghvx4 , \CORTEXM0DS_INST/u_logic/Rghvx4 ,
         \CORTEXM0DS_INST/u_logic/Mhhvx4 , \CORTEXM0DS_INST/u_logic/Thhvx4 ,
         \CORTEXM0DS_INST/u_logic/Aihvx4 , \CORTEXM0DS_INST/u_logic/Hihvx4 ,
         \CORTEXM0DS_INST/u_logic/Oihvx4 , \CORTEXM0DS_INST/u_logic/Vihvx4 ,
         \CORTEXM0DS_INST/u_logic/Cjhvx4 , \CORTEXM0DS_INST/u_logic/Jjhvx4 ,
         \CORTEXM0DS_INST/u_logic/Qjhvx4 , \CORTEXM0DS_INST/u_logic/Xjhvx4 ,
         \CORTEXM0DS_INST/u_logic/Ekhvx4 , \CORTEXM0DS_INST/u_logic/Lkhvx4 ,
         \CORTEXM0DS_INST/u_logic/Skhvx4 , \CORTEXM0DS_INST/u_logic/Zkhvx4 ,
         \CORTEXM0DS_INST/u_logic/Glhvx4 , \CORTEXM0DS_INST/u_logic/Nlhvx4 ,
         \CORTEXM0DS_INST/u_logic/Ulhvx4 , \CORTEXM0DS_INST/u_logic/Bmhvx4 ,
         \CORTEXM0DS_INST/u_logic/Imhvx4 , \CORTEXM0DS_INST/u_logic/Lrhvx4 ,
         \CORTEXM0DS_INST/u_logic/Ithvx4 , \CORTEXM0DS_INST/u_logic/Pthvx4 ,
         \CORTEXM0DS_INST/u_logic/Wthvx4 , \CORTEXM0DS_INST/u_logic/Duhvx4 ,
         \CORTEXM0DS_INST/u_logic/Kuhvx4 , \CORTEXM0DS_INST/u_logic/Ruhvx4 ,
         \CORTEXM0DS_INST/u_logic/Yuhvx4 , \CORTEXM0DS_INST/u_logic/Fvhvx4 ,
         \CORTEXM0DS_INST/u_logic/Mvhvx4 , \CORTEXM0DS_INST/u_logic/Tvhvx4 ,
         \CORTEXM0DS_INST/u_logic/Awhvx4 , \CORTEXM0DS_INST/u_logic/Hwhvx4 ,
         \CORTEXM0DS_INST/u_logic/Owhvx4 , \CORTEXM0DS_INST/u_logic/Vwhvx4 ,
         \CORTEXM0DS_INST/u_logic/Cxhvx4 , \CORTEXM0DS_INST/u_logic/Jxhvx4 ,
         \CORTEXM0DS_INST/u_logic/Qxhvx4 , \CORTEXM0DS_INST/u_logic/Xxhvx4 ,
         \CORTEXM0DS_INST/u_logic/Eyhvx4 , \CORTEXM0DS_INST/u_logic/Lyhvx4 ,
         \CORTEXM0DS_INST/u_logic/Bq5wx4 , \CORTEXM0DS_INST/u_logic/Owgvx4 ,
         \CORTEXM0DS_INST/u_logic/T2ivx4 , \CORTEXM0DS_INST/u_logic/F2ivx4 ,
         \CORTEXM0DS_INST/u_logic/Y1ivx4 , \CORTEXM0DS_INST/u_logic/M2ivx4 ,
         \CORTEXM0DS_INST/u_logic/K1ivx4 , \CORTEXM0DS_INST/u_logic/D1ivx4 ,
         \CORTEXM0DS_INST/u_logic/R1ivx4 , \CORTEXM0DS_INST/u_logic/P0ivx4 ,
         \CORTEXM0DS_INST/u_logic/I0ivx4 , \CORTEXM0DS_INST/u_logic/W0ivx4 ,
         \CORTEXM0DS_INST/u_logic/B0ivx4 , \CORTEXM0DS_INST/u_logic/Uzhvx4 ,
         \CORTEXM0DS_INST/u_logic/Gzhvx4 , \CORTEXM0DS_INST/u_logic/Zyhvx4 ,
         \CORTEXM0DS_INST/u_logic/Nzhvx4 , \CORTEXM0DS_INST/u_logic/Syhvx4 ,
         \CORTEXM0DS_INST/u_logic/O24wx4 , \CORTEXM0DS_INST/u_logic/Sx3wx4 ,
         \CORTEXM0DS_INST/u_logic/H3ivx4 , \CORTEXM0DS_INST/u_logic/V3ivx4 ,
         \CORTEXM0DS_INST/u_logic/C4ivx4 , \CORTEXM0DS_INST/u_logic/J4ivx4 ,
         \CORTEXM0DS_INST/u_logic/Q4ivx4 , \CORTEXM0DS_INST/u_logic/X4ivx4 ,
         \CORTEXM0DS_INST/u_logic/E5ivx4 , \CORTEXM0DS_INST/u_logic/L5ivx4 ,
         \CORTEXM0DS_INST/u_logic/S5ivx4 , \CORTEXM0DS_INST/u_logic/Z5ivx4 ,
         \CORTEXM0DS_INST/u_logic/G6ivx4 , \CORTEXM0DS_INST/u_logic/N6ivx4 ,
         \CORTEXM0DS_INST/u_logic/U6ivx4 , \CORTEXM0DS_INST/u_logic/B7ivx4 ,
         \CORTEXM0DS_INST/u_logic/I7ivx4 , \CORTEXM0DS_INST/u_logic/P7ivx4 ,
         \CORTEXM0DS_INST/u_logic/W7ivx4 , \CORTEXM0DS_INST/u_logic/D8ivx4 ,
         \CORTEXM0DS_INST/u_logic/Y92wx4 , \CORTEXM0DS_INST/u_logic/R8ivx4 ,
         \CORTEXM0DS_INST/u_logic/Y8ivx4 , \CORTEXM0DS_INST/u_logic/F9ivx4 ,
         \CORTEXM0DS_INST/u_logic/M9ivx4 , \CORTEXM0DS_INST/u_logic/T9ivx4 ,
         \CORTEXM0DS_INST/u_logic/Aaivx4 , \CORTEXM0DS_INST/u_logic/Haivx4 ,
         \CORTEXM0DS_INST/u_logic/Oaivx4 , \CORTEXM0DS_INST/u_logic/Vaivx4 ,
         \CORTEXM0DS_INST/u_logic/Cbivx4 , \CORTEXM0DS_INST/u_logic/Jbivx4 ,
         \CORTEXM0DS_INST/u_logic/Qbivx4 , \CORTEXM0DS_INST/u_logic/Xbivx4 ,
         \CORTEXM0DS_INST/u_logic/Ecivx4 , \CORTEXM0DS_INST/u_logic/Lcivx4 ,
         \CORTEXM0DS_INST/u_logic/Scivx4 , \CORTEXM0DS_INST/u_logic/Gdivx4 ,
         \CORTEXM0DS_INST/u_logic/Ndivx4 , \CORTEXM0DS_INST/u_logic/Udivx4 ,
         \CORTEXM0DS_INST/u_logic/Beivx4 , \CORTEXM0DS_INST/u_logic/Ieivx4 ,
         \CORTEXM0DS_INST/u_logic/Peivx4 , \CORTEXM0DS_INST/u_logic/Weivx4 ,
         \CORTEXM0DS_INST/u_logic/Dfivx4 , \CORTEXM0DS_INST/u_logic/Kfivx4 ,
         \CORTEXM0DS_INST/u_logic/Rfivx4 , \CORTEXM0DS_INST/u_logic/Yfivx4 ,
         \CORTEXM0DS_INST/u_logic/Fgivx4 , \CORTEXM0DS_INST/u_logic/Mgivx4 ,
         \CORTEXM0DS_INST/u_logic/Tgivx4 , \CORTEXM0DS_INST/u_logic/Ahivx4 ,
         \CORTEXM0DS_INST/u_logic/Hhivx4 , \CORTEXM0DS_INST/u_logic/Vhivx4 ,
         \CORTEXM0DS_INST/u_logic/Ciivx4 , \CORTEXM0DS_INST/u_logic/Jiivx4 ,
         \CORTEXM0DS_INST/u_logic/Qiivx4 , \CORTEXM0DS_INST/u_logic/Xiivx4 ,
         \CORTEXM0DS_INST/u_logic/Ejivx4 , \CORTEXM0DS_INST/u_logic/Ljivx4 ,
         \CORTEXM0DS_INST/u_logic/Sjivx4 , \CORTEXM0DS_INST/u_logic/Zjivx4 ,
         \CORTEXM0DS_INST/u_logic/Gkivx4 , \CORTEXM0DS_INST/u_logic/Nkivx4 ,
         \CORTEXM0DS_INST/u_logic/Ukivx4 , \CORTEXM0DS_INST/u_logic/Blivx4 ,
         \CORTEXM0DS_INST/u_logic/Ilivx4 , \CORTEXM0DS_INST/u_logic/Plivx4 ,
         \CORTEXM0DS_INST/u_logic/Wlivx4 , \CORTEXM0DS_INST/u_logic/Kmivx4 ,
         \CORTEXM0DS_INST/u_logic/Rmivx4 , \CORTEXM0DS_INST/u_logic/Ymivx4 ,
         \CORTEXM0DS_INST/u_logic/Fnivx4 , \CORTEXM0DS_INST/u_logic/Mnivx4 ,
         \CORTEXM0DS_INST/u_logic/Tnivx4 , \CORTEXM0DS_INST/u_logic/Aoivx4 ,
         \CORTEXM0DS_INST/u_logic/Hoivx4 , \CORTEXM0DS_INST/u_logic/Ooivx4 ,
         \CORTEXM0DS_INST/u_logic/Voivx4 , \CORTEXM0DS_INST/u_logic/Cpivx4 ,
         \CORTEXM0DS_INST/u_logic/Jpivx4 , \CORTEXM0DS_INST/u_logic/Qpivx4 ,
         \CORTEXM0DS_INST/u_logic/Xpivx4 , \CORTEXM0DS_INST/u_logic/Eqivx4 ,
         \CORTEXM0DS_INST/u_logic/Lqivx4 , \CORTEXM0DS_INST/u_logic/Sqivx4 ,
         \CORTEXM0DS_INST/u_logic/Zqivx4 , \CORTEXM0DS_INST/u_logic/Grivx4 ,
         \CORTEXM0DS_INST/u_logic/Nrivx4 , \CORTEXM0DS_INST/u_logic/Urivx4 ,
         \CORTEXM0DS_INST/u_logic/Bsivx4 , \CORTEXM0DS_INST/u_logic/Isivx4 ,
         \CORTEXM0DS_INST/u_logic/Psivx4 , \CORTEXM0DS_INST/u_logic/Wsivx4 ,
         \CORTEXM0DS_INST/u_logic/Dtivx4 , \CORTEXM0DS_INST/u_logic/Ktivx4 ,
         \CORTEXM0DS_INST/u_logic/Rtivx4 , \CORTEXM0DS_INST/u_logic/Ytivx4 ,
         \CORTEXM0DS_INST/u_logic/Fuivx4 , \CORTEXM0DS_INST/u_logic/Muivx4 ,
         \CORTEXM0DS_INST/u_logic/Tuivx4 , \CORTEXM0DS_INST/u_logic/Avivx4 ,
         \CORTEXM0DS_INST/u_logic/Ovivx4 , \CORTEXM0DS_INST/u_logic/Vvivx4 ,
         \CORTEXM0DS_INST/u_logic/Cwivx4 , \CORTEXM0DS_INST/u_logic/Jwivx4 ,
         \CORTEXM0DS_INST/u_logic/Qwivx4 , \CORTEXM0DS_INST/u_logic/Xwivx4 ,
         \CORTEXM0DS_INST/u_logic/Exivx4 , \CORTEXM0DS_INST/u_logic/Lxivx4 ,
         \CORTEXM0DS_INST/u_logic/Sxivx4 , \CORTEXM0DS_INST/u_logic/Zxivx4 ,
         \CORTEXM0DS_INST/u_logic/Gyivx4 , \CORTEXM0DS_INST/u_logic/Nyivx4 ,
         \CORTEXM0DS_INST/u_logic/Uyivx4 , \CORTEXM0DS_INST/u_logic/Bzivx4 ,
         \CORTEXM0DS_INST/u_logic/Izivx4 , \CORTEXM0DS_INST/u_logic/Pzivx4 ,
         \CORTEXM0DS_INST/u_logic/D0jvx4 , \CORTEXM0DS_INST/u_logic/K0jvx4 ,
         \CORTEXM0DS_INST/u_logic/R0jvx4 , \CORTEXM0DS_INST/u_logic/Y0jvx4 ,
         \CORTEXM0DS_INST/u_logic/F1jvx4 , \CORTEXM0DS_INST/u_logic/M1jvx4 ,
         \CORTEXM0DS_INST/u_logic/T1jvx4 , \CORTEXM0DS_INST/u_logic/A2jvx4 ,
         \CORTEXM0DS_INST/u_logic/H2jvx4 , \CORTEXM0DS_INST/u_logic/O2jvx4 ,
         \CORTEXM0DS_INST/u_logic/V2jvx4 , \CORTEXM0DS_INST/u_logic/C3jvx4 ,
         \CORTEXM0DS_INST/u_logic/J3jvx4 , \CORTEXM0DS_INST/u_logic/Q3jvx4 ,
         \CORTEXM0DS_INST/u_logic/X3jvx4 , \CORTEXM0DS_INST/u_logic/E4jvx4 ,
         \CORTEXM0DS_INST/u_logic/S4jvx4 , \CORTEXM0DS_INST/u_logic/Z4jvx4 ,
         \CORTEXM0DS_INST/u_logic/G5jvx4 , \CORTEXM0DS_INST/u_logic/N5jvx4 ,
         \CORTEXM0DS_INST/u_logic/U5jvx4 , \CORTEXM0DS_INST/u_logic/B6jvx4 ,
         \CORTEXM0DS_INST/u_logic/I6jvx4 , \CORTEXM0DS_INST/u_logic/P6jvx4 ,
         \CORTEXM0DS_INST/u_logic/W6jvx4 , \CORTEXM0DS_INST/u_logic/D7jvx4 ,
         \CORTEXM0DS_INST/u_logic/K7jvx4 , \CORTEXM0DS_INST/u_logic/R7jvx4 ,
         \CORTEXM0DS_INST/u_logic/Y7jvx4 , \CORTEXM0DS_INST/u_logic/F8jvx4 ,
         \CORTEXM0DS_INST/u_logic/M8jvx4 , \CORTEXM0DS_INST/u_logic/T8jvx4 ,
         \CORTEXM0DS_INST/u_logic/H9jvx4 , \CORTEXM0DS_INST/u_logic/O9jvx4 ,
         \CORTEXM0DS_INST/u_logic/V9jvx4 , \CORTEXM0DS_INST/u_logic/Cajvx4 ,
         \CORTEXM0DS_INST/u_logic/Jajvx4 , \CORTEXM0DS_INST/u_logic/Qajvx4 ,
         \CORTEXM0DS_INST/u_logic/Xajvx4 , \CORTEXM0DS_INST/u_logic/Ebjvx4 ,
         \CORTEXM0DS_INST/u_logic/Lbjvx4 , \CORTEXM0DS_INST/u_logic/Sbjvx4 ,
         \CORTEXM0DS_INST/u_logic/Zbjvx4 , \CORTEXM0DS_INST/u_logic/Gcjvx4 ,
         \CORTEXM0DS_INST/u_logic/Ncjvx4 , \CORTEXM0DS_INST/u_logic/Ucjvx4 ,
         \CORTEXM0DS_INST/u_logic/Bdjvx4 , \CORTEXM0DS_INST/u_logic/Idjvx4 ,
         \CORTEXM0DS_INST/u_logic/Wdjvx4 , \CORTEXM0DS_INST/u_logic/Dejvx4 ,
         \CORTEXM0DS_INST/u_logic/Kejvx4 , \CORTEXM0DS_INST/u_logic/Rejvx4 ,
         \CORTEXM0DS_INST/u_logic/Yejvx4 , \CORTEXM0DS_INST/u_logic/Ffjvx4 ,
         \CORTEXM0DS_INST/u_logic/Mfjvx4 , \CORTEXM0DS_INST/u_logic/Tfjvx4 ,
         \CORTEXM0DS_INST/u_logic/Agjvx4 , \CORTEXM0DS_INST/u_logic/Hgjvx4 ,
         \CORTEXM0DS_INST/u_logic/Ogjvx4 , \CORTEXM0DS_INST/u_logic/Vgjvx4 ,
         \CORTEXM0DS_INST/u_logic/Chjvx4 , \CORTEXM0DS_INST/u_logic/Jhjvx4 ,
         \CORTEXM0DS_INST/u_logic/Qhjvx4 , \CORTEXM0DS_INST/u_logic/Xhjvx4 ,
         \CORTEXM0DS_INST/u_logic/Lijvx4 , \CORTEXM0DS_INST/u_logic/Sijvx4 ,
         \CORTEXM0DS_INST/u_logic/Zijvx4 , \CORTEXM0DS_INST/u_logic/Gjjvx4 ,
         \CORTEXM0DS_INST/u_logic/Njjvx4 , \CORTEXM0DS_INST/u_logic/Ujjvx4 ,
         \CORTEXM0DS_INST/u_logic/Bkjvx4 , \CORTEXM0DS_INST/u_logic/Ikjvx4 ,
         \CORTEXM0DS_INST/u_logic/Pkjvx4 , \CORTEXM0DS_INST/u_logic/Wkjvx4 ,
         \CORTEXM0DS_INST/u_logic/Dljvx4 , \CORTEXM0DS_INST/u_logic/Kljvx4 ,
         \CORTEXM0DS_INST/u_logic/Rljvx4 , \CORTEXM0DS_INST/u_logic/Yljvx4 ,
         \CORTEXM0DS_INST/u_logic/Fmjvx4 , \CORTEXM0DS_INST/u_logic/Mmjvx4 ,
         \CORTEXM0DS_INST/u_logic/Bv0wx4 , \CORTEXM0DS_INST/u_logic/Anjvx4 ,
         \CORTEXM0DS_INST/u_logic/Hnjvx4 , \CORTEXM0DS_INST/u_logic/Onjvx4 ,
         \CORTEXM0DS_INST/u_logic/Vnjvx4 , \CORTEXM0DS_INST/u_logic/Cojvx4 ,
         \CORTEXM0DS_INST/u_logic/Jojvx4 , \CORTEXM0DS_INST/u_logic/Qojvx4 ,
         \CORTEXM0DS_INST/u_logic/Xojvx4 , \CORTEXM0DS_INST/u_logic/Epjvx4 ,
         \CORTEXM0DS_INST/u_logic/Lpjvx4 , \CORTEXM0DS_INST/u_logic/Spjvx4 ,
         \CORTEXM0DS_INST/u_logic/Zpjvx4 , \CORTEXM0DS_INST/u_logic/Gqjvx4 ,
         \CORTEXM0DS_INST/u_logic/Nqjvx4 , \CORTEXM0DS_INST/u_logic/Uqjvx4 ,
         \CORTEXM0DS_INST/u_logic/Brjvx4 , \CORTEXM0DS_INST/u_logic/Fq0wx4 ,
         \CORTEXM0DS_INST/u_logic/Prjvx4 , \CORTEXM0DS_INST/u_logic/Wrjvx4 ,
         \CORTEXM0DS_INST/u_logic/Dsjvx4 , \CORTEXM0DS_INST/u_logic/Ksjvx4 ,
         \CORTEXM0DS_INST/u_logic/Rsjvx4 , \CORTEXM0DS_INST/u_logic/Ysjvx4 ,
         \CORTEXM0DS_INST/u_logic/Ftjvx4 , \CORTEXM0DS_INST/u_logic/Mtjvx4 ,
         \CORTEXM0DS_INST/u_logic/Ttjvx4 , \CORTEXM0DS_INST/u_logic/Aujvx4 ,
         \CORTEXM0DS_INST/u_logic/Hujvx4 , \CORTEXM0DS_INST/u_logic/Oujvx4 ,
         \CORTEXM0DS_INST/u_logic/Vujvx4 , \CORTEXM0DS_INST/u_logic/Cvjvx4 ,
         \CORTEXM0DS_INST/u_logic/Jvjvx4 , \CORTEXM0DS_INST/u_logic/Qvjvx4 ,
         \CORTEXM0DS_INST/u_logic/Ql0wx4 , \CORTEXM0DS_INST/u_logic/Ewjvx4 ,
         \CORTEXM0DS_INST/u_logic/Lwjvx4 , \CORTEXM0DS_INST/u_logic/Swjvx4 ,
         \CORTEXM0DS_INST/u_logic/Zwjvx4 , \CORTEXM0DS_INST/u_logic/Gxjvx4 ,
         \CORTEXM0DS_INST/u_logic/Nxjvx4 , \CORTEXM0DS_INST/u_logic/Uxjvx4 ,
         \CORTEXM0DS_INST/u_logic/Byjvx4 , \CORTEXM0DS_INST/u_logic/Iyjvx4 ,
         \CORTEXM0DS_INST/u_logic/Pyjvx4 , \CORTEXM0DS_INST/u_logic/Wyjvx4 ,
         \CORTEXM0DS_INST/u_logic/Dzjvx4 , \CORTEXM0DS_INST/u_logic/Kzjvx4 ,
         \CORTEXM0DS_INST/u_logic/Rzjvx4 , \CORTEXM0DS_INST/u_logic/Yzjvx4 ,
         \CORTEXM0DS_INST/u_logic/F0kvx4 , \CORTEXM0DS_INST/u_logic/Ug0wx4 ,
         \CORTEXM0DS_INST/u_logic/T0kvx4 , \CORTEXM0DS_INST/u_logic/A1kvx4 ,
         \CORTEXM0DS_INST/u_logic/H1kvx4 , \CORTEXM0DS_INST/u_logic/O1kvx4 ,
         \CORTEXM0DS_INST/u_logic/V1kvx4 , \CORTEXM0DS_INST/u_logic/C2kvx4 ,
         \CORTEXM0DS_INST/u_logic/J2kvx4 , \CORTEXM0DS_INST/u_logic/Q2kvx4 ,
         \CORTEXM0DS_INST/u_logic/X2kvx4 , \CORTEXM0DS_INST/u_logic/E3kvx4 ,
         \CORTEXM0DS_INST/u_logic/L3kvx4 , \CORTEXM0DS_INST/u_logic/S3kvx4 ,
         \CORTEXM0DS_INST/u_logic/Z3kvx4 , \CORTEXM0DS_INST/u_logic/G4kvx4 ,
         \CORTEXM0DS_INST/u_logic/N4kvx4 , \CORTEXM0DS_INST/u_logic/U4kvx4 ,
         \CORTEXM0DS_INST/u_logic/Fc0wx4 , \CORTEXM0DS_INST/u_logic/I5kvx4 ,
         \CORTEXM0DS_INST/u_logic/P5kvx4 , \CORTEXM0DS_INST/u_logic/W5kvx4 ,
         \CORTEXM0DS_INST/u_logic/D6kvx4 , \CORTEXM0DS_INST/u_logic/K6kvx4 ,
         \CORTEXM0DS_INST/u_logic/R6kvx4 , \CORTEXM0DS_INST/u_logic/Y6kvx4 ,
         \CORTEXM0DS_INST/u_logic/F7kvx4 , \CORTEXM0DS_INST/u_logic/M7kvx4 ,
         \CORTEXM0DS_INST/u_logic/T7kvx4 , \CORTEXM0DS_INST/u_logic/A8kvx4 ,
         \CORTEXM0DS_INST/u_logic/H8kvx4 , \CORTEXM0DS_INST/u_logic/O8kvx4 ,
         \CORTEXM0DS_INST/u_logic/V8kvx4 , \CORTEXM0DS_INST/u_logic/C9kvx4 ,
         \CORTEXM0DS_INST/u_logic/J9kvx4 , \CORTEXM0DS_INST/u_logic/C70wx4 ,
         \CORTEXM0DS_INST/u_logic/X9kvx4 , \CORTEXM0DS_INST/u_logic/Eakvx4 ,
         \CORTEXM0DS_INST/u_logic/Lakvx4 , \CORTEXM0DS_INST/u_logic/Sakvx4 ,
         \CORTEXM0DS_INST/u_logic/Zakvx4 , \CORTEXM0DS_INST/u_logic/Gbkvx4 ,
         \CORTEXM0DS_INST/u_logic/Nbkvx4 , \CORTEXM0DS_INST/u_logic/Ubkvx4 ,
         \CORTEXM0DS_INST/u_logic/Bckvx4 , \CORTEXM0DS_INST/u_logic/Ickvx4 ,
         \CORTEXM0DS_INST/u_logic/Pckvx4 , \CORTEXM0DS_INST/u_logic/Wckvx4 ,
         \CORTEXM0DS_INST/u_logic/Ddkvx4 , \CORTEXM0DS_INST/u_logic/Kdkvx4 ,
         \CORTEXM0DS_INST/u_logic/Rdkvx4 , \CORTEXM0DS_INST/u_logic/Ydkvx4 ,
         \CORTEXM0DS_INST/u_logic/Fekvx4 , \CORTEXM0DS_INST/u_logic/Tekvx4 ,
         \CORTEXM0DS_INST/u_logic/Afkvx4 , \CORTEXM0DS_INST/u_logic/Hfkvx4 ,
         \CORTEXM0DS_INST/u_logic/Ofkvx4 , \CORTEXM0DS_INST/u_logic/Vfkvx4 ,
         \CORTEXM0DS_INST/u_logic/Cgkvx4 , \CORTEXM0DS_INST/u_logic/Jgkvx4 ,
         \CORTEXM0DS_INST/u_logic/Qgkvx4 , \CORTEXM0DS_INST/u_logic/Xgkvx4 ,
         \CORTEXM0DS_INST/u_logic/Ehkvx4 , \CORTEXM0DS_INST/u_logic/Lhkvx4 ,
         \CORTEXM0DS_INST/u_logic/Shkvx4 , \CORTEXM0DS_INST/u_logic/Zhkvx4 ,
         \CORTEXM0DS_INST/u_logic/Gikvx4 , \CORTEXM0DS_INST/u_logic/Nikvx4 ,
         \CORTEXM0DS_INST/u_logic/Uikvx4 , \CORTEXM0DS_INST/u_logic/Ijkvx4 ,
         \CORTEXM0DS_INST/u_logic/Pjkvx4 , \CORTEXM0DS_INST/u_logic/Wjkvx4 ,
         \CORTEXM0DS_INST/u_logic/Dkkvx4 , \CORTEXM0DS_INST/u_logic/Kkkvx4 ,
         \CORTEXM0DS_INST/u_logic/Rkkvx4 , \CORTEXM0DS_INST/u_logic/Ykkvx4 ,
         \CORTEXM0DS_INST/u_logic/Flkvx4 , \CORTEXM0DS_INST/u_logic/Mlkvx4 ,
         \CORTEXM0DS_INST/u_logic/Tlkvx4 , \CORTEXM0DS_INST/u_logic/Amkvx4 ,
         \CORTEXM0DS_INST/u_logic/Hmkvx4 , \CORTEXM0DS_INST/u_logic/Omkvx4 ,
         \CORTEXM0DS_INST/u_logic/Vmkvx4 , \CORTEXM0DS_INST/u_logic/Cnkvx4 ,
         \CORTEXM0DS_INST/u_logic/Jnkvx4 , \CORTEXM0DS_INST/u_logic/Rxzvx4 ,
         \CORTEXM0DS_INST/u_logic/Xnkvx4 , \CORTEXM0DS_INST/u_logic/Eokvx4 ,
         \CORTEXM0DS_INST/u_logic/Lokvx4 , \CORTEXM0DS_INST/u_logic/Sokvx4 ,
         \CORTEXM0DS_INST/u_logic/Zokvx4 , \CORTEXM0DS_INST/u_logic/Gpkvx4 ,
         \CORTEXM0DS_INST/u_logic/Npkvx4 , \CORTEXM0DS_INST/u_logic/Upkvx4 ,
         \CORTEXM0DS_INST/u_logic/Bqkvx4 , \CORTEXM0DS_INST/u_logic/Iqkvx4 ,
         \CORTEXM0DS_INST/u_logic/Pqkvx4 , \CORTEXM0DS_INST/u_logic/Wqkvx4 ,
         \CORTEXM0DS_INST/u_logic/Drkvx4 , \CORTEXM0DS_INST/u_logic/Krkvx4 ,
         \CORTEXM0DS_INST/u_logic/Rrkvx4 , \CORTEXM0DS_INST/u_logic/Yrkvx4 ,
         \CORTEXM0DS_INST/u_logic/Hszvx4 , \CORTEXM0DS_INST/u_logic/Mskvx4 ,
         \CORTEXM0DS_INST/u_logic/Tskvx4 , \CORTEXM0DS_INST/u_logic/Atkvx4 ,
         \CORTEXM0DS_INST/u_logic/Htkvx4 , \CORTEXM0DS_INST/u_logic/Otkvx4 ,
         \CORTEXM0DS_INST/u_logic/Vtkvx4 , \CORTEXM0DS_INST/u_logic/Cukvx4 ,
         \CORTEXM0DS_INST/u_logic/Jukvx4 , \CORTEXM0DS_INST/u_logic/Qukvx4 ,
         \CORTEXM0DS_INST/u_logic/Xukvx4 , \CORTEXM0DS_INST/u_logic/Evkvx4 ,
         \CORTEXM0DS_INST/u_logic/Lvkvx4 , \CORTEXM0DS_INST/u_logic/Svkvx4 ,
         \CORTEXM0DS_INST/u_logic/Zvkvx4 , \CORTEXM0DS_INST/u_logic/Gwkvx4 ,
         \CORTEXM0DS_INST/u_logic/Nwkvx4 , \CORTEXM0DS_INST/u_logic/Uwkvx4 ,
         \CORTEXM0DS_INST/u_logic/Bxkvx4 , \CORTEXM0DS_INST/u_logic/Ixkvx4 ,
         \CORTEXM0DS_INST/u_logic/Pxkvx4 , \CORTEXM0DS_INST/u_logic/Wxkvx4 ,
         \CORTEXM0DS_INST/u_logic/Dykvx4 , \CORTEXM0DS_INST/u_logic/Kykvx4 ,
         \CORTEXM0DS_INST/u_logic/Rykvx4 , \CORTEXM0DS_INST/u_logic/Yykvx4 ,
         \CORTEXM0DS_INST/u_logic/Fzkvx4 , \CORTEXM0DS_INST/u_logic/Mzkvx4 ,
         \CORTEXM0DS_INST/u_logic/Tzkvx4 , \CORTEXM0DS_INST/u_logic/A0lvx4 ,
         \CORTEXM0DS_INST/u_logic/H0lvx4 , \CORTEXM0DS_INST/u_logic/O0lvx4 ,
         \CORTEXM0DS_INST/u_logic/V0lvx4 , \CORTEXM0DS_INST/u_logic/J1lvx4 ,
         \CORTEXM0DS_INST/u_logic/Q1lvx4 , \CORTEXM0DS_INST/u_logic/X1lvx4 ,
         \CORTEXM0DS_INST/u_logic/E2lvx4 , \CORTEXM0DS_INST/u_logic/L2lvx4 ,
         \CORTEXM0DS_INST/u_logic/S2lvx4 , \CORTEXM0DS_INST/u_logic/Z2lvx4 ,
         \CORTEXM0DS_INST/u_logic/G3lvx4 , \CORTEXM0DS_INST/u_logic/N3lvx4 ,
         \CORTEXM0DS_INST/u_logic/U3lvx4 , \CORTEXM0DS_INST/u_logic/B4lvx4 ,
         \CORTEXM0DS_INST/u_logic/I4lvx4 , \CORTEXM0DS_INST/u_logic/P4lvx4 ,
         \CORTEXM0DS_INST/u_logic/W4lvx4 , \CORTEXM0DS_INST/u_logic/D5lvx4 ,
         \CORTEXM0DS_INST/u_logic/K5lvx4 , \CORTEXM0DS_INST/u_logic/Nhzvx4 ,
         \CORTEXM0DS_INST/u_logic/Y5lvx4 , \CORTEXM0DS_INST/u_logic/F6lvx4 ,
         \CORTEXM0DS_INST/u_logic/M6lvx4 , \CORTEXM0DS_INST/u_logic/T6lvx4 ,
         \CORTEXM0DS_INST/u_logic/A7lvx4 , \CORTEXM0DS_INST/u_logic/H7lvx4 ,
         \CORTEXM0DS_INST/u_logic/O7lvx4 , \CORTEXM0DS_INST/u_logic/V7lvx4 ,
         \CORTEXM0DS_INST/u_logic/C8lvx4 , \CORTEXM0DS_INST/u_logic/J8lvx4 ,
         \CORTEXM0DS_INST/u_logic/Q8lvx4 , \CORTEXM0DS_INST/u_logic/X8lvx4 ,
         \CORTEXM0DS_INST/u_logic/E9lvx4 , \CORTEXM0DS_INST/u_logic/L9lvx4 ,
         \CORTEXM0DS_INST/u_logic/S9lvx4 , \CORTEXM0DS_INST/u_logic/Z9lvx4 ,
         \CORTEXM0DS_INST/u_logic/Vezvx4 , \CORTEXM0DS_INST/u_logic/Nalvx4 ,
         \CORTEXM0DS_INST/u_logic/Ualvx4 , \CORTEXM0DS_INST/u_logic/Bblvx4 ,
         \CORTEXM0DS_INST/u_logic/Iblvx4 , \CORTEXM0DS_INST/u_logic/Pblvx4 ,
         \CORTEXM0DS_INST/u_logic/Wblvx4 , \CORTEXM0DS_INST/u_logic/Dclvx4 ,
         \CORTEXM0DS_INST/u_logic/Kclvx4 , \CORTEXM0DS_INST/u_logic/Rclvx4 ,
         \CORTEXM0DS_INST/u_logic/Yclvx4 , \CORTEXM0DS_INST/u_logic/Fdlvx4 ,
         \CORTEXM0DS_INST/u_logic/Mdlvx4 , \CORTEXM0DS_INST/u_logic/Tdlvx4 ,
         \CORTEXM0DS_INST/u_logic/Aelvx4 , \CORTEXM0DS_INST/u_logic/Helvx4 ,
         \CORTEXM0DS_INST/u_logic/Oelvx4 , \CORTEXM0DS_INST/u_logic/Cflvx4 ,
         \CORTEXM0DS_INST/u_logic/Jflvx4 , \CORTEXM0DS_INST/u_logic/Qflvx4 ,
         \CORTEXM0DS_INST/u_logic/Xflvx4 , \CORTEXM0DS_INST/u_logic/Eglvx4 ,
         \CORTEXM0DS_INST/u_logic/Lglvx4 , \CORTEXM0DS_INST/u_logic/Sglvx4 ,
         \CORTEXM0DS_INST/u_logic/Zglvx4 , \CORTEXM0DS_INST/u_logic/Ghlvx4 ,
         \CORTEXM0DS_INST/u_logic/Nhlvx4 , \CORTEXM0DS_INST/u_logic/Uhlvx4 ,
         \CORTEXM0DS_INST/u_logic/Bilvx4 , \CORTEXM0DS_INST/u_logic/Iilvx4 ,
         \CORTEXM0DS_INST/u_logic/Pilvx4 , \CORTEXM0DS_INST/u_logic/Wilvx4 ,
         \CORTEXM0DS_INST/u_logic/Djlvx4 , \CORTEXM0DS_INST/u_logic/Kjlvx4 ,
         \CORTEXM0DS_INST/u_logic/Rjlvx4 , \CORTEXM0DS_INST/u_logic/Yjlvx4 ,
         \CORTEXM0DS_INST/u_logic/Fklvx4 , \CORTEXM0DS_INST/u_logic/Mklvx4 ,
         \CORTEXM0DS_INST/u_logic/Tklvx4 , \CORTEXM0DS_INST/u_logic/Allvx4 ,
         \CORTEXM0DS_INST/u_logic/Hllvx4 , \CORTEXM0DS_INST/u_logic/Ollvx4 ,
         \CORTEXM0DS_INST/u_logic/Cmlvx4 , \CORTEXM0DS_INST/u_logic/Jmlvx4 ,
         \CORTEXM0DS_INST/u_logic/Qmlvx4 , \CORTEXM0DS_INST/u_logic/Xmlvx4 ,
         \CORTEXM0DS_INST/u_logic/Enlvx4 , \CORTEXM0DS_INST/u_logic/Lnlvx4 ,
         \CORTEXM0DS_INST/u_logic/Snlvx4 , \CORTEXM0DS_INST/u_logic/Znlvx4 ,
         \CORTEXM0DS_INST/u_logic/Golvx4 , \CORTEXM0DS_INST/u_logic/Nolvx4 ,
         \CORTEXM0DS_INST/u_logic/Uolvx4 , \CORTEXM0DS_INST/u_logic/Bplvx4 ,
         \CORTEXM0DS_INST/u_logic/Iplvx4 , \CORTEXM0DS_INST/u_logic/Pplvx4 ,
         \CORTEXM0DS_INST/u_logic/Wplvx4 , \CORTEXM0DS_INST/u_logic/Dqlvx4 ,
         \CORTEXM0DS_INST/u_logic/Kqlvx4 , \CORTEXM0DS_INST/u_logic/Rqlvx4 ,
         \CORTEXM0DS_INST/u_logic/Yqlvx4 , \CORTEXM0DS_INST/u_logic/Frlvx4 ,
         \CORTEXM0DS_INST/u_logic/Mrlvx4 , \CORTEXM0DS_INST/u_logic/Trlvx4 ,
         \CORTEXM0DS_INST/u_logic/Aslvx4 , \CORTEXM0DS_INST/u_logic/Hslvx4 ,
         \CORTEXM0DS_INST/u_logic/Oslvx4 , \CORTEXM0DS_INST/u_logic/Vslvx4 ,
         \CORTEXM0DS_INST/u_logic/Ctlvx4 , \CORTEXM0DS_INST/u_logic/Jtlvx4 ,
         \CORTEXM0DS_INST/u_logic/Qtlvx4 , \CORTEXM0DS_INST/u_logic/Xtlvx4 ,
         \CORTEXM0DS_INST/u_logic/Eulvx4 , \CORTEXM0DS_INST/u_logic/Lulvx4 ,
         \CORTEXM0DS_INST/u_logic/Sulvx4 , \CORTEXM0DS_INST/u_logic/Zulvx4 ,
         \CORTEXM0DS_INST/u_logic/Gvlvx4 , \CORTEXM0DS_INST/u_logic/Nvlvx4 ,
         \CORTEXM0DS_INST/u_logic/Uvlvx4 , \CORTEXM0DS_INST/u_logic/Bwlvx4 ,
         \CORTEXM0DS_INST/u_logic/Iwlvx4 , \CORTEXM0DS_INST/u_logic/Pwlvx4 ,
         \CORTEXM0DS_INST/u_logic/Wwlvx4 , \CORTEXM0DS_INST/u_logic/Dxlvx4 ,
         \CORTEXM0DS_INST/u_logic/Kxlvx4 , \CORTEXM0DS_INST/u_logic/Rxlvx4 ,
         \CORTEXM0DS_INST/u_logic/Yxlvx4 , \CORTEXM0DS_INST/u_logic/Fylvx4 ,
         \CORTEXM0DS_INST/u_logic/Mylvx4 , \CORTEXM0DS_INST/u_logic/Tylvx4 ,
         \CORTEXM0DS_INST/u_logic/Azlvx4 , \CORTEXM0DS_INST/u_logic/Hzlvx4 ,
         \CORTEXM0DS_INST/u_logic/Ozlvx4 , \CORTEXM0DS_INST/u_logic/Vzlvx4 ,
         \CORTEXM0DS_INST/u_logic/C0mvx4 , \CORTEXM0DS_INST/u_logic/J0mvx4 ,
         \CORTEXM0DS_INST/u_logic/Q0mvx4 , \CORTEXM0DS_INST/u_logic/X0mvx4 ,
         \CORTEXM0DS_INST/u_logic/E1mvx4 , \CORTEXM0DS_INST/u_logic/L1mvx4 ,
         \CORTEXM0DS_INST/u_logic/S1mvx4 , \CORTEXM0DS_INST/u_logic/Z1mvx4 ,
         \CORTEXM0DS_INST/u_logic/G2mvx4 , \CORTEXM0DS_INST/u_logic/N2mvx4 ,
         \CORTEXM0DS_INST/u_logic/U2mvx4 , \CORTEXM0DS_INST/u_logic/L8mvx4 ,
         \CORTEXM0DS_INST/u_logic/U9mvx4 , \CORTEXM0DS_INST/u_logic/Pamvx4 ,
         \CORTEXM0DS_INST/u_logic/Wamvx4 , \CORTEXM0DS_INST/u_logic/Jemvx4 ,
         \CORTEXM0DS_INST/u_logic/Qemvx4 , \CORTEXM0DS_INST/u_logic/Xemvx4 ,
         \CORTEXM0DS_INST/u_logic/Efmvx4 , \CORTEXM0DS_INST/u_logic/Lfmvx4 ,
         \CORTEXM0DS_INST/u_logic/Sfmvx4 , \CORTEXM0DS_INST/u_logic/Zfmvx4 ,
         \CORTEXM0DS_INST/u_logic/Ggmvx4 , \CORTEXM0DS_INST/u_logic/Ngmvx4 ,
         \CORTEXM0DS_INST/u_logic/Ugmvx4 , \CORTEXM0DS_INST/u_logic/Bhmvx4 ,
         \CORTEXM0DS_INST/u_logic/Ihmvx4 , \CORTEXM0DS_INST/u_logic/Phmvx4 ,
         \CORTEXM0DS_INST/u_logic/Whmvx4 , \CORTEXM0DS_INST/u_logic/Dimvx4 ,
         \CORTEXM0DS_INST/u_logic/Kimvx4 , \CORTEXM0DS_INST/u_logic/Rimvx4 ,
         \CORTEXM0DS_INST/u_logic/Yimvx4 , \CORTEXM0DS_INST/u_logic/Fjmvx4 ,
         \CORTEXM0DS_INST/u_logic/Mjmvx4 , \CORTEXM0DS_INST/u_logic/Tjmvx4 ,
         \CORTEXM0DS_INST/u_logic/Akmvx4 , \CORTEXM0DS_INST/u_logic/Hkmvx4 ,
         \CORTEXM0DS_INST/u_logic/Okmvx4 , \CORTEXM0DS_INST/u_logic/Vkmvx4 ,
         \CORTEXM0DS_INST/u_logic/Clmvx4 , \CORTEXM0DS_INST/u_logic/Jlmvx4 ,
         \CORTEXM0DS_INST/u_logic/Qlmvx4 , \CORTEXM0DS_INST/u_logic/Xlmvx4 ,
         \CORTEXM0DS_INST/u_logic/Emmvx4 , \CORTEXM0DS_INST/u_logic/Lmmvx4 ,
         \CORTEXM0DS_INST/u_logic/Smmvx4 , \CORTEXM0DS_INST/u_logic/F4nvx4 ,
         \CORTEXM0DS_INST/u_logic/G8nvx4 , \CORTEXM0DS_INST/u_logic/Acnvx4 ,
         \CORTEXM0DS_INST/u_logic/Ocnvx4 , \CORTEXM0DS_INST/u_logic/Jdnvx4 ,
         \CORTEXM0DS_INST/u_logic/Eenvx4 , \CORTEXM0DS_INST/u_logic/Lenvx4 ,
         \CORTEXM0DS_INST/u_logic/Senvx4 , \CORTEXM0DS_INST/u_logic/Zenvx4 ,
         \CORTEXM0DS_INST/u_logic/Gfnvx4 , \CORTEXM0DS_INST/u_logic/Ufnvx4 ,
         \CORTEXM0DS_INST/u_logic/Bgnvx4 , \CORTEXM0DS_INST/u_logic/Ignvx4 ,
         \CORTEXM0DS_INST/u_logic/S4qvx4 , \CORTEXM0DS_INST/u_logic/Wgnvx4 ,
         \CORTEXM0DS_INST/u_logic/Dhnvx4 , \CORTEXM0DS_INST/u_logic/V2qvx4 ,
         \CORTEXM0DS_INST/u_logic/Rhnvx4 , \CORTEXM0DS_INST/u_logic/Finvx4 ,
         \CORTEXM0DS_INST/u_logic/Minvx4 , \CORTEXM0DS_INST/u_logic/Tinvx4 ,
         \CORTEXM0DS_INST/u_logic/Ojnvx4 , \CORTEXM0DS_INST/u_logic/Y1pvx4 ,
         \CORTEXM0DS_INST/u_logic/Xxovx4 , \CORTEXM0DS_INST/u_logic/Jxovx4 ,
         \CORTEXM0DS_INST/u_logic/Owovx4 , \CORTEXM0DS_INST/u_logic/Fvovx4 ,
         \CORTEXM0DS_INST/u_logic/Yuovx4 , \CORTEXM0DS_INST/u_logic/Cqovx4 ,
         \CORTEXM0DS_INST/u_logic/Vpovx4 , \CORTEXM0DS_INST/u_logic/Rnovx4 ,
         \CORTEXM0DS_INST/u_logic/Ekovx4 , \CORTEXM0DS_INST/u_logic/Llnvx4 ,
         \CORTEXM0DS_INST/u_logic/Slnvx4 , \CORTEXM0DS_INST/u_logic/Z6ovx4 ,
         \CORTEXM0DS_INST/u_logic/Pxdvx4 , \CORTEXM0DS_INST/u_logic/H0gvx4 ,
         \CORTEXM0DS_INST/u_logic/W1evx4 , \CORTEXM0DS_INST/u_logic/Itdvx4 ,
         \CORTEXM0DS_INST/u_logic/Mqdvx4 , \CORTEXM0DS_INST/u_logic/Rddvx4 ,
         \CORTEXM0DS_INST/u_logic/Gcdvx4 , \CORTEXM0DS_INST/u_logic/Oy8vx4 ,
         \CORTEXM0DS_INST/u_logic/Fs8vx4 , \CORTEXM0DS_INST/u_logic/Vu8vx4 ,
         \CORTEXM0DS_INST/u_logic/Y3dvx4 , \CORTEXM0DS_INST/u_logic/S0hvx4 ,
         \CORTEXM0DS_INST/u_logic/F2hvx4 , \CORTEXM0DS_INST/u_logic/N6hvx4 ,
         \CORTEXM0DS_INST/u_logic/O2dvx4 , \CORTEXM0DS_INST/u_logic/E1dvx4 ,
         \CORTEXM0DS_INST/u_logic/Ukdvx4 , \CORTEXM0DS_INST/u_logic/C8dvx4 ,
         \CORTEXM0DS_INST/u_logic/S6dvx4 , \CORTEXM0DS_INST/u_logic/Nt8vx4 ,
         \CORTEXM0DS_INST/u_logic/Ks9vx4 , \CORTEXM0DS_INST/u_logic/Gr9vx4 ,
         \CORTEXM0DS_INST/u_logic/Cq9vx4 , \CORTEXM0DS_INST/u_logic/Uzcvx4 ,
         \CORTEXM0DS_INST/u_logic/Bx9vx4 , \CORTEXM0DS_INST/u_logic/Wv9vx4 ,
         \CORTEXM0DS_INST/u_logic/Cf9vx4 , \CORTEXM0DS_INST/u_logic/Ud9vx4 ,
         \CORTEXM0DS_INST/u_logic/Mc9vx4 , \CORTEXM0DS_INST/u_logic/Fb9vx4 ,
         \CORTEXM0DS_INST/u_logic/Y99vx4 , \CORTEXM0DS_INST/u_logic/R89vx4 ,
         \CORTEXM0DS_INST/u_logic/K79vx4 , \CORTEXM0DS_INST/u_logic/D69vx4 ,
         \CORTEXM0DS_INST/u_logic/W49vx4 , \CORTEXM0DS_INST/u_logic/P39vx4 ,
         \CORTEXM0DS_INST/u_logic/I29vx4 , \CORTEXM0DS_INST/u_logic/V8evx4 ,
         \CORTEXM0DS_INST/u_logic/G8fvx4 , \CORTEXM0DS_INST/u_logic/V6fvx4 ,
         \CORTEXM0DS_INST/u_logic/Z3fvx4 , \CORTEXM0DS_INST/u_logic/O2fvx4 ,
         \CORTEXM0DS_INST/u_logic/D1fvx4 , \CORTEXM0DS_INST/u_logic/Tzevx4 ,
         \CORTEXM0DS_INST/u_logic/Jyevx4 , \CORTEXM0DS_INST/u_logic/Zwevx4 ,
         \CORTEXM0DS_INST/u_logic/Pvevx4 , \CORTEXM0DS_INST/u_logic/R9fvx4 ,
         \CORTEXM0DS_INST/u_logic/Fuevx4 , \CORTEXM0DS_INST/u_logic/I4gvx4 ,
         \CORTEXM0DS_INST/u_logic/A3gvx4 , \CORTEXM0DS_INST/u_logic/Mk8vx4 ,
         \CORTEXM0DS_INST/u_logic/Aj9vx4 , \CORTEXM0DS_INST/u_logic/Bwfvx4 ,
         \CORTEXM0DS_INST/u_logic/Qufvx4 , \CORTEXM0DS_INST/u_logic/Ftfvx4 ,
         \CORTEXM0DS_INST/u_logic/Urfvx4 , \CORTEXM0DS_INST/u_logic/Jqfvx4 ,
         \CORTEXM0DS_INST/u_logic/Yofvx4 , \CORTEXM0DS_INST/u_logic/Onfvx4 ,
         \CORTEXM0DS_INST/u_logic/Emfvx4 , \CORTEXM0DS_INST/u_logic/Ukfvx4 ,
         \CORTEXM0DS_INST/u_logic/Kjfvx4 , \CORTEXM0DS_INST/u_logic/Aifvx4 ,
         \CORTEXM0DS_INST/u_logic/Qgfvx4 , \CORTEXM0DS_INST/u_logic/Gffvx4 ,
         \CORTEXM0DS_INST/u_logic/Wdfvx4 , \CORTEXM0DS_INST/u_logic/Mcfvx4 ,
         \CORTEXM0DS_INST/u_logic/Cbfvx4 , \CORTEXM0DS_INST/u_logic/Mxfvx4 ,
         \CORTEXM0DS_INST/u_logic/Xyfvx4 , \CORTEXM0DS_INST/u_logic/Ki8vx4 ,
         \CORTEXM0DS_INST/u_logic/Krgvx4 , \CORTEXM0DS_INST/u_logic/Ul8vx4 ,
         \CORTEXM0DS_INST/u_logic/Rkgvx4 , \CORTEXM0DS_INST/u_logic/Wtgvx4 ,
         \CORTEXM0DS_INST/u_logic/Hx8vx4 , \CORTEXM0DS_INST/u_logic/Vogvx4 ,
         \CORTEXM0DS_INST/u_logic/Nngvx4 , \CORTEXM0DS_INST/u_logic/Pp8vx4 ,
         \CORTEXM0DS_INST/u_logic/Mj8vx4 , \CORTEXM0DS_INST/u_logic/Q5gvx4 ,
         \CORTEXM0DS_INST/u_logic/Fjgvx4 , \CORTEXM0DS_INST/u_logic/Dmgvx4 ,
         \CORTEXM0DS_INST/u_logic/Ot9vx4 , \CORTEXM0DS_INST/u_logic/Eg8vx4 ,
         \CORTEXM0DS_INST/u_logic/Z7hvx4 , \CORTEXM0DS_INST/u_logic/Wadvx4 ,
         \CORTEXM0DS_INST/u_logic/M9dvx4 , \CORTEXM0DS_INST/u_logic/Ngdvx4 ,
         \CORTEXM0DS_INST/u_logic/Cfdvx4 , \CORTEXM0DS_INST/u_logic/Ik9vx4 ,
         \CORTEXM0DS_INST/u_logic/Yo9vx4 , \CORTEXM0DS_INST/u_logic/Vsevx4 ,
         \CORTEXM0DS_INST/u_logic/Xrdvx4 , \CORTEXM0DS_INST/u_logic/Jjdvx4 ,
         \CORTEXM0DS_INST/u_logic/Yhdvx4 , \CORTEXM0DS_INST/u_logic/Kycvx4 ,
         \CORTEXM0DS_INST/u_logic/Un9vx4 , \CORTEXM0DS_INST/u_logic/Lrevx4 ,
         \CORTEXM0DS_INST/u_logic/L9hvx4 , \CORTEXM0DS_INST/u_logic/I5dvx4 ,
         \CORTEXM0DS_INST/u_logic/Bpdvx4 , \CORTEXM0DS_INST/u_logic/Qndvx4 ,
         \CORTEXM0DS_INST/u_logic/Fmdvx4 , \CORTEXM0DS_INST/u_logic/H3evx4 ,
         \CORTEXM0DS_INST/u_logic/Izgvx4 , \CORTEXM0DS_INST/u_logic/Qm9vx4 ,
         \CORTEXM0DS_INST/u_logic/Bqevx4 , \CORTEXM0DS_INST/u_logic/Kg9vx4 ,
         \CORTEXM0DS_INST/u_logic/K5fvx4 , \CORTEXM0DS_INST/u_logic/Xlevx4 ,
         \CORTEXM0DS_INST/u_logic/Ml9vx4 , \CORTEXM0DS_INST/u_logic/B19vx4 ,
         \CORTEXM0DS_INST/u_logic/Roevx4 , \CORTEXM0DS_INST/u_logic/B5hvx4 ,
         \CORTEXM0DS_INST/u_logic/Mf8vx4 , \CORTEXM0DS_INST/u_logic/D6evx4 ,
         \CORTEXM0DS_INST/u_logic/Xq8vx4 , \CORTEXM0DS_INST/u_logic/Su9vx4 ,
         \CORTEXM0DS_INST/u_logic/Vdgvx4 , \CORTEXM0DS_INST/u_logic/Z6gvx4 ,
         \CORTEXM0DS_INST/u_logic/U9gvx4 , \CORTEXM0DS_INST/u_logic/Dbgvx4 ,
         \CORTEXM0DS_INST/u_logic/Qsgvx4 , \CORTEXM0DS_INST/u_logic/L0evx4 ,
         \CORTEXM0DS_INST/u_logic/Azdvx4 , \CORTEXM0DS_INST/u_logic/R3hvx4 ,
         \CORTEXM0DS_INST/u_logic/Mcgvx4 , \CORTEXM0DS_INST/u_logic/Efgvx4 ,
         \CORTEXM0DS_INST/u_logic/Nggvx4 , \CORTEXM0DS_INST/u_logic/Ho8vx4 ,
         \CORTEXM0DS_INST/u_logic/Ewdvx4 , \CORTEXM0DS_INST/u_logic/Tudvx4 ,
         \CORTEXM0DS_INST/u_logic/O7evx4 , \CORTEXM0DS_INST/u_logic/Uz8vx4 ,
         \CORTEXM0DS_INST/u_logic/Hnevx4 , \CORTEXM0DS_INST/u_logic/Eqgvx4 ,
         \CORTEXM0DS_INST/u_logic/Whgvx4 , \CORTEXM0DS_INST/u_logic/Cn8vx4 ,
         \CORTEXM0DS_INST/u_logic/Ih8vx4 , \CORTEXM0DS_INST/u_logic/S4evx4 ,
         \CORTEXM0DS_INST/u_logic/O8gvx4 , \CORTEXM0DS_INST/u_logic/Dw8vx4 ,
         \CORTEXM0DS_INST/u_logic/Sh9vx4 , \CORTEXM0DS_INST/u_logic/Xahvx4 ,
         n1, n2, n449, n487, n488, n1059, n1060, n1061, n1075, n1078, n1080,
         n1083, n1085, n1088, n1090, n1093, n1095, n1100, n1103, n1105, n1108,
         n1110, n1113, n1115, n1118, n1120, n1123, n1125, n1128, n1130, n1133,
         n1135, n1138, n1140, n1143, n1144, n1146, n1147, n1153, n1154, n1156,
         n1159, n1161, n1163, n1165, n1167, n1168, n1171, n1173, n1175, n1177,
         n1179, n1181, n1183, n1184, n1185, n1187, n1402, n1472, n1475, n1478,
         n1481, n1484, n1487, n1490, n1494, n1496, n1500, n1504, n1505, n1509,
         n1513, n1514, n1520, n1628, n1629, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1669, n1670, n1671, n1674, n1675, n1676, n1677, n1684,
         n1686, n1690, n1708, n1743, n1769, n1788, n1812, n1850, n1869, n1943,
         n2056, n2059, n2064, n2068, n2094, n2118, n2119, n2121, n2134, n2135,
         n2139, n2167, n2196, n2197, n2204, n2207, n2208, n2211, n2212, n2213,
         n2214, n2215, n2216, n2265, n2266, n2269, n2270, n2326, n2328, n2460,
         n2463, n2464, n2490, n2492, n2500, n2502, n2511, n2512, n2513, n2514,
         n2528, n2531, n2533, n2541, n2543, n2544, n2577, n2620, n2623, n2624,
         n2626, n2627, n2641, n2644, n2645, n2647, n2648, n2683, n2686, n2711,
         n2713, n2714, n2754, n2757, n2774, n2776, n2785, n2786, n2790, n2791,
         n2792, n2974, n2994, n2995, n3008, n3009, n3017, n3018, n3020, n3030,
         n3045, n3068, n3082, n3083, n3085, n3102, n3128, n3129, n3166, n3187,
         n3197, n3212, n3217, n3223, n3224, n3226, n3227, n3228, n3229, n3230,
         n3231, n3233, n3276, n3317, n3348, n3369, n3393, n3420, n3485, n3514,
         n3554, n3958, n3959, n3966, n3970, n3973, n4087, n4092, n4097, n4106,
         n4130, n4149, n4175, n4180, n4185, n4190, n4203, n4227, n4237, n4241,
         n4243, n4263, n4286, n4578, n4619, n4620, n4697, n4699, n4701, n4704,
         n4705, n4806, n4807, n4808, n4823, n5013, n5014, n5092, n5420, n5639,
         n5656, n5772, n5814, n5880, n5881, n5885, n5886, n5906, n5907, n5908,
         n5913, n5914, n5917, n5919, n5920, n5921, n5924, n5925, n5926, n5928,
         n5929, n5932, n5933, n5934, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6141, n6143, n6147, n6150, n6151, n6153, n6156,
         n6157, n6158, n6160, n6161, n6165, n6166, n6167, n6169, n6170, n6171,
         n6174, n6175, n6176, n6177, n6183, n6184, n6186, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748;
  wire   [31:0] PID_haddr_top;
  wire   [3:0] PID_hprot_top;
  wire   [2:0] PID_hsize_top;
  wire   [31:0] PID_hwdata_top;
  wire   [31:0] RAM_hrdata_top;
  wire   [2:0] \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state ;
  wire   [2:0] \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_nextstate ;
  wire   [4:1] \interconnect_ip_inst/i_ahb_U_mux_hsel_prev ;
  wire   [5:0] \CORTEXM0DS_INST/vis_ipsr ;
  wire   [3:0] \CORTEXM0DS_INST/vis_apsr ;
  wire   [30:0] \CORTEXM0DS_INST/vis_pc ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r14 ;
  wire   [29:0] \CORTEXM0DS_INST/vis_psp ;
  wire   [29:0] \CORTEXM0DS_INST/vis_msp ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r12 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r11 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r10 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r09 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r08 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r07 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r06 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r05 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r04 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r03 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r02 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r01 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r00 ;
  wire   [15:0] \CORTEXM0DS_INST/u_logic/L0i2z4 ;
  wire   [1:0] \CORTEXM0DS_INST/u_logic/Uth2z4 ;
  wire   [1:0] \CORTEXM0DS_INST/u_logic/Zph2z4 ;
  wire   [1:0] \CORTEXM0DS_INST/u_logic/Txh2z4 ;
  wire   [23:0] \CORTEXM0DS_INST/u_logic/Irh2z4 ;
  wire   [23:0] \CORTEXM0DS_INST/u_logic/Czh2z4 ;
  wire   [31:0] \CORTEXM0DS_INST/u_logic/Zuh2z4 ;
  wire   [15:0] \CORTEXM0DS_INST/u_logic/T1i2z4 ;
  wire   [1:0] \CORTEXM0DS_INST/u_logic/Psh2z4 ;
  wire   [3:0] \CORTEXM0DS_INST/u_logic/Tjh2z4 ;
  wire   UNCONNECTED_0;

  CPU_stub CPU_stub_inst ( .i_ssi_rxd(), .i_ssi_ss_in_n(), .i_ssi_ssi_clk(
        i_ssi_ssi_clk_top), .i_ssi_ssi_rst_n(i_ssi_ssi_rst_n_top), 
        .i_ssi_sclk_out(i_ssi_sclk_out_top), .i_ssi_ss_0_n(i_ssi_ss_0_n_top), 
        .i_ssi_ssi_mst_intr_n(i_ssi_ssi_mst_intr_n_top), .i_ssi_ssi_oe_n(
        i_ssi_ssi_oe_n_top), .i_ssi_ssi_rxf_intr_n(i_ssi_ssi_rxf_intr_n_top), 
        .i_ssi_ssi_rxo_intr_n(i_ssi_ssi_rxo_intr_n_top), 
        .i_ssi_ssi_rxu_intr_n(i_ssi_ssi_rxu_intr_n_top), .i_ssi_ssi_sleep(
        i_ssi_ssi_sleep_top), .i_ssi_ssi_txe_intr_n(i_ssi_ssi_txe_intr_n_top), 
        .i_ssi_ssi_txo_intr_n(i_ssi_ssi_intr_n_top), .i_ssi_txd(i_ssi_txd_top), 
        .HCLK(HCLK_top), .HRESETn(HRESETn_top) );
  cortexM0RAM ram2ahb_wrapper_inst ( .HCLK(HCLK_top), .HRESETn(HRESETn_top), 
        .ex_i_ahb_AHB_Slave_RAM_hrdata(RAM_hrdata_top), 
        .ex_i_ahb_AHB_Slave_RAM_hready_resp(RAM_hready_resp_top), 
        .ex_i_ahb_AHB_Slave_RAM_hresp({UNCONNECTED_0, \RAM_hresp_top[0] }), 
        .ex_i_ahb_AHB_Slave_RAM_haddr(PID_haddr_top), 
        .ex_i_ahb_AHB_Slave_RAM_hburst({1'b0, 1'b0, 1'b0}), 
        .ex_i_ahb_AHB_Slave_RAM_hmastlock(PID_hmastlock_top), 
        .ex_i_ahb_AHB_Slave_RAM_hprot({PID_hprot_top[3:2], 1'b1, 
        PID_hprot_top[0]}), .ex_i_ahb_AHB_Slave_RAM_hready(HREADY_top), 
        .ex_i_ahb_AHB_Slave_RAM_hsel(RAM_hsel_top), 
        .ex_i_ahb_AHB_Slave_RAM_hsize({1'b0, PID_hsize_top[1:0]}), 
        .ex_i_ahb_AHB_Slave_RAM_htrans({\PID_htrans_top[1] , 1'b0}), 
        .ex_i_ahb_AHB_Slave_RAM_hwdata(PID_hwdata_top), 
        .ex_i_ahb_AHB_Slave_RAM_hwrite(PID_hwrite_top) );
  nand2_1 \interconnect_ip_inst/U11942  ( .ip1(1'b0), .ip2(1'b1), .op(
        i_ssi_ssi_rxf_intr_n_top) );
  nand2_1 \interconnect_ip_inst/U11875  ( .ip1(1'b0), .ip2(1'b1), .op(
        i_ssi_ssi_txe_intr_n_top) );
  nand2_1 \interconnect_ip_inst/U11802  ( .ip1(1'b0), .ip2(1'b1), .op(
        i_ssi_ssi_rxo_intr_n_top) );
  nand2_1 \interconnect_ip_inst/U11791  ( .ip1(1'b0), .ip2(1'b1), .op(
        i_ssi_ssi_intr_n_top) );
  nand2_1 \interconnect_ip_inst/U11778  ( .ip1(1'b0), .ip2(1'b1), .op(
        i_ssi_ssi_rxu_intr_n_top) );
  nand2_1 \interconnect_ip_inst/U10788  ( .ip1(1'b0), .ip2(1'b1), .op(
        i_ssi_ssi_mst_intr_n_top) );
  nor2_1 \interconnect_ip_inst/U7231  ( .ip1(PID_haddr_top[17]), .ip2(n6111), 
        .op(RAM_hsel_top) );
  inv_1 \interconnect_ip_inst/U6038  ( .ip(1'b0), .op(i_ssi_ss_0_n_top) );
  nand2_1 \interconnect_ip_inst/U5634  ( .ip1(\interconnect_ip_inst/n6491 ), 
        .ip2(\interconnect_ip_inst/n5991 ), .op(HREADY_top) );
  drsp_1 \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_hready_resp_reg  ( .ip(
        \interconnect_ip_inst/n4829 ), .ck(HCLK_top), .rb(1'b1), .s(n12693), 
        .q(\interconnect_ip_inst/i_apb_hready_resp ) );
  drp_1 \interconnect_ip_inst/i_ssi_U_regfile_ssi_sleep_ir_reg  ( .ip(
        \interconnect_ip_inst/i_ssi_fsm_sleep ), .ck(HCLK_top), .rb(
        HRESETn_top), .q(i_ssi_ssi_sleep_top) );
  drp_1 \interconnect_ip_inst/i_ssi_U_mstfsm_fsm_sleep_reg  ( .ip(
        \interconnect_ip_inst/i_ssi_U_mstfsm_c_state[3] ), .ck(
        i_ssi_ssi_clk_top), .rb(i_ssi_ssi_rst_n_top), .q(
        \interconnect_ip_inst/i_ssi_fsm_sleep ) );
  drp_1 \interconnect_ip_inst/i_ssi_U_sclkgen_sclk_out_reg  ( .ip(1'b0), .ck(
        i_ssi_ssi_clk_top), .rb(i_ssi_ssi_rst_n_top), .q(i_ssi_sclk_out_top)
         );
  drp_1 \interconnect_ip_inst/i_ssi_U_shift_U_tx_shifter_txd_reg  ( .ip(
        i_ssi_txd_top), .ck(i_ssi_ssi_clk_top), .rb(i_ssi_ssi_rst_n_top), .q(
        i_ssi_txd_top) );
  drp_1 \interconnect_ip_inst/i_ssi_U_mstfsm_c_state_reg_3_  ( .ip(1'b1), .ck(
        i_ssi_ssi_clk_top), .rb(i_ssi_ssi_rst_n_top), .q(
        \interconnect_ip_inst/i_ssi_U_mstfsm_c_state[3] ) );
  drp_1 \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state_reg_2_  ( .ip(
        \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_nextstate [2]), .ck(
        HCLK_top), .rb(HRESETn_top), .q(
        \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state [2]) );
  drp_1 \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state_reg_0_  ( .ip(
        \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_nextstate [0]), .ck(
        HCLK_top), .rb(HRESETn_top), .q(
        \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state [0]) );
  drp_1 \interconnect_ip_inst/i_ahb_U_arblite_hmastlock_reg  ( .ip(
        \interconnect_ip_inst/n4860 ), .ck(HCLK_top), .rb(HRESETn_top), .q(
        PID_hmastlock_top) );
  drp_1 \interconnect_ip_inst/i_ahb_U_mux_hsel_prev_reg_1_  ( .ip(
        \interconnect_ip_inst/n4861 ), .ck(HCLK_top), .rb(HRESETn_top), .q(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [1]) );
  drp_1 \interconnect_ip_inst/i_ahb_U_mux_hsel_prev_reg_2_  ( .ip(
        \interconnect_ip_inst/n4862 ), .ck(HCLK_top), .rb(HRESETn_top), .q(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [2]) );
  drp_1 \interconnect_ip_inst/i_ahb_U_mux_hsel_prev_reg_3_  ( .ip(
        \interconnect_ip_inst/n4863 ), .ck(HCLK_top), .rb(HRESETn_top), .q(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [3]) );
  drp_1 \interconnect_ip_inst/i_ahb_U_mux_hsel_prev_reg_4_  ( .ip(
        \interconnect_ip_inst/n4864 ), .ck(HCLK_top), .rb(HRESETn_top), .q(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [4]) );
  drp_1 \interconnect_ip_inst/i_ahb_U_dfltslv_hresp_none_reg_0_  ( .ip(
        \interconnect_ip_inst/i_ahb_U_dfltslv_N4 ), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\interconnect_ip_inst/i_ahb_hresp_none_0_ ) );
  drp_1 \interconnect_ip_inst/i_ahb_U_dfltslv_current_state_reg  ( .ip(
        \interconnect_ip_inst/n10765 ), .ck(HCLK_top), .rb(HRESETn_top), .q(
        \interconnect_ip_inst/i_ahb_U_dfltslv_current_state ) );
  drsp_1 \interconnect_ip_inst/i_ssi_U_mstfsm_ssi_oe_n_reg  ( .ip(1'b1), .ck(
        i_ssi_ssi_clk_top), .rb(1'b1), .s(\interconnect_ip_inst/n11572 ), .q(
        i_ssi_ssi_oe_n_top) );
  drp_1 \CORTEXM0DS_INST/u_logic/J6i2z4_reg  ( .ip(n6061), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Xahvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/A4t2z4_reg  ( .ip(n6009), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Dmgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Pet2z4_reg  ( .ip(n6001), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Hx8vx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Mjl2z4_reg  ( .ip(n6060), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/B5hvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Jhy2z4_reg  ( .ip(n6042), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/V8evx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Emi2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qxhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Whgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Uqi2z4_reg  ( .ip(n6005), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Psh2z4 [1]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Zei2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Finvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/vis_apsr [1]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Gji2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/H3ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Ih8vx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Tki2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xxhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Cn8vx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Hzj2z4_reg  ( .ip(n6113), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/R3hvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Y6t2z4_reg  ( .ip(n6003), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Q5gvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/I6w2z4_reg  ( .ip(n6065), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Ul8vx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Qrp2z4_reg  ( .ip(n6007), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Txh2z4 [1]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Kop2z4_reg  ( .ip(n6062), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L9hvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/P2a3z4_reg  ( .ip(n6008), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Uth2z4 [1]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Vve3z4_reg  ( .ip(n6151), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [9]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Wbk2z4_reg  ( .ip(n6143), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Qsgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/S4w2z4_reg  ( .ip(n6002), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Rkgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/U7w2z4_reg  ( .ip(n6158), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Krgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Fed3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Efmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [4]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Nnc3z4_reg  ( .ip(n6156), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [10]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ble3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uzhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [11]) );
  drp_1 \CORTEXM0DS_INST/u_logic/D4g3z4_reg  ( .ip(n6147), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [13]) );
  drp_1 \CORTEXM0DS_INST/u_logic/T8f3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/P0ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [8]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Sgj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Owhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Efgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Vaw2z4_reg  ( .ip(n6059), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Xyfvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ffj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vwhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Nggvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Aok2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mvhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Dbgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Fij2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hwhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Mcgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/L8t2z4_reg  ( .ip(n6108), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Mj8vx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ark2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yuhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Z6gvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Nsk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ruhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Vdgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Nbm2z4_reg  ( .ip(n6109), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Xlevx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Cam2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/L8mvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/vis_ipsr [3]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Trq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pamvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/vis_ipsr [4]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Tdp2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wamvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/vis_ipsr [5]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Npk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fvhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/U9gvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Y9t2z4_reg  ( .ip(n6000), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Pp8vx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Thm2z4_reg  ( .ip(n6058), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/cm0_primask[0] ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Wxp2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/X9kvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zph2z4 [1]) );
  drp_1 \CORTEXM0DS_INST/u_logic/C3w2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ufnvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zph2z4 [0]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Dpc3z4_reg  ( .ip(n6171), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [12]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ffs2z4_reg  ( .ip(n6063), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Z7hvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/U5x2z4_reg  ( .ip(n6066), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Mk8vx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Uaj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/U9mvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/vis_ipsr [2]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Uyv2z4_reg  ( .ip(n6157), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Wtgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Nen2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ollvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/cm0_control[1] ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Idk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rhnvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/vis_apsr [0]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Lz93z4_reg  ( .ip(n6064), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/N6hvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ywi2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Owgvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Eqgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/K3l2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/F4nvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Mf8vx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Cps2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vkmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [31]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Uls2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jlmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [29]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Dks2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qlmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [28]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Tib3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lmmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [25]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Pab3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Smmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [24]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Azs2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rimvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [23]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Svs2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fjmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [21]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Bus2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mjmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [20]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Kkb3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hkmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [17]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Gcb3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Okmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [16]) );
  drp_1 \CORTEXM0DS_INST/u_logic/H8l2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ngmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [15]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Z4l2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bhmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [13]) );
  drp_1 \CORTEXM0DS_INST/u_logic/G8n2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ihmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [12]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Bmb3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dimvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [9]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Xdb3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kimvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [8]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Bjd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jemvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [7]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Vfd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xemvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [5]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Zad3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zfmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [1]) );
  drp_1 \CORTEXM0DS_INST/u_logic/J9d3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ggmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [0]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Gxk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/T2ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [0]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Vac3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/M2ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [1]) );
  drp_1 \CORTEXM0DS_INST/u_logic/F4c3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/D1ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [6]) );
  drp_1 \CORTEXM0DS_INST/u_logic/N7c3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/K1ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [5]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Oar2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nzhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [12]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ipb3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/R1ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [4]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Hub3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Y1ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [3]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Pxb3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/F2ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [2]) );
  drp_1 \CORTEXM0DS_INST/u_logic/X0c3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/W0ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [7]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ipn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/B0ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [10]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Y9l2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/I0ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [9]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Wuq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gzhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [13]) );
  drp_1 \CORTEXM0DS_INST/u_logic/V3o2z4_reg  ( .ip(n6139), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Izgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ztc3z4_reg  ( .ip(n6186), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [0]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Mcc3z4_reg  ( .ip(n6183), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [1]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Jkc3z4_reg  ( .ip(n6176), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [6]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Uic3z4_reg  ( .ip(n6174), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [5]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Fhc3z4_reg  ( .ip(n6169), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [4]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Qfc3z4_reg  ( .ip(n6167), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [3]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Bec3z4_reg  ( .ip(n6165), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [2]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ylc3z4_reg  ( .ip(n6160), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [7]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Lee3z4_reg  ( .ip(n6153), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [11]) );
  drp_1 \CORTEXM0DS_INST/u_logic/H2f3z4_reg  ( .ip(n6150), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [8]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Lns2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Clmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [30]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Jxs2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yimvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [22]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Q6l2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ugmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [14]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Lhd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qemvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [6]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Mis2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Emmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [26]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Kss2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Akmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [18]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Axm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Whmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [10]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Pcd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sfmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [2]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Tqc3z4_reg  ( .ip(n6177), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [14]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Rym2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zyhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [14]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Vgs2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xlmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [27]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Tqs2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tjmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [19]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Usl2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Phmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [11]) );
  drp_1 \CORTEXM0DS_INST/u_logic/T7d3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lfmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [3]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Lul2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Syhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [15]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Jsc3z4_reg  ( .ip(n6141), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [15]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ypi3z4_reg  ( .ip(n6112), .ck(HCLK_top), .rb(
        HRESETn_top), .q(SYSRESETREQ_top_out) );
  drp_1 \CORTEXM0DS_INST/u_logic/Aqp2z4_reg  ( .ip(n5969), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Txh2z4 [0]) );
  drp_1 \CORTEXM0DS_INST/u_logic/B1a3z4_reg  ( .ip(n5968), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Uth2z4 [0]) );
  drp_1 \CORTEXM0DS_INST/u_logic/X9n2z4_reg  ( .ip(n5967), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Psh2z4 [0]) );
  drp_1 \CORTEXM0DS_INST/u_logic/R0t2z4_reg  ( .ip(n5966), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Eg8vx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Mbt2z4_reg  ( .ip(n5965), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Nngvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Adt2z4_reg  ( .ip(n5964), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Vogvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Tna3z4_reg  ( .ip(n5963), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/F2hvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/S5b3z4_reg  ( .ip(n5962), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/S0hvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/H9i2z4_reg  ( .ip(n6010), .ck(HCLK_top), 
        .rb(1'b1), .s(\CORTEXM0DS_INST/u_logic/N586 ), .q(
        \CORTEXM0DS_INST/u_logic/Sh9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hxx2z4_reg  ( .ip(n6004), .ck(HCLK_top), 
        .rb(1'b1), .s(n12694), .q(\CORTEXM0DS_INST/u_logic/A3gvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tyx2z4_reg  ( .ip(n6104), .ck(HCLK_top), 
        .rb(1'b1), .s(\CORTEXM0DS_INST/u_logic/N586 ), .q(
        \CORTEXM0DS_INST/u_logic/I4gvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hyy2z4_reg  ( .ip(n6011), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/Cf9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I2t2z4_reg  ( .ip(n6067), .ck(HCLK_top), 
        .rb(1'b1), .s(\CORTEXM0DS_INST/u_logic/N586 ), .q(
        \CORTEXM0DS_INST/u_logic/Ot9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cqo2z4_reg  ( .ip(n6072), .ck(HCLK_top), 
        .rb(1'b1), .s(n12694), .q(\CORTEXM0DS_INST/u_logic/H3evx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Igi2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cflvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12693), .q(\CORTEXM0DS_INST/vis_apsr [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rhi2z4_reg  ( .ip(n6078), .ck(HCLK_top), 
        .rb(1'b1), .s(n12695), .q(\CORTEXM0DS_INST/u_logic/S4evx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ft73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xflvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/cm0_r02 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Iwp2z4_reg  ( .ip(n6076), .ck(HCLK_top), 
        .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/u_logic/Kycvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U4z2z4_reg  ( .ip(n6077), .ck(HCLK_top), 
        .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/u_logic/Uzcvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/S3i3z4_reg  ( .ip(n6121), .ck(HCLK_top), 
        .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bdm2z4_reg  ( .ip(n6044), .ck(HCLK_top), 
        .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/u_logic/K5fvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fcj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cxhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/vis_pc [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Swy2z4_reg  ( .ip(n6012), .ck(HCLK_top), 
        .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/u_logic/Ud9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cyq2z4_reg  ( .ip(n6105), .ck(HCLK_top), 
        .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/u_logic/Yo9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Svk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kuhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/u_logic/Xq8vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gci2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/V3ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/vis_apsr [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/V1l2z4_reg  ( .ip(n6102), .ck(HCLK_top), 
        .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/u_logic/D6evx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pdi2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Eyhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/u_logic/O8gvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/C183z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Atkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/cm0_r02 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Q7j2z4_reg  ( .ip(n6071), .ck(HCLK_top), 
        .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/Ewdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ogo2z4_reg  ( .ip(n6117), .ck(HCLK_top), 
        .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F483z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wjkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/cm0_r02 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jca3z4_reg  ( .ip(n6006), .ck(HCLK_top), 
        .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z7i2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ojnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/cm0_xpsr[24] ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/T1y2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Slnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/R9fvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jcw2z4_reg  ( .ip(n5999), .ck(HCLK_top), 
        .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/Mxfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qdj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Llnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/Ho8vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Auk2z4_reg  ( .ip(n6069), .ck(HCLK_top), 
        .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/Su9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yaz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pfhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/Nt8vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wbf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/C4ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/cm0_r00 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/G6d3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sqivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/Oy8vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/G1s2z4_reg  ( .ip(n6098), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/Wadvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kyi2z4_reg  ( .ip(n6057), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/Hnevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yzi2z4_reg  ( .ip(n6023), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/Uz8vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dq73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/E1mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/cm0_r02 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/An73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/S1mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/cm0_r02 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ohh3z4_reg  ( .ip(n6073), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/W1evx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/T583z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hfkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/cm0_r02 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z2h3z4_reg  ( .ip(n6118), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rdg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Swjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/cm0_r02 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tzg3z4_reg  ( .ip(n6088), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/Mqdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Llq2z4_reg  ( .ip(n6087), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/Xrdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ka83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/H1kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/cm0_r02 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/G0w2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Acnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/vis_ipsr [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/G9w2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lrhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Ki8vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/H3d3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/G2mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Fs8vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lbn2z4_reg  ( .ip(n6055), .ck(HCLK_top), 
        .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Bqevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Viy2z4_reg  ( .ip(n6021), .ck(HCLK_top), 
        .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/I29vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/K1z2z4_reg  ( .ip(n6070), .ck(HCLK_top), 
        .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Wv9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/An83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nrivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/cm0_r02 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yx73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/X1lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/cm0_r02 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/S8k2z4_reg  ( .ip(n6080), .ck(HCLK_top), 
        .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Azdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hak2z4_reg  ( .ip(n6079), .ck(HCLK_top), 
        .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/L0evx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jw73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/M6lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/cm0_r02 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nz73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ixkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/cm0_r02 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/H783z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sakvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/cm0_r02 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zb83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dsjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/cm0_r02 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wj83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/G5jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/cm0_r02 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dwl2z4_reg  ( .ip(n6056), .ck(HCLK_top), 
        .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/u_logic/Roevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rxl2z4_reg  ( .ip(n6022), .ck(HCLK_top), 
        .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/u_logic/B19vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Po83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ymivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/cm0_r02 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/O0o2z4_reg  ( .ip(n6120), .ck(HCLK_top), 
        .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Od83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Onjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/cm0_r02 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/E0d3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/R8ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/cm0_r00 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Df83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zijvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/cm0_r02 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qyc3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gdivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/cm0_r00 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rr73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/X0mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/cm0_r02 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wqd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cwivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r02 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wce3z4_reg  ( .ip(n6096), .ck(HCLK_top), 
        .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/u_logic/Rddvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ufy2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/G8nvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/u_logic/G8fvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gtp2z4_reg  ( .ip(n6054), .ck(HCLK_top), 
        .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/u_logic/Lrevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Owq2z4_reg  ( .ip(n6053), .ck(HCLK_top), 
        .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/u_logic/Vsevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F0y2z4_reg  ( .ip(n6052), .ck(HCLK_top), 
        .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/u_logic/Fuevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I3y2z4_reg  ( .ip(n6051), .ck(HCLK_top), 
        .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/u_logic/Pvevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/W4y2z4_reg  ( .ip(n6050), .ck(HCLK_top), 
        .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/u_logic/Zwevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/K6y2z4_reg  ( .ip(n6049), .ck(HCLK_top), 
        .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/u_logic/Jyevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Y7y2z4_reg  ( .ip(n6048), .ck(HCLK_top), 
        .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/u_logic/Tzevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M9y2z4_reg  ( .ip(n6047), .ck(HCLK_top), 
        .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/u_logic/D1fvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bby2z4_reg  ( .ip(n6046), .ck(HCLK_top), 
        .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/u_logic/O2fvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qcy2z4_reg  ( .ip(n6045), .ck(HCLK_top), 
        .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/u_logic/Z3fvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fey2z4_reg  ( .ip(n6043), .ck(HCLK_top), 
        .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/u_logic/V6fvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F1x2z4_reg  ( .ip(n6026), .ck(HCLK_top), 
        .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/u_logic/Bwfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U2x2z4_reg  ( .ip(n6025), .ck(HCLK_top), 
        .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/u_logic/Aj9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ydw2z4_reg  ( .ip(n6041), .ck(HCLK_top), 
        .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/u_logic/Cbfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mfw2z4_reg  ( .ip(n6040), .ck(HCLK_top), 
        .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/u_logic/Mcfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ahw2z4_reg  ( .ip(n6039), .ck(HCLK_top), 
        .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/u_logic/Wdfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Oiw2z4_reg  ( .ip(n6038), .ck(HCLK_top), 
        .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/u_logic/Gffvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jky2z4_reg  ( .ip(n6020), .ck(HCLK_top), 
        .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/u_logic/P39vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ckw2z4_reg  ( .ip(n6037), .ck(HCLK_top), 
        .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/u_logic/Qgfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xly2z4_reg  ( .ip(n6019), .ck(HCLK_top), 
        .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/u_logic/W49vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qlw2z4_reg  ( .ip(n6036), .ck(HCLK_top), 
        .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/u_logic/Aifvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lny2z4_reg  ( .ip(n6018), .ck(HCLK_top), 
        .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/u_logic/D69vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Enw2z4_reg  ( .ip(n6035), .ck(HCLK_top), 
        .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/u_logic/Kjfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zoy2z4_reg  ( .ip(n6017), .ck(HCLK_top), 
        .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/u_logic/K79vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sow2z4_reg  ( .ip(n6034), .ck(HCLK_top), 
        .rb(1'b1), .s(n12693), .q(\CORTEXM0DS_INST/u_logic/Ukfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nqy2z4_reg  ( .ip(n6016), .ck(HCLK_top), 
        .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/u_logic/R89vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gqw2z4_reg  ( .ip(n6033), .ck(HCLK_top), 
        .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/u_logic/Emfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bsy2z4_reg  ( .ip(n6015), .ck(HCLK_top), 
        .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Y99vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Urw2z4_reg  ( .ip(n6032), .ck(HCLK_top), 
        .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/u_logic/Onfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pty2z4_reg  ( .ip(n6014), .ck(HCLK_top), 
        .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/u_logic/Fb9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Itw2z4_reg  ( .ip(n6031), .ck(HCLK_top), 
        .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/u_logic/Yofvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dvy2z4_reg  ( .ip(n6013), .ck(HCLK_top), 
        .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/u_logic/Mc9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xuw2z4_reg  ( .ip(n6030), .ck(HCLK_top), 
        .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/u_logic/Jqfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mww2z4_reg  ( .ip(n6029), .ck(HCLK_top), 
        .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/u_logic/Urfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Byw2z4_reg  ( .ip(n6028), .ck(HCLK_top), 
        .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/u_logic/Ftfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qem2z4_reg  ( .ip(n6024), .ck(HCLK_top), 
        .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/u_logic/Kg9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/O5t2z4_reg  ( .ip(n6103), .ck(HCLK_top), 
        .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/u_logic/Fjgvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/R1w2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ocnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/vis_ipsr [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fgm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pthvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/u_logic/Tjh2z4 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wzy2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rghvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/u_logic/Tjh2z4 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sjj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Awhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/u_logic/Tjh2z4 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rni2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jxhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/u_logic/Tjh2z4 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/K9z2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wfhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/u_logic/Ks9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/W7z2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dghvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/u_logic/Gr9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I6z2z4_reg  ( .ip(n6106), .ck(HCLK_top), 
        .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/u_logic/Cq9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jwf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sdhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/vis_pc [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tme3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nehvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/vis_pc [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gmd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uehvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/vis_pc [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/V4d3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bfhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/vis_pc [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vvx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mhhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/vis_pc [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jux2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Thhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/vis_pc [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lrx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hihvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/vis_pc [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zpx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Oihvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/vis_pc [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jex2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Skhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/vis_pc [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cax2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nlhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/vis_pc [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/R8x2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ulhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/vis_pc [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/G7x2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bmhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/vis_pc [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J0l2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wthvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/vis_pc [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qzq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tinvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/u_logic/Ik9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fzl2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jdnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/u_logic/Ml9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zcn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/U2mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/u_logic/Qm9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Uup2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/N2mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/u_logic/Un9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lgi3z4_reg  ( .ip(n6081), .ck(HCLK_top), 
        .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/u_logic/Pxdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qzw2z4_reg  ( .ip(n6027), .ck(HCLK_top), 
        .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/u_logic/Qufvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wai2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lyhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/u_logic/Dw8vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/C3z2z4_reg  ( .ip(n6068), .ck(HCLK_top), 
        .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/u_logic/Bx9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/T1d3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ifhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/u_logic/Vu8vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ftf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/P7ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/cm0_r14 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Arh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ecivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r14 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/E913z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tgivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r14 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Q713z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xpivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r14 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/B613z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Muivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r14 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F8e3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bzivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r14 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kzf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/F8jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r14 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tz03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yljvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r14 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ey03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nqjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r14 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ixh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cvjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r14 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Avg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rzjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r14 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/P9h3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/G4kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r14 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bv03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rdkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r14 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nt03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gikvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r14 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zr03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vmkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r14 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fli3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zvkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r14 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wo03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/H0lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r14 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hn03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/W4lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r14 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Skh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/L9lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r14 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sl03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Aelvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r14 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Y6i3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wilvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r14 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ek03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vslvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r14 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qi03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ctlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r14 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nf03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qtlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r14 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yd03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xtlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r14 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wa03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qpivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r12 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/H903z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fuivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r12 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Q6e3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uyivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r12 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vxf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Y7jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r12 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z203z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rljvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r12 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/K103z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gqjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r12 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tvh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vujvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r12 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ltg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kzjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r12 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/A8h3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Z3kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r12 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hyz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kdkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r12 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Twz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zhkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r12 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fvz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Omkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r12 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qji3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Svkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r12 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Csz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/A0lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/cm0_r12 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nqz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/P4lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r12 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Djh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/E9lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r12 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yoz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tdlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/cm0_r12 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J5i3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pilvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/cm0_r12 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Knz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mrlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/cm0_r12 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wlz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Trlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r12 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tiz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hslvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r12 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ehz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Oslvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/cm0_r12 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qrf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/I7ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r12 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lph3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xbivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r12 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kc03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mgivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r12 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wd23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hoivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r11 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hc23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wsivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r11 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tyd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lxivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r11 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/D923z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/P6jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r11 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/K423z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ikjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r11 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/V223z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xojvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r11 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/G123z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mtjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r11 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Olg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Byjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r11 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rz13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Q2kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r11 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ow13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bckvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r11 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Av13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qgkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r11 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mt13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Flkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r11 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jq13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jukvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r11 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Uo13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rykvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r11 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fn13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/G3lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r11 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ql13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/V7lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r11 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bk13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kclvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r11 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mi13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ghlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r11 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yg13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Eulvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r11 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kf13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lulvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r11 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hc13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zulvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r11 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sa13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gvlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r11 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ilf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Z5ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r11 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mi23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Oaivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r11 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yg23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dfivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r11 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tjf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/S5ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r10 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vr33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Haivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r10 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hq33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Weivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r10 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fn33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Aoivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r10 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ql33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Psivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r10 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Exd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Exivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r10 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mi33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/I6jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r10 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Td33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bkjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r10 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ec33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qojvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r10 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pa33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ftjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r10 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zjg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uxjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r10 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/A933z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/J2kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r10 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/X533z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ubkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r10 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J433z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jgkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r10 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/V233z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ykkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r10 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sz23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cukvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r10 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dy23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kykvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r10 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ow23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Z2lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r10 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zu23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/O7lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r10 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kt23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dclvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r10 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vr23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zglvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r10 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hq23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nvlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r10 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/To23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uvlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r10 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ql23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Iwlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r10 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bk23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pwlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r10 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ow43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tnivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r09 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zu43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Isivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r09 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pvd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xwivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r09 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vr43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/B6jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r09 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cn43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ujjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r09 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nl43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jojvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r09 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yj43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ysjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r09 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kig3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nxjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r09 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ji43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/C2kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r09 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gf43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nbkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r09 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sd43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cgkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12695), .q(\CORTEXM0DS_INST/cm0_r09 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ec43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rkkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r09 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/B943z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vtkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r09 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M743z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dykvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12693), .q(\CORTEXM0DS_INST/cm0_r09 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/X543z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/S2lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r09 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I443z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/H7lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r09 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/T243z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wblvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r09 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/E143z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sglvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r09 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qz33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wwlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/cm0_r09 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cy33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dxlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/cm0_r09 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zu33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rxlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/cm0_r09 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kt33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yxlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r09 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Eif3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/L5ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r09 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/E153z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Aaivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r09 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qz43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Peivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r09 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/X563z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mnivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r08 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I463z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bsivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r08 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Aud3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qwivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r08 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/E163z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/U5jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r08 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lw53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Njjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r08 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wu53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cojvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r08 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ht53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rsjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r08 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vgg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gxjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r08 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sr53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/V1kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r08 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Po53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gbkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/cm0_r08 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bn53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vfkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r08 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nl53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kkkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/cm0_r08 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ki53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Otkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r08 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vg53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wxkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/cm0_r08 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gf53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/L2lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/cm0_r08 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rd53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/A7lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r08 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cc53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pblvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r08 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Na53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lglvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r08 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z853z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fylvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/cm0_r08 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/L753z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mylvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/cm0_r08 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I453z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Azlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12695), .q(\CORTEXM0DS_INST/cm0_r08 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/T253z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hzlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r08 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pgf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/E5ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r08 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Na63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/T9ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r08 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z863z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ieivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r08 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ajn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jpivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r07 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Oas2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ytivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r07 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/B5e3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nyivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r07 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lqr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/R7jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r07 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ozo2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kljvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r07 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Eun2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zpjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r07 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ecp2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Oujvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r07 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wrg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dzjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r07 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Eqq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/S3kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r07 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/V3m2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ddkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r07 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/G4r2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Shkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r07 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ujp2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hmkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r07 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F9j2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lvkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r07 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tel2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tzkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r07 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z3k2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/I4lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r07 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kiq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/X8lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r07 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jlo2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mdlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r07 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vuo2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Iilvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r07 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Skm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dqlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r07 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ruj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kqlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r07 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vhk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yqlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r07 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Isi2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Frlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r07 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fpi2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/B7ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r07 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rdq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qbivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r07 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cvr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fgivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r07 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bqf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/U6ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r06 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wnu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jbivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r06 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Imu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yfivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r06 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gju2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cpivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r06 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rhu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rtivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r06 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M3e3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gyivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r06 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Neu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/K7jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r06 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U9u2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dljvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r06 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F8u2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Spjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r06 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Q6u2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hujvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r06 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hqg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wyjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r06 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/B5u2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/L3kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r06 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Y1u2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wckvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r06 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/K0u2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lhkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r06 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wyt2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Amkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r06 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tvt2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Evkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r06 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Eut2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mzkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r06 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pst2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/B4lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r06 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Art2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Q8lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r06 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lpt2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fdlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r06 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wnt2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bilvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r06 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Imt2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uolvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r06 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ukt2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bplvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r06 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rht2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pplvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r06 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cgt2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wplvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r06 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mhn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Voivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r05 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z8s2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ktivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r05 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/X1e3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zxivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r05 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wor2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/D7jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r05 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zxo2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wkjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r05 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Psn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lpjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r05 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pap2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Aujvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r05 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sog3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pyjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r05 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Poq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/E3kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r05 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/H2m2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pckvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r05 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/S2r2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ehkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r05 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gip2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tlkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r05 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vmj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xukvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r05 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Edl2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fzkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r05 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/K2k2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/U3lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r05 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vgq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/J8lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r05 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ujo2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yclvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r05 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gto2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uhlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r05 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ejm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lnlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r05 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dtj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Snlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r05 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ggk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Golvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r05 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Glj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nolvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r05 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mof3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/N6ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r05 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ccq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cbivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r05 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Otr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rfivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r05 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Psv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ooivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r04 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Arv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dtivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r04 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I0e3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sxivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r04 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wnv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/W6jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r04 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Djv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pkjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r04 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ohv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Epjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r04 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zfv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ttjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r04 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dng3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Iyjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r04 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kev2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/X2kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r04 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hbv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ickvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r04 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/T9v2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xgkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r04 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F8v2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mlkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r04 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/C5v2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qukvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r04 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/N3v2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yykvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r04 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Y1v2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/N3lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r04 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J0v2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/C8lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r04 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Uyu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rclvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r04 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fxu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nhlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r04 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rvu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cmlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r04 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Duu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jmlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r04 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Aru2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xmlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r04 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lpu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Enlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r04 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xmf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/G6ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r04 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fxv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vaivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r04 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rvv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kfivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r04 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gf73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fnivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r03 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rd73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Urivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r03 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lsd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jwivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r03 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Na73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/N5jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r03 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U573z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gjjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/cm0_r03 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F473z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vnjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_r03 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Q273z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ksjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(
        \CORTEXM0DS_INST/u_logic/N586 ), .q(\CORTEXM0DS_INST/cm0_r03 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gfg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zwjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/cm0_r03 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/B173z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/O1kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_r03 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yx63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zakvx4 ), .ck(HCLK_top), .rb(1'b1), .s(
        \CORTEXM0DS_INST/u_logic/N586 ), .q(\CORTEXM0DS_INST/cm0_r03 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kw63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ofkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r03 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wu63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dkkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_r03 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tr63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Htkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(
        \CORTEXM0DS_INST/u_logic/N586 ), .q(\CORTEXM0DS_INST/cm0_r03 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Eq63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pxkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r03 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Po63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/E2lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_r03 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/An63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/T6lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(
        \CORTEXM0DS_INST/u_logic/N586 ), .q(\CORTEXM0DS_INST/cm0_r03 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ll63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Iblvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r03 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wj63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Eglvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r03 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ii63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ozlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r03 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ug63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vzlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r03 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rd63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/J0mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r03 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cc63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Q0mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r03 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Aff3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/X4ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r03 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wj73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/M9ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r03 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ii73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Beivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r03 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ldf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Q4ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r02 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ft83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/F9ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r02 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rr83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Udivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r02 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Uu73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bblvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r02 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ll73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Z1mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r02 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yfn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rmivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r01 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/K7s2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Grivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r01 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hpd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vvivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r01 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hnr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Z4jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r01 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kwo2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sijvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r01 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Arn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hnjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r01 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/A9p2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wrjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r01 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ccg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lwjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r01 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Anq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/A1kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r01 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/T0m2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lakvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r01 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/E1r2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Afkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/cm0_r01 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sgp2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pjkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/cm0_r01 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zpj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tskvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r01 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pbl2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bxkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r01 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/V0k2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Q1lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r01 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gfq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/F6lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/cm0_r01 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fio2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ualvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/cm0_r01 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rro2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qflvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/cm0_r01 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gmm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Eenvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/cm0_r01 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fwj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lenvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/cm0_r01 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kjk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zenvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/cm0_r01 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Koj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gfnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/cm0_r01 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Orj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/J4ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r01 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Naq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Y8ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r01 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Asr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ndivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r01 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vu93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kmivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r00 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gt93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zqivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r00 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Snd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ovivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r00 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cq93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/S4jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r00 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Uj93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lijvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r00 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fi93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Anjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r00 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qg93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Prjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r00 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nag3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ewjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r00 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bf93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/T0kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r00 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yb93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Eakvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/cm0_r00 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ka93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tekvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r00 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/W893z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ijkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/cm0_r00 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/R293z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mskvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/cm0_r00 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/C193z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uwkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/cm0_r00 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nz83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/J1lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r00 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yx83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Y5lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r00 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jw83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nalvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r00 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Uu83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jflvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r00 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Unm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bgnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/cm0_r00 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xti2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wgnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r00 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zkk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dhnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r00 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Txj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Minvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/cm0_r00 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/B9g3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ldhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/vis_pc [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bnx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cjhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/vis_pc [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Plx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jjhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/vis_pc [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zjq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ithvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/vis_pc [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fhx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ekhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/vis_pc [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dkr2z4_reg  ( .ip(n6095), .ck(HCLK_top), 
        .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/u_logic/Cfdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/S703z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/J3jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/cm0_r12 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kfr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/C3jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/cm0_r07 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vdr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/O2jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/cm0_r05 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lpv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/H2jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/cm0_r04 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sa23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/A2jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/cm0_r11 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kt43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/M1jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/cm0_r09 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/T263z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/F1jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/cm0_r08 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cc73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Y0jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/cm0_r03 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gcr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/K0jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/cm0_r01 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rr93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/D0jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/cm0_r00 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M413z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Q3jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/cm0_r14 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cgu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/V2jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/cm0_r06 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bk33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/T1jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/cm0_r10 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ll83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/R0jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/cm0_r02 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ycx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zkhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/vis_pc [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ikz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Aslvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/cm0_r12 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Eol2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rqlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/cm0_r07 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qml2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Znlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/cm0_r05 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Psu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qmlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/cm0_r04 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wd13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sulvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/cm0_r11 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ow33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kxlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/cm0_r09 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/X553z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tylvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/cm0_r08 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gf63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/C0mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/cm0_r03 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Spl2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Senvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/cm0_r01 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Grl2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ignvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/cm0_r00 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ch03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jtlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/cm0_r14 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gjt2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Iplvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/cm0_r06 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fn23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bwlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/cm0_r10 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Po73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/L1mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/cm0_r02 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I793z4_reg  ( .ip(n6074), .ck(HCLK_top), 
        .rb(1'b1), .s(n12694), .q(\CORTEXM0DS_INST/u_logic/C8dvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Szr2z4_reg  ( .ip(n6099), .ck(HCLK_top), 
        .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/M9dvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rpe3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Blivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12693), .q(\CORTEXM0DS_INST/cm0_r12 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/W5s2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ukivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12695), .q(\CORTEXM0DS_INST/cm0_r07 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I4s2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gkivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r05 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Duv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zjivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r04 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kf23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sjivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r11 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cy43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ejivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r09 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/L763z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xiivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r08 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ug73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qiivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r03 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U2s2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ciivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r01 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cxc3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vhivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r00 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fre3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ilivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/cm0_r14 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Uku2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nkivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/cm0_r06 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/To33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ljivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/cm0_r10 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dq83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jiivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/cm0_r02 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ufx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lkhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/vis_pc [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rkd3z4_reg  ( .ip(n6097), .ck(HCLK_top), 
        .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/u_logic/Gcdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J4x2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Imhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/vis_pc [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M1j2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hllvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/u_logic/O7evx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Eyr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hhivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/vis_psp [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hue3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wlivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/vis_psp [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cmn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lqivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/vis_psp [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rds2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Avivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/vis_psp [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ibe3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pzivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_psp [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Oir2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/E4jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_psp [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/O2g3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/T8jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_psp [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/S2p2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mmjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_psp [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ixn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Brjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_psp [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M0i3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qvjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_psp [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Eyg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/F0kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_psp [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tch3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/U4kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_psp [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/X6m2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fekvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_psp [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I7r2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uikvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_psp [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wmp2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jnkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_psp [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Joi3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nwkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_psp [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xhl2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/V0lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/vis_psp [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/D7k2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/K5lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/vis_psp [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wnh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Z9lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/vis_psp [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Noo2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Oelvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/vis_psp [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cai3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kjlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/vis_psp [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pfz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mklvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/vis_psp [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Aez2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tklvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/vis_psp [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mcz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Allvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/vis_psp [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Uuf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/D8ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/vis_psp [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Euh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Scivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/vis_psp [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tse3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Plivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/vis_msp [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Okn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Eqivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/vis_msp [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dcs2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tuivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/vis_msp [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U9e3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Izivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/vis_msp [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zgr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/X3jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/vis_msp [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z0g3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/M8jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/vis_msp [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/D1p2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fmjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/vis_msp [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tvn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uqjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/vis_msp [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xyh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jvjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/vis_msp [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pwg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yzjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/vis_msp [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ebh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/N4kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/vis_msp [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J5m2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ydkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/vis_msp [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U5r2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nikvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/vis_msp [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ilp2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cnkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/vis_msp [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Umi3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gwkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/vis_msp [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Igl2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/O0lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/vis_msp [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/O5k2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/D5lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/vis_msp [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hmh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/S9lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/vis_msp [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ymo2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Helvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/vis_msp [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/N8i3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Djlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/vis_msp [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/X2j2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rjlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/vis_msp [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rek2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yjlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/vis_msp [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cll2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fklvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/vis_msp [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M4j2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/W7ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/vis_msp [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Psh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lcivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/vis_msp [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qwr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ahivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/vis_msp [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Slr2z4_reg  ( .ip(n6094), .ck(HCLK_top), 
        .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/u_logic/Ngdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rbi3z4_reg  ( .ip(n6107), .ck(HCLK_top), 
        .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/u_logic/H0gvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jw93z4_reg  ( .ip(n6075), .ck(HCLK_top), 
        .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/u_logic/E1dvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xx93z4_reg  ( .ip(n6085), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/O2dvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ovc3z4_reg  ( .ip(n6084), .ck(HCLK_top), 
        .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/u_logic/Y3dvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Efp2z4_reg  ( .ip(n6083), .ck(HCLK_top), 
        .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/u_logic/I5dvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F2o2z4_reg  ( .ip(n6138), .ck(HCLK_top), 
        .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/C4b3z4_reg  ( .ip(n6137), .ck(HCLK_top), 
        .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M2b3z4_reg  ( .ip(n6136), .ck(HCLK_top), 
        .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/W0b3z4_reg  ( .ip(n6135), .ck(HCLK_top), 
        .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gza3z4_reg  ( .ip(n6134), .ck(HCLK_top), 
        .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qxa3z4_reg  ( .ip(n6133), .ck(HCLK_top), 
        .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z8b3z4_reg  ( .ip(n6132), .ck(HCLK_top), 
        .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dhb3z4_reg  ( .ip(n6131), .ck(HCLK_top), 
        .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M5f3z4_reg  ( .ip(n6130), .ck(HCLK_top), 
        .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Aze3z4_reg  ( .ip(n6129), .ck(HCLK_top), 
        .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zva3z4_reg  ( .ip(n6128), .ck(HCLK_top), 
        .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/She3z4_reg  ( .ip(n6127), .ck(HCLK_top), 
        .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Iua3z4_reg  ( .ip(n6126), .ck(HCLK_top), 
        .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/K7g3z4_reg  ( .ip(n6125), .ck(HCLK_top), 
        .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ddi3z4_reg  ( .ip(n6116), .ck(HCLK_top), 
        .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Uei3z4_reg  ( .ip(n6115), .ck(HCLK_top), 
        .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nbx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Glhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/vis_pc [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ytm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rrkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/vis_msp [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rtz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Drkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r12 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ksm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wqkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/cm0_r07 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wqm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Iqkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/cm0_r05 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/R6v2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bqkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/cm0_r04 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yr13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Upkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r11 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qa43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gpkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/cm0_r09 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zj53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zokvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r08 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/It63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sokvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/cm0_r03 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ipm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Eokvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r01 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/G493z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xnkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r00 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mvm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yrkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(
        \CORTEXM0DS_INST/u_logic/N586 ), .q(\CORTEXM0DS_INST/vis_psp [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lq03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Krkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r14 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ixt2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pqkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/cm0_r06 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/H133z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Npkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/cm0_r10 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/R283z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lokvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/cm0_r02 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dkx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qjhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/vis_pc [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cao2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qhjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/vis_msp [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/O403z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Chjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/cm0_r12 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/N8o2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vgjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/cm0_r07 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Y6o2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hgjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/cm0_r05 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Skv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Agjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/cm0_r04 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z523z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tfjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/cm0_r11 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ro43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ffjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/cm0_r09 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ay53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yejvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/cm0_r08 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J773z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rejvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/cm0_r03 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J5o2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dejvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/cm0_r01 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jl93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wdjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r00 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rbo2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xhjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(
        \CORTEXM0DS_INST/u_logic/N586 ), .q(\CORTEXM0DS_INST/vis_psp [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I113z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jhjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r14 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jbu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ogjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r06 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/If33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mfjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r10 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sg83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kejvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r02 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nox2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vihvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/vis_pc [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/C5n2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/C9kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_msp [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vzz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/O8kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r12 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/N3n2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/H8kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r07 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Y1n2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/T7kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/cm0_r05 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vcv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/M7kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/cm0_r04 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cy13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/F7kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/cm0_r11 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ug43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/R6kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/cm0_r09 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dq53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/K6kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/cm0_r08 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mz63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/D6kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/cm0_r03 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J0n2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/P5kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/cm0_r01 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Md93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/I5kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/cm0_r00 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/R6n2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/J9kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/vis_psp [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pw03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/V8kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/cm0_r14 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M3u2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/A8kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/cm0_r06 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/L733z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Y6kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/cm0_r10 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/V883z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/W5kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/cm0_r02 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rix2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xjhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/vis_pc [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F4q2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bdjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/vis_msp [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/D603z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ncjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r12 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Q2q2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gcjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r07 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/B1q2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sbjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r05 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hmv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lbjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/cm0_r04 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/O723z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ebjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r11 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gq43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qajvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/cm0_r09 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pz53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jajvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/cm0_r08 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Y873z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cajvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/cm0_r03 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mzp2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/O9jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r01 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/No93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/H9jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/cm0_r00 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U5q2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Idjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/vis_psp [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/X213z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ucjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/cm0_r14 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ycu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zbjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/cm0_r06 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xg33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xajvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/cm0_r10 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hi83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/V9jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/cm0_r02 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J7q2z4_reg  ( .ip(n6093), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/Yhdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Y8q2z4_reg  ( .ip(n6100), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/Jjdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rsa3z4_reg  ( .ip(n6124), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zfh3z4_reg  ( .ip(n6086), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/Itdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ym93z4_reg  ( .ip(n6092), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/Ukdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xeo2z4_reg  ( .ip(n6122), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xyk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Duhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12695), .q(\CORTEXM0DS_INST/vis_pc [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U593z4_reg  ( .ip(n6082), .ck(HCLK_top), 
        .rb(1'b1), .s(n12695), .q(\CORTEXM0DS_INST/u_logic/S6dvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kaf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zdhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12695), .q(\CORTEXM0DS_INST/vis_pc [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/H4p2z4_reg  ( .ip(n6091), .ck(HCLK_top), 
        .rb(1'b1), .s(n12695), .q(\CORTEXM0DS_INST/u_logic/Fmdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ara3z4_reg  ( .ip(n6123), .ck(HCLK_top), 
        .rb(1'b1), .s(n12695), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/W5p2z4_reg  ( .ip(n6090), .ck(HCLK_top), 
        .rb(1'b1), .s(n12695), .q(\CORTEXM0DS_INST/u_logic/Qndvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Foe3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gehvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12695), .q(\CORTEXM0DS_INST/vis_pc [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/L7p2z4_reg  ( .ip(n6089), .ck(HCLK_top), 
        .rb(1'b1), .s(n12695), .q(\CORTEXM0DS_INST/u_logic/Bpdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jpa3z4_reg  ( .ip(n6119), .ck(HCLK_top), 
        .rb(1'b1), .s(n12695), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xsx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Aihvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12695), .q(\CORTEXM0DS_INST/vis_pc [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Omk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tvhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12695), .q(\CORTEXM0DS_INST/vis_pc [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/B6j2z4_reg  ( .ip(n6101), .ck(HCLK_top), 
        .rb(1'b1), .s(n12695), .q(\CORTEXM0DS_INST/u_logic/Tudvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/B2i3z4_reg  ( .ip(n5961), .ck(HCLK_top), 
        .rb(1'b1), .s(n12694), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ieh3z4_reg  ( .ip(n5960), .ck(HCLK_top), 
        .rb(1'b1), .s(n12694), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kxe3z4_reg  ( .ip(n5959), .ck(HCLK_top), 
        .rb(1'b1), .s(n12694), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I1h3z4_reg  ( .ip(n5958), .ck(HCLK_top), 
        .rb(1'b1), .s(n12694), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cma3z4_reg  ( .ip(n5957), .ck(HCLK_top), 
        .rb(1'b1), .s(n12694), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/C9a3z4_reg  ( .ip(n5956), .ck(HCLK_top), 
        .rb(1'b1), .s(n12694), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bge3z4_reg  ( .ip(n5955), .ck(HCLK_top), 
        .rb(1'b1), .s(n12694), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/T5g3z4_reg  ( .ip(n5954), .ck(HCLK_top), 
        .rb(1'b1), .s(n12694), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xyn2z4_reg  ( .ip(n5953), .ck(HCLK_top), 
        .rb(1'b1), .s(n12694), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/W3f3z4_reg  ( .ip(n5952), .ck(HCLK_top), 
        .rb(1'b1), .s(n12694), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Aea3z4_reg  ( .ip(n5951), .ck(HCLK_top), 
        .rb(1'b1), .s(n12694), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wia3z4_reg  ( .ip(n5950), .ck(HCLK_top), 
        .rb(1'b1), .s(n12694), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J7b3z4_reg  ( .ip(n5949), .ck(HCLK_top), 
        .rb(1'b1), .s(n12693), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qfa3z4_reg  ( .ip(n5948), .ck(HCLK_top), 
        .rb(1'b1), .s(n12693), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mka3z4_reg  ( .ip(n5947), .ck(HCLK_top), 
        .rb(1'b1), .s(n12693), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Taa3z4_reg  ( .ip(n5946), .ck(HCLK_top), 
        .rb(1'b1), .s(n12693), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gha3z4_reg  ( .ip(n5945), .ck(HCLK_top), 
        .rb(1'b1), .s(n12693), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nfb3z4_reg  ( .ip(n5944), .ck(HCLK_top), 
        .rb(1'b1), .s(n12693), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/L7a3z4_reg  ( .ip(n5943), .ck(HCLK_top), 
        .rb(1'b1), .s(n12693), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U5a3z4_reg  ( .ip(n5942), .ck(HCLK_top), 
        .rb(1'b1), .s(n12693), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gdo2z4_reg  ( .ip(n5941), .ck(HCLK_top), 
        .rb(1'b1), .s(n12693), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/D4a3z4_reg  ( .ip(n5940), .ck(HCLK_top), 
        .rb(1'b1), .s(n12693), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/L8m2z4_reg  ( .ip(n5939), .ck(HCLK_top), 
        .rb(1'b1), .s(n12693), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [19]) );
  mux2_1 U8 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [19]), .ip2(
        PID_hwdata_top[19]), .s(n12691), .op(n5939) );
  mux2_1 U10 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [15]), .ip2(
        PID_hwdata_top[15]), .s(n12692), .op(n5940) );
  mux2_1 U11 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [16]), .ip2(
        PID_hwdata_top[16]), .s(n12691), .op(n5941) );
  mux2_1 U12 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [14]), .ip2(
        PID_hwdata_top[14]), .s(n12691), .op(n5942) );
  mux2_1 U13 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [12]), .ip2(
        PID_hwdata_top[12]), .s(n12691), .op(n5943) );
  mux2_1 U14 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [7]), .ip2(
        PID_hwdata_top[7]), .s(n12691), .op(n5944) );
  mux2_1 U15 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [2]), .ip2(
        PID_hwdata_top[2]), .s(n12691), .op(n5945) );
  mux2_1 U16 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [4]), .ip2(
        PID_hwdata_top[4]), .s(n12691), .op(n5946) );
  mux2_1 U17 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [5]), .ip2(
        PID_hwdata_top[5]), .s(n12691), .op(n5947) );
  mux2_1 U18 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [1]), .ip2(
        PID_hwdata_top[1]), .s(n12691), .op(n5948) );
  mux2_1 U19 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [6]), .ip2(
        PID_hwdata_top[6]), .s(n12691), .op(n5949) );
  mux2_1 U20 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [3]), .ip2(
        PID_hwdata_top[3]), .s(n12691), .op(n5950) );
  mux2_1 U21 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [0]), .ip2(
        PID_hwdata_top[0]), .s(n12692), .op(n5951) );
  mux2_1 U22 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [8]), .ip2(
        PID_hwdata_top[8]), .s(n12692), .op(n5952) );
  mux2_1 U23 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [18]), .ip2(
        PID_hwdata_top[18]), .s(n12692), .op(n5953) );
  mux2_1 U24 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [13]), .ip2(
        PID_hwdata_top[13]), .s(n12692), .op(n5954) );
  mux2_1 U25 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [11]), .ip2(
        PID_hwdata_top[11]), .s(n12692), .op(n5955) );
  mux2_1 U26 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [10]), .ip2(
        PID_hwdata_top[10]), .s(n12692), .op(n5956) );
  mux2_1 U27 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [22]), .ip2(
        PID_hwdata_top[22]), .s(n12692), .op(n5957) );
  mux2_1 U28 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [20]), .ip2(
        PID_hwdata_top[20]), .s(n12692), .op(n5958) );
  mux2_1 U29 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [9]), .ip2(
        PID_hwdata_top[9]), .s(n12692), .op(n5959) );
  mux2_1 U30 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [21]), .ip2(
        PID_hwdata_top[21]), .s(n12692), .op(n5960) );
  mux2_1 U31 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [17]), .ip2(
        PID_hwdata_top[17]), .s(n12692), .op(n5961) );
  mux2_1 U35 ( .ip1(\CORTEXM0DS_INST/u_logic/S0hvx4 ), .ip2(PID_hwdata_top[1]), 
        .s(n1), .op(n5962) );
  inv_1 U36 ( .ip(HRESETn_top), .op(\CORTEXM0DS_INST/u_logic/N586 ) );
  mux2_1 U37 ( .ip1(\CORTEXM0DS_INST/u_logic/F2hvx4 ), .ip2(PID_hwdata_top[0]), 
        .s(n1), .op(n5963) );
  mux2_1 U41 ( .ip1(\CORTEXM0DS_INST/u_logic/Vogvx4 ), .ip2(PID_hwdata_top[4]), 
        .s(n2), .op(n5964) );
  mux2_1 U42 ( .ip1(\CORTEXM0DS_INST/u_logic/Nngvx4 ), .ip2(PID_hwdata_top[2]), 
        .s(n2), .op(n5965) );
  mux2_1 U43 ( .ip1(\CORTEXM0DS_INST/u_logic/Eg8vx4 ), .ip2(PID_hwdata_top[1]), 
        .s(n2), .op(n5966) );
  mux2_1 U47 ( .ip1(PID_hwdata_top[22]), .ip2(
        \CORTEXM0DS_INST/u_logic/Psh2z4 [0]), .s(n487), .op(n5967) );
  mux2_1 U52 ( .ip1(\CORTEXM0DS_INST/u_logic/Uth2z4 [0]), .ip2(
        PID_hwdata_top[30]), .s(n488), .op(n5968) );
  mux2_1 U53 ( .ip1(PID_hwdata_top[30]), .ip2(
        \CORTEXM0DS_INST/u_logic/Txh2z4 [0]), .s(n487), .op(n5969) );
  mux2_1 U646 ( .ip1(\RAM_hresp_top[0] ), .ip2(
        \interconnect_ip_inst/i_ahb_hresp_none_0_ ), .s(n5920), .op(n449) );
  nand2_1 U649 ( .ip1(HREADY_top), .ip2(\CORTEXM0DS_INST/u_logic/Xyfvx4 ), 
        .op(n1185) );
  inv_1 U651 ( .ip(HREADY_top), .op(n5932) );
  mux2_1 U652 ( .ip1(PID_hwrite_top), .ip2(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), 
        .s(n5932), .op(n6000) );
  nand2_1 U798 ( .ip1(\CORTEXM0DS_INST/u_logic/Mf8vx4 ), .ip2(
        PID_hwdata_top[23]), .op(n3226) );
  nand2_1 U802 ( .ip1(\CORTEXM0DS_INST/u_logic/Mf8vx4 ), .ip2(
        PID_hwdata_top[31]), .op(n3227) );
  nand2_1 U994 ( .ip1(HREADY_top), .ip2(PID_hprot_top[0]), .op(n4578) );
  ab_or_c_or_d U1586 ( .ip1(n1060), .ip2(n5639), .ip3(HREADY_top), .ip4(n1059), 
        .op(n1061) );
  nand2_1 U1595 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(HREADY_top), 
        .op(n1708) );
  nand2_1 U1599 ( .ip1(RAM_hrdata_top[14]), .ip2(n1147), .op(n1075) );
  inv_1 U1602 ( .ip(RAM_hrdata_top[30]), .op(n1156) );
  nand2_1 U1612 ( .ip1(RAM_hrdata_top[12]), .ip2(n1147), .op(n1080) );
  nand2_1 U1616 ( .ip1(RAM_hrdata_top[28]), .ip2(n1143), .op(n1078) );
  nand2_1 U1618 ( .ip1(RAM_hrdata_top[27]), .ip2(n1143), .op(n1085) );
  nand2_1 U1623 ( .ip1(RAM_hrdata_top[11]), .ip2(n1147), .op(n1083) );
  nand2_1 U1625 ( .ip1(RAM_hrdata_top[26]), .ip2(n1143), .op(n1090) );
  nand2_1 U1630 ( .ip1(RAM_hrdata_top[10]), .ip2(n1147), .op(n1088) );
  nand2_1 U1632 ( .ip1(RAM_hrdata_top[9]), .ip2(n1147), .op(n1095) );
  nand2_1 U1638 ( .ip1(RAM_hrdata_top[25]), .ip2(n1143), .op(n1093) );
  nand2_1 U1640 ( .ip1(RAM_hrdata_top[8]), .ip2(n1147), .op(n1100) );
  inv_1 U1641 ( .ip(RAM_hrdata_top[24]), .op(n1168) );
  nand2_1 U1648 ( .ip1(RAM_hrdata_top[23]), .ip2(n1143), .op(n1105) );
  nand2_1 U1652 ( .ip1(RAM_hrdata_top[7]), .ip2(n1147), .op(n1103) );
  nand2_1 U1654 ( .ip1(RAM_hrdata_top[22]), .ip2(n1143), .op(n1110) );
  nand2_1 U1659 ( .ip1(RAM_hrdata_top[6]), .ip2(n1147), .op(n1108) );
  nand2_1 U1661 ( .ip1(RAM_hrdata_top[21]), .ip2(n1143), .op(n1115) );
  nand2_1 U1667 ( .ip1(RAM_hrdata_top[5]), .ip2(n1147), .op(n1113) );
  nand2_1 U1669 ( .ip1(RAM_hrdata_top[20]), .ip2(n1143), .op(n1120) );
  nand2_1 U1675 ( .ip1(RAM_hrdata_top[4]), .ip2(n1147), .op(n1118) );
  nand2_1 U1677 ( .ip1(RAM_hrdata_top[19]), .ip2(n1143), .op(n1125) );
  nand2_1 U1683 ( .ip1(RAM_hrdata_top[3]), .ip2(n1147), .op(n1123) );
  nand2_1 U1685 ( .ip1(RAM_hrdata_top[18]), .ip2(n1143), .op(n1130) );
  nand2_1 U1691 ( .ip1(RAM_hrdata_top[2]), .ip2(n1147), .op(n1128) );
  nand2_1 U1693 ( .ip1(RAM_hrdata_top[17]), .ip2(n1143), .op(n1135) );
  nand2_1 U1699 ( .ip1(RAM_hrdata_top[1]), .ip2(n1147), .op(n1133) );
  nand2_1 U1701 ( .ip1(RAM_hrdata_top[16]), .ip2(n1143), .op(n1140) );
  nand2_1 U1707 ( .ip1(RAM_hrdata_top[0]), .ip2(n1147), .op(n1138) );
  nand2_1 U1709 ( .ip1(RAM_hrdata_top[13]), .ip2(n1147), .op(n1146) );
  nand2_1 U1714 ( .ip1(RAM_hrdata_top[29]), .ip2(n1143), .op(n1144) );
  nand2_1 U1716 ( .ip1(RAM_hrdata_top[15]), .ip2(n1147), .op(n1153) );
  inv_1 U1717 ( .ip(RAM_hrdata_top[31]), .op(n1154) );
  nand2_1 U1728 ( .ip1(RAM_hrdata_top[29]), .ip2(n1184), .op(n1159) );
  nand2_1 U1731 ( .ip1(RAM_hrdata_top[28]), .ip2(n1184), .op(n1161) );
  nand2_1 U1734 ( .ip1(RAM_hrdata_top[27]), .ip2(n1184), .op(n1163) );
  nand2_1 U1737 ( .ip1(RAM_hrdata_top[26]), .ip2(n1184), .op(n1165) );
  nand2_1 U1740 ( .ip1(RAM_hrdata_top[25]), .ip2(n1184), .op(n1167) );
  nand2_1 U1745 ( .ip1(RAM_hrdata_top[23]), .ip2(n1184), .op(n1171) );
  nand2_1 U1748 ( .ip1(RAM_hrdata_top[22]), .ip2(n1184), .op(n1173) );
  nand2_1 U1751 ( .ip1(RAM_hrdata_top[21]), .ip2(n1184), .op(n1175) );
  nand2_1 U1754 ( .ip1(RAM_hrdata_top[20]), .ip2(n1184), .op(n1177) );
  nand2_1 U1757 ( .ip1(RAM_hrdata_top[19]), .ip2(n1184), .op(n1179) );
  nand2_1 U1760 ( .ip1(RAM_hrdata_top[18]), .ip2(n1184), .op(n1181) );
  nand2_1 U1763 ( .ip1(RAM_hrdata_top[17]), .ip2(n1184), .op(n1183) );
  nand2_1 U1766 ( .ip1(RAM_hrdata_top[16]), .ip2(n1184), .op(n1187) );
  nand2_1 U2030 ( .ip1(n1513), .ip2(RAM_hrdata_top[14]), .op(n1402) );
  nand2_1 U2032 ( .ip1(RAM_hrdata_top[13]), .ip2(n1513), .op(n1472) );
  nand2_1 U2082 ( .ip1(RAM_hrdata_top[12]), .ip2(n1513), .op(n1475) );
  nand2_1 U2086 ( .ip1(RAM_hrdata_top[11]), .ip2(n1513), .op(n1478) );
  nand2_1 U2090 ( .ip1(RAM_hrdata_top[10]), .ip2(n1513), .op(n1481) );
  nand2_1 U2094 ( .ip1(RAM_hrdata_top[9]), .ip2(n1513), .op(n1484) );
  nand2_1 U2098 ( .ip1(RAM_hrdata_top[8]), .ip2(n1513), .op(n1487) );
  nand2_1 U2102 ( .ip1(RAM_hrdata_top[7]), .ip2(n1513), .op(n1490) );
  nand2_1 U2106 ( .ip1(RAM_hrdata_top[6]), .ip2(n1513), .op(n1494) );
  nand2_1 U2113 ( .ip1(n1513), .ip2(RAM_hrdata_top[5]), .op(n1496) );
  nand2_1 U2115 ( .ip1(RAM_hrdata_top[4]), .ip2(n1513), .op(n1500) );
  nand2_1 U2119 ( .ip1(RAM_hrdata_top[3]), .ip2(n1513), .op(n1504) );
  nand2_1 U2125 ( .ip1(RAM_hrdata_top[2]), .ip2(n1513), .op(n1505) );
  nand2_1 U2128 ( .ip1(RAM_hrdata_top[1]), .ip2(n1513), .op(n1509) );
  nand2_1 U2133 ( .ip1(RAM_hrdata_top[0]), .ip2(n1513), .op(n1514) );
  nor2_1 U2139 ( .ip1(PID_hprot_top[0]), .ip2(n1520), .op(n2211) );
  nand3_1 U2265 ( .ip1(PID_haddr_top[29]), .ip2(PID_haddr_top[30]), .ip3(
        PID_haddr_top[31]), .op(n2207) );
  nor3_1 U2270 ( .ip1(PID_haddr_top[5]), .ip2(PID_haddr_top[9]), .ip3(
        PID_haddr_top[7]), .op(n1671) );
  inv_1 U2271 ( .ip(PID_haddr_top[8]), .op(n1629) );
  nor3_1 U2273 ( .ip1(PID_haddr_top[3]), .ip2(PID_haddr_top[4]), .ip3(n2068), 
        .op(n1628) );
  not_ab_or_c_or_d U2274 ( .ip1(PID_haddr_top[11]), .ip2(n1629), .ip3(n1628), 
        .ip4(PID_haddr_top[6]), .op(n1663) );
  nand3_1 U2310 ( .ip1(n2064), .ip2(PID_haddr_top[10]), .ip3(n1850), .op(n1661) );
  nand2_1 U2311 ( .ip1(PID_haddr_top[8]), .ip2(n1661), .op(n1662) );
  nor2_1 U2313 ( .ip1(PID_haddr_top[8]), .ip2(PID_haddr_top[9]), .op(n1664) );
  not_ab_or_c_or_d U2314 ( .ip1(PID_haddr_top[8]), .ip2(PID_haddr_top[9]), 
        .ip3(PID_haddr_top[6]), .ip4(n1664), .op(n1674) );
  nor2_1 U2315 ( .ip1(PID_haddr_top[9]), .ip2(PID_haddr_top[7]), .op(n1665) );
  nand3_1 U2316 ( .ip1(n1665), .ip2(PID_haddr_top[11]), .ip3(PID_haddr_top[10]), .op(n1669) );
  inv_1 U2318 ( .ip(PID_haddr_top[2]), .op(n1666) );
  nor2_1 U2322 ( .ip1(PID_haddr_top[2]), .ip2(n1943), .op(n1670) );
  nor3_1 U2325 ( .ip1(PID_haddr_top[23]), .ip2(PID_haddr_top[27]), .ip3(
        PID_haddr_top[26]), .op(n2212) );
  nor3_1 U2326 ( .ip1(PID_haddr_top[24]), .ip2(PID_haddr_top[22]), .ip3(
        PID_haddr_top[17]), .op(n1675) );
  nor2_1 U2336 ( .ip1(PID_haddr_top[7]), .ip2(PID_haddr_top[2]), .op(n1684) );
  nor2_1 U2339 ( .ip1(PID_haddr_top[3]), .ip2(PID_haddr_top[5]), .op(n1686) );
  inv_1 U2342 ( .ip(PID_haddr_top[10]), .op(n1690) );
  nand2_1 U2362 ( .ip1(HREADY_top), .ip2(n3217), .op(n4823) );
  nand2_1 U2474 ( .ip1(HREADY_top), .ip2(n1743), .op(n1769) );
  nand2_1 U2530 ( .ip1(HREADY_top), .ip2(n1788), .op(n2119) );
  nand2_1 U2563 ( .ip1(PID_haddr_top[29]), .ip2(n2118), .op(n1812) );
  nand2_1 U2636 ( .ip1(PID_haddr_top[30]), .ip2(n2118), .op(n1869) );
  nand2_1 U2857 ( .ip1(PID_haddr_top[14]), .ip2(n2118), .op(n2056) );
  nand2_1 U2861 ( .ip1(PID_haddr_top[13]), .ip2(n2118), .op(n2059) );
  nand2_1 U2903 ( .ip1(PID_haddr_top[15]), .ip2(n2118), .op(n2094) );
  nand2_1 U2928 ( .ip1(PID_haddr_top[31]), .ip2(n2118), .op(n2121) );
  nand2_1 U2944 ( .ip1(HREADY_top), .ip2(n2134), .op(n2135) );
  nand2_1 U2949 ( .ip1(n2139), .ip2(HREADY_top), .op(n5814) );
  nand2_1 U2983 ( .ip1(HREADY_top), .ip2(n2167), .op(n5772) );
  inv_1 U3025 ( .ip(PID_hprot_top[3]), .op(n2196) );
  nand2_1 U3027 ( .ip1(HREADY_top), .ip2(n2211), .op(n2197) );
  nand2_1 U3040 ( .ip1(n3276), .ip2(HREADY_top), .op(n2204) );
  or4_1 U3096 ( .ip1(PID_hwdata_top[30]), .ip2(PID_hwdata_top[29]), .ip3(
        PID_hwdata_top[27]), .ip4(PID_hwdata_top[25]), .op(n3231) );
  nand3_1 U3097 ( .ip1(PID_hwdata_top[26]), .ip2(n4704), .ip3(
        PID_hwdata_top[22]), .op(n2270) );
  inv_1 U3102 ( .ip(PID_hwdata_top[18]), .op(n2265) );
  and4_1 U3103 ( .ip1(PID_hwdata_top[19]), .ip2(PID_hwdata_top[24]), .ip3(
        PID_hwdata_top[17]), .ip4(n2265), .op(n2266) );
  nand2_1 U3187 ( .ip1(n3224), .ip2(PID_hwdata_top[25]), .op(n2328) );
  nand2_1 U3353 ( .ip1(n2785), .ip2(PID_hwdata_top[15]), .op(n2460) );
  not_ab_or_c_or_d U3361 ( .ip1(n2792), .ip2(PID_hwdata_top[15]), .ip3(n2464), 
        .ip4(n2463), .op(\CORTEXM0DS_INST/u_logic/Syhvx4 ) );
  nand2_1 U3389 ( .ip1(n3224), .ip2(PID_hwdata_top[27]), .op(n2490) );
  nand2_1 U3391 ( .ip1(n3224), .ip2(PID_hwdata_top[28]), .op(n2492) );
  nand2_1 U3404 ( .ip1(n2785), .ip2(PID_hwdata_top[13]), .op(n2500) );
  and2_1 U3406 ( .ip1(n2792), .ip2(PID_hwdata_top[13]), .op(n2502) );
  not_ab_or_c_or_d U3417 ( .ip1(n2792), .ip2(PID_hwdata_top[8]), .ip3(n2512), 
        .ip4(n2511), .op(\CORTEXM0DS_INST/u_logic/P0ivx4 ) );
  nand2_1 U3418 ( .ip1(n2785), .ip2(PID_hwdata_top[8]), .op(n2513) );
  nand2_1 U3420 ( .ip1(n2785), .ip2(PID_hwdata_top[9]), .op(n2514) );
  and2_1 U3437 ( .ip1(n2792), .ip2(PID_hwdata_top[9]), .op(n2528) );
  and2_1 U3440 ( .ip1(n2792), .ip2(PID_hwdata_top[11]), .op(n2531) );
  nand2_1 U3443 ( .ip1(n2785), .ip2(PID_hwdata_top[11]), .op(n2533) );
  nand2_1 U3452 ( .ip1(n2785), .ip2(PID_hwdata_top[10]), .op(n2541) );
  not_ab_or_c_or_d U3456 ( .ip1(n2792), .ip2(PID_hwdata_top[10]), .ip3(n2544), 
        .ip4(n2543), .op(\CORTEXM0DS_INST/u_logic/B0ivx4 ) );
  nand2_1 U3496 ( .ip1(n2785), .ip2(PID_hwdata_top[7]), .op(n2577) );
  nand2_1 U3544 ( .ip1(n2792), .ip2(PID_hwdata_top[2]), .op(n2620) );
  nand2_1 U3548 ( .ip1(n2785), .ip2(PID_hwdata_top[2]), .op(n2623) );
  nand2_1 U3550 ( .ip1(n2785), .ip2(PID_hwdata_top[3]), .op(n2624) );
  not_ab_or_c_or_d U3554 ( .ip1(n2792), .ip2(PID_hwdata_top[3]), .ip3(n2627), 
        .ip4(n2626), .op(\CORTEXM0DS_INST/u_logic/Y1ivx4 ) );
  nand2_1 U3568 ( .ip1(n2792), .ip2(PID_hwdata_top[4]), .op(n2641) );
  nand2_1 U3572 ( .ip1(n2785), .ip2(PID_hwdata_top[4]), .op(n2644) );
  nand2_1 U3574 ( .ip1(n2785), .ip2(PID_hwdata_top[12]), .op(n2645) );
  not_ab_or_c_or_d U3578 ( .ip1(n2792), .ip2(PID_hwdata_top[12]), .ip3(n2648), 
        .ip4(n2647), .op(\CORTEXM0DS_INST/u_logic/Nzhvx4 ) );
  nand2_1 U3613 ( .ip1(n2792), .ip2(PID_hwdata_top[5]), .op(n2683) );
  nand2_1 U3617 ( .ip1(n2785), .ip2(PID_hwdata_top[5]), .op(n2686) );
  nand2_1 U3641 ( .ip1(n2785), .ip2(PID_hwdata_top[6]), .op(n2711) );
  not_ab_or_c_or_d U3645 ( .ip1(n2792), .ip2(PID_hwdata_top[6]), .ip3(n2714), 
        .ip4(n2713), .op(\CORTEXM0DS_INST/u_logic/D1ivx4 ) );
  nand2_1 U3670 ( .ip1(PID_hwdata_top[14]), .ip2(n2792), .op(n2754) );
  nand2_1 U3674 ( .ip1(n2785), .ip2(PID_hwdata_top[14]), .op(n2757) );
  nand2_1 U3694 ( .ip1(n2785), .ip2(PID_hwdata_top[1]), .op(n2774) );
  nand2_1 U3697 ( .ip1(n2792), .ip2(PID_hwdata_top[1]), .op(n2776) );
  nand2_1 U3705 ( .ip1(n2785), .ip2(PID_hwdata_top[0]), .op(n2786) );
  not_ab_or_c_or_d U3709 ( .ip1(n2792), .ip2(PID_hwdata_top[0]), .ip3(n2791), 
        .ip4(n2790), .op(\CORTEXM0DS_INST/u_logic/T2ivx4 ) );
  nand2_1 U3963 ( .ip1(n12690), .ip2(RAM_hrdata_top[13]), .op(n2974) );
  not_ab_or_c_or_d U3989 ( .ip1(RAM_hrdata_top[7]), .ip2(n12690), .ip3(n2995), 
        .ip4(n2994), .op(n4149) );
  not_ab_or_c_or_d U4010 ( .ip1(n12690), .ip2(RAM_hrdata_top[31]), .ip3(n3009), 
        .ip4(n3008), .op(n4130) );
  not_ab_or_c_or_d U4022 ( .ip1(n12690), .ip2(RAM_hrdata_top[23]), .ip3(n3018), 
        .ip4(n3017), .op(n3020) );
  not_ab_or_c_or_d U4036 ( .ip1(RAM_hrdata_top[15]), .ip2(n12690), .ip3(n3030), 
        .ip4(n4241), .op(n3045) );
  nand2_1 U4078 ( .ip1(n12690), .ip2(RAM_hrdata_top[29]), .op(n3068) );
  not_ab_or_c_or_d U4100 ( .ip1(RAM_hrdata_top[5]), .ip2(n12690), .ip3(n3083), 
        .ip4(n3082), .op(n3085) );
  nand2_1 U4121 ( .ip1(n12690), .ip2(RAM_hrdata_top[21]), .op(n3102) );
  mux2_1 U4147 ( .ip1(n3129), .ip2(PID_hwrite_top), .s(n3128), .op(
        \CORTEXM0DS_INST/u_logic/F4nvx4 ) );
  nand2_1 U4189 ( .ip1(n12690), .ip2(RAM_hrdata_top[9]), .op(n3166) );
  nand2_1 U4221 ( .ip1(n12690), .ip2(RAM_hrdata_top[1]), .op(n3187) );
  nand2_1 U4234 ( .ip1(n12690), .ip2(RAM_hrdata_top[17]), .op(n3197) );
  nand2_1 U4249 ( .ip1(n12690), .ip2(RAM_hrdata_top[25]), .op(n3212) );
  nand2_1 U4354 ( .ip1(HREADY_top), .ip2(n3317), .op(n3348) );
  nand2_1 U4416 ( .ip1(HREADY_top), .ip2(n3369), .op(n3393) );
  nand2_1 U4466 ( .ip1(n12690), .ip2(RAM_hrdata_top[14]), .op(n3420) );
  nand2_1 U4500 ( .ip1(n12690), .ip2(RAM_hrdata_top[30]), .op(n3485) );
  nand2_1 U4534 ( .ip1(n12690), .ip2(RAM_hrdata_top[6]), .op(n3514) );
  nand2_1 U4549 ( .ip1(n12690), .ip2(RAM_hrdata_top[22]), .op(n3554) );
  not_ab_or_c_or_d U4937 ( .ip1(n12690), .ip2(RAM_hrdata_top[8]), .ip3(n3959), 
        .ip4(n3958), .op(n4286) );
  nand2_1 U4946 ( .ip1(n12690), .ip2(RAM_hrdata_top[16]), .op(n3966) );
  and2_1 U4948 ( .ip1(n12690), .ip2(RAM_hrdata_top[24]), .op(n3970) );
  nand2_1 U4955 ( .ip1(n12690), .ip2(RAM_hrdata_top[0]), .op(n3973) );
  nand2_1 U5053 ( .ip1(n12690), .ip2(RAM_hrdata_top[12]), .op(n4087) );
  nand2_1 U5057 ( .ip1(n12690), .ip2(RAM_hrdata_top[28]), .op(n4092) );
  nand2_1 U5066 ( .ip1(n12690), .ip2(RAM_hrdata_top[4]), .op(n4097) );
  nand2_1 U5072 ( .ip1(n12690), .ip2(RAM_hrdata_top[20]), .op(n4106) );
  nand2_1 U5133 ( .ip1(n12690), .ip2(RAM_hrdata_top[27]), .op(n4175) );
  not_ab_or_c_or_d U5136 ( .ip1(n12690), .ip2(RAM_hrdata_top[19]), .ip3(n4180), 
        .ip4(n4241), .op(n4185) );
  nand2_1 U5146 ( .ip1(n12690), .ip2(RAM_hrdata_top[11]), .op(n4190) );
  nand2_1 U5156 ( .ip1(n12690), .ip2(RAM_hrdata_top[3]), .op(n4203) );
  nand2_1 U5170 ( .ip1(n12690), .ip2(RAM_hrdata_top[26]), .op(n4227) );
  nand2_1 U5180 ( .ip1(n12690), .ip2(RAM_hrdata_top[10]), .op(n4237) );
  nand2_1 U5186 ( .ip1(n12690), .ip2(RAM_hrdata_top[18]), .op(n4243) );
  nand2_1 U5197 ( .ip1(n12690), .ip2(RAM_hrdata_top[2]), .op(n4263) );
  nand2_1 U5935 ( .ip1(HREADY_top), .ip2(n4619), .op(n4620) );
  mux2_1 U5991 ( .ip1(PID_hwdata_top[6]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [0]), .s(n4697), .op(
        \CORTEXM0DS_INST/u_logic/Ggmvx4 ) );
  mux2_1 U5992 ( .ip1(PID_hwdata_top[7]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [1]), .s(n4697), .op(
        \CORTEXM0DS_INST/u_logic/Zfmvx4 ) );
  mux2_1 U5993 ( .ip1(PID_hwdata_top[14]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [2]), .s(n4697), .op(
        \CORTEXM0DS_INST/u_logic/Sfmvx4 ) );
  mux2_1 U5994 ( .ip1(PID_hwdata_top[15]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [3]), .s(n4697), .op(
        \CORTEXM0DS_INST/u_logic/Lfmvx4 ) );
  mux2_1 U5995 ( .ip1(PID_hwdata_top[22]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [4]), .s(n4697), .op(
        \CORTEXM0DS_INST/u_logic/Efmvx4 ) );
  mux2_1 U5997 ( .ip1(PID_hwdata_top[30]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [6]), .s(n4697), .op(
        \CORTEXM0DS_INST/u_logic/Qemvx4 ) );
  mux2_1 U6000 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [8]), .ip2(
        PID_hwdata_top[6]), .s(n4699), .op(\CORTEXM0DS_INST/u_logic/Kimvx4 )
         );
  mux2_1 U6001 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [9]), .ip2(
        PID_hwdata_top[7]), .s(n4699), .op(\CORTEXM0DS_INST/u_logic/Dimvx4 )
         );
  mux2_1 U6002 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [10]), .ip2(
        PID_hwdata_top[14]), .s(n4699), .op(\CORTEXM0DS_INST/u_logic/Whmvx4 )
         );
  mux2_1 U6003 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [11]), .ip2(
        PID_hwdata_top[15]), .s(n4699), .op(\CORTEXM0DS_INST/u_logic/Phmvx4 )
         );
  mux2_1 U6004 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [12]), .ip2(
        PID_hwdata_top[22]), .s(n4699), .op(\CORTEXM0DS_INST/u_logic/Ihmvx4 )
         );
  mux2_1 U6006 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [14]), .ip2(
        PID_hwdata_top[30]), .s(n4699), .op(\CORTEXM0DS_INST/u_logic/Ugmvx4 )
         );
  mux2_1 U6009 ( .ip1(PID_hwdata_top[6]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [16]), .s(n4701), .op(
        \CORTEXM0DS_INST/u_logic/Okmvx4 ) );
  mux2_1 U6010 ( .ip1(PID_hwdata_top[7]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [17]), .s(n4701), .op(
        \CORTEXM0DS_INST/u_logic/Hkmvx4 ) );
  mux2_1 U6011 ( .ip1(PID_hwdata_top[14]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [18]), .s(n4701), .op(
        \CORTEXM0DS_INST/u_logic/Akmvx4 ) );
  mux2_1 U6012 ( .ip1(PID_hwdata_top[15]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [19]), .s(n4701), .op(
        \CORTEXM0DS_INST/u_logic/Tjmvx4 ) );
  mux2_1 U6013 ( .ip1(PID_hwdata_top[22]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [20]), .s(n4701), .op(
        \CORTEXM0DS_INST/u_logic/Mjmvx4 ) );
  mux2_1 U6015 ( .ip1(PID_hwdata_top[30]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [22]), .s(n4701), .op(
        \CORTEXM0DS_INST/u_logic/Yimvx4 ) );
  mux2_1 U6018 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [24]), .ip2(
        PID_hwdata_top[6]), .s(n4705), .op(\CORTEXM0DS_INST/u_logic/Smmvx4 )
         );
  mux2_1 U6019 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [25]), .ip2(
        PID_hwdata_top[7]), .s(n4705), .op(\CORTEXM0DS_INST/u_logic/Lmmvx4 )
         );
  mux2_1 U6020 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [26]), .ip2(
        PID_hwdata_top[14]), .s(n4705), .op(\CORTEXM0DS_INST/u_logic/Emmvx4 )
         );
  mux2_1 U6021 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [27]), .ip2(
        PID_hwdata_top[15]), .s(n4705), .op(\CORTEXM0DS_INST/u_logic/Xlmvx4 )
         );
  mux2_1 U6022 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [28]), .ip2(
        PID_hwdata_top[22]), .s(n4705), .op(\CORTEXM0DS_INST/u_logic/Qlmvx4 )
         );
  mux2_1 U6024 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [30]), .ip2(
        PID_hwdata_top[30]), .s(n4705), .op(\CORTEXM0DS_INST/u_logic/Clmvx4 )
         );
  nand3_1 U6117 ( .ip1(n4807), .ip2(RAM_hrdata_top[15]), .ip3(n4806), .op(
        n4808) );
  mux2_1 U6700 ( .ip1(\CORTEXM0DS_INST/u_logic/Ki8vx4 ), .ip2(n5656), .s(
        HREADY_top), .op(\CORTEXM0DS_INST/u_logic/Lrhvx4 ) );
  not_ab_or_c_or_d U6877 ( .ip1(PID_haddr_top[29]), .ip2(n5881), .ip3(
        \CORTEXM0DS_INST/u_logic/Q462z4 ), .ip4(n5880), .op(n5885) );
  and2_1 U6882 ( .ip1(PID_hprot_top[2]), .ip2(n5886), .op(
        \CORTEXM0DS_INST/u_logic/N4422 ) );
  inv_1 U6897 ( .ip(PID_haddr_top[14]), .op(n5906) );
  nand2_1 U6898 ( .ip1(PID_haddr_top[17]), .ip2(n5906), .op(n5907) );
  inv_1 U6900 ( .ip(\PID_htrans_top[1] ), .op(n5908) );
  or4_1 U6901 ( .ip1(n5925), .ip2(RAM_hsel_top), .ip3(n5932), .ip4(n5908), 
        .op(n5921) );
  nand2_1 U6909 ( .ip1(n5913), .ip2(RAM_hready_resp_top), .op(
        \interconnect_ip_inst/n5991 ) );
  nand2_1 U6910 ( .ip1(HREADY_top), .ip2(n5925), .op(n5914) );
  nor2_1 U6911 ( .ip1(PID_haddr_top[13]), .ip2(n5914), .op(n5929) );
  nand2_1 U6912 ( .ip1(n5929), .ip2(\PID_htrans_top[1] ), .op(n5934) );
  nor2_1 U6913 ( .ip1(PID_hwrite_top), .ip2(n5934), .op(n5933) );
  inv_1 U6917 ( .ip(PID_hwrite_top), .op(n5917) );
  nor2_1 U6920 ( .ip1(RAM_hsel_top), .ip2(n5932), .op(n5919) );
  inv_1 U6922 ( .ip(i_ssi_ssi_rst_n_top), .op(\interconnect_ip_inst/n11572 )
         );
  nand3_1 U6927 ( .ip1(HREADY_top), .ip2(PID_haddr_top[13]), .ip3(n5925), .op(
        n5926) );
  or2_1 U6928 ( .ip1(PID_haddr_top[12]), .ip2(n5926), .op(n5928) );
  and2_1 U6934 ( .ip1(PID_hmastlock_top), .ip2(n5932), .op(
        \interconnect_ip_inst/n4860 ) );
  inv_1 U6939 ( .ip(\CORTEXM0DS_INST/u_logic/N4816 ), .op(PID_haddr_top[0]) );
  inv_1 U6940 ( .ip(\CORTEXM0DS_INST/u_logic/Jxovx4 ), .op(PID_haddr_top[10])
         );
  inv_1 U6941 ( .ip(\CORTEXM0DS_INST/u_logic/Cqovx4 ), .op(PID_haddr_top[12])
         );
  inv_1 U6942 ( .ip(\CORTEXM0DS_INST/u_logic/N4767 ), .op(PID_haddr_top[13])
         );
  inv_1 U6943 ( .ip(\CORTEXM0DS_INST/u_logic/N4751 ), .op(PID_haddr_top[14])
         );
  inv_1 U6944 ( .ip(\CORTEXM0DS_INST/u_logic/Vpovx4 ), .op(PID_haddr_top[16])
         );
  inv_1 U6945 ( .ip(\CORTEXM0DS_INST/u_logic/Bv0wx4 ), .op(PID_haddr_top[17])
         );
  inv_1 U6946 ( .ip(\CORTEXM0DS_INST/u_logic/Fq0wx4 ), .op(PID_haddr_top[18])
         );
  inv_1 U6947 ( .ip(\CORTEXM0DS_INST/u_logic/Ql0wx4 ), .op(PID_haddr_top[19])
         );
  inv_1 U6948 ( .ip(\CORTEXM0DS_INST/u_logic/N4674 ), .op(PID_haddr_top[1]) );
  inv_1 U6949 ( .ip(\CORTEXM0DS_INST/u_logic/Ug0wx4 ), .op(PID_haddr_top[20])
         );
  inv_1 U6950 ( .ip(\CORTEXM0DS_INST/u_logic/Fc0wx4 ), .op(PID_haddr_top[21])
         );
  inv_1 U6951 ( .ip(\CORTEXM0DS_INST/u_logic/C70wx4 ), .op(PID_haddr_top[22])
         );
  inv_1 U6952 ( .ip(\CORTEXM0DS_INST/u_logic/Y92wx4 ), .op(PID_haddr_top[23])
         );
  inv_1 U6953 ( .ip(\CORTEXM0DS_INST/u_logic/Y1pvx4 ), .op(PID_haddr_top[24])
         );
  inv_1 U6954 ( .ip(\CORTEXM0DS_INST/u_logic/Rnovx4 ), .op(PID_haddr_top[25])
         );
  inv_1 U6955 ( .ip(\CORTEXM0DS_INST/u_logic/Nhzvx4 ), .op(PID_haddr_top[26])
         );
  inv_1 U6956 ( .ip(\CORTEXM0DS_INST/u_logic/Vezvx4 ), .op(PID_haddr_top[27])
         );
  inv_1 U6957 ( .ip(\CORTEXM0DS_INST/u_logic/V2qvx4 ), .op(PID_haddr_top[28])
         );
  inv_1 U6958 ( .ip(\CORTEXM0DS_INST/u_logic/N4518 ), .op(PID_haddr_top[31])
         );
  inv_1 U6959 ( .ip(\CORTEXM0DS_INST/u_logic/Yuovx4 ), .op(PID_haddr_top[4])
         );
  inv_1 U6960 ( .ip(\CORTEXM0DS_INST/u_logic/Rxzvx4 ), .op(PID_haddr_top[5])
         );
  inv_1 U6961 ( .ip(\CORTEXM0DS_INST/u_logic/Hszvx4 ), .op(PID_haddr_top[6])
         );
  inv_1 U6962 ( .ip(\CORTEXM0DS_INST/u_logic/S4qvx4 ), .op(PID_haddr_top[7])
         );
  inv_1 U6963 ( .ip(\CORTEXM0DS_INST/u_logic/N4439 ), .op(PID_haddr_top[30])
         );
  or2_1 U6964 ( .ip1(\CORTEXM0DS_INST/u_logic/E562z4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Q462z4 ), .op(PID_haddr_top[29]) );
  or2_1 U6965 ( .ip1(PID_haddr_top[30]), .ip2(PID_haddr_top[29]), .op(
        PID_hprot_top[2]) );
  inv_1 U6966 ( .ip(\CORTEXM0DS_INST/u_logic/N4422 ), .op(PID_hprot_top[3]) );
  and2_1 U6967 ( .ip1(\CORTEXM0DS_INST/u_logic/A362z4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Oq42z4 ), .op(PID_hsize_top[0]) );
  inv_1 U6968 ( .ip(\CORTEXM0DS_INST/u_logic/N4421 ), .op(PID_hsize_top[1]) );
  inv_1 U6969 ( .ip(\CORTEXM0DS_INST/u_logic/N4396 ), .op(PID_hprot_top[0]) );
  and2_1 U6970 ( .ip1(n6110), .ip2(\CORTEXM0DS_INST/u_logic/Xmywx4 ), .op(
        \PID_htrans_top[1] ) );
  inv_1 U6971 ( .ip(\CORTEXM0DS_INST/u_logic/N4359 ), .op(PID_hwdata_top[0])
         );
  inv_1 U6972 ( .ip(\CORTEXM0DS_INST/u_logic/N4282 ), .op(PID_hwdata_top[24])
         );
  inv_1 U6973 ( .ip(\CORTEXM0DS_INST/u_logic/N4227 ), .op(PID_hwdata_top[25])
         );
  inv_1 U6974 ( .ip(\CORTEXM0DS_INST/u_logic/N4170 ), .op(PID_hwdata_top[26])
         );
  inv_1 U6975 ( .ip(\CORTEXM0DS_INST/u_logic/N4116 ), .op(PID_hwdata_top[27])
         );
  inv_1 U6976 ( .ip(\CORTEXM0DS_INST/u_logic/Sx3wx4 ), .op(PID_hwdata_top[28])
         );
  inv_1 U6977 ( .ip(\CORTEXM0DS_INST/u_logic/N4005 ), .op(PID_hwdata_top[29])
         );
  inv_1 U6978 ( .ip(\CORTEXM0DS_INST/u_logic/N3967 ), .op(PID_hwdata_top[31])
         );
  inv_1 U6979 ( .ip(\CORTEXM0DS_INST/u_logic/N3966 ), .op(PID_hwdata_top[3])
         );
  inv_1 U6980 ( .ip(n6170), .op(PID_hwdata_top[4]) );
  inv_1 U6981 ( .ip(n6175), .op(PID_hwdata_top[5]) );
  inv_1 U6982 ( .ip(\CORTEXM0DS_INST/u_logic/N3946 ), .op(PID_hwdata_top[6])
         );
  inv_1 U6983 ( .ip(n6161), .op(PID_hwdata_top[7]) );
  inv_1 U6984 ( .ip(n6166), .op(PID_hwdata_top[2]) );
  inv_1 U6985 ( .ip(\CORTEXM0DS_INST/u_logic/N3783 ), .op(PID_hwdata_top[30])
         );
  inv_1 U6986 ( .ip(\CORTEXM0DS_INST/u_logic/N2678 ), .op(PID_hwrite_top) );
  inv_1 U6987 ( .ip(\CORTEXM0DS_INST/u_logic/Bq5wx4 ), .op(PID_hwdata_top[14])
         );
  inv_1 U6988 ( .ip(n6184), .op(PID_hwdata_top[1]) );
  inv_1 U6989 ( .ip(\CORTEXM0DS_INST/u_logic/O24wx4 ), .op(PID_hwdata_top[16])
         );
  inv_1 U6990 ( .ip(\CORTEXM0DS_INST/u_logic/N1447 ), .op(PID_haddr_top[15])
         );
  inv_1 U6991 ( .ip(\CORTEXM0DS_INST/u_logic/Xxovx4 ), .op(PID_haddr_top[9])
         );
  inv_1 U6992 ( .ip(\CORTEXM0DS_INST/u_logic/Ekovx4 ), .op(PID_haddr_top[3])
         );
  inv_1 U6993 ( .ip(\CORTEXM0DS_INST/u_logic/Owovx4 ), .op(PID_haddr_top[11])
         );
  inv_1 U6994 ( .ip(\CORTEXM0DS_INST/u_logic/Z6ovx4 ), .op(PID_haddr_top[8])
         );
  inv_1 U6995 ( .ip(\CORTEXM0DS_INST/u_logic/Fvovx4 ), .op(PID_haddr_top[2])
         );
  nand2_1 U6996 ( .ip1(n5972), .ip2(n5971), .op(PID_hwdata_top[23]) );
  nand2_1 U6997 ( .ip1(n5974), .ip2(n5973), .op(PID_hwdata_top[22]) );
  nand2_1 U6998 ( .ip1(n5976), .ip2(n5975), .op(PID_hwdata_top[21]) );
  nand2_1 U6999 ( .ip1(n5978), .ip2(n5977), .op(PID_hwdata_top[19]) );
  nand2_1 U7000 ( .ip1(n5980), .ip2(n5979), .op(PID_hwdata_top[20]) );
  nand2_1 U7001 ( .ip1(n5982), .ip2(n5981), .op(PID_hwdata_top[17]) );
  nand2_1 U7002 ( .ip1(n5984), .ip2(n5983), .op(PID_hwdata_top[18]) );
  nand2_1 U7003 ( .ip1(n5986), .ip2(n5985), .op(PID_hwdata_top[15]) );
  nand2_1 U7004 ( .ip1(n5988), .ip2(n5987), .op(PID_hwdata_top[13]) );
  nand2_1 U7005 ( .ip1(n5990), .ip2(n5989), .op(PID_hwdata_top[12]) );
  nand2_1 U7006 ( .ip1(n5992), .ip2(n5991), .op(PID_hwdata_top[11]) );
  nand2_1 U7007 ( .ip1(n5994), .ip2(n5993), .op(PID_hwdata_top[10]) );
  nand2_1 U7008 ( .ip1(n5996), .ip2(n5995), .op(PID_hwdata_top[9]) );
  nand2_1 U7009 ( .ip1(n5998), .ip2(n5997), .op(PID_hwdata_top[8]) );
  nand4_1 U7010 ( .ip1(n6693), .ip2(n6692), .ip3(n6691), .ip4(n6690), .op(
        n6694) );
  nand4_1 U7011 ( .ip1(n6547), .ip2(n6546), .ip3(n6545), .ip4(n6544), .op(
        n6548) );
  nand4_1 U7012 ( .ip1(n6711), .ip2(n6710), .ip3(n6709), .ip4(n6708), .op(
        n6712) );
  nand4_1 U7013 ( .ip1(n6529), .ip2(n6528), .ip3(n6527), .ip4(n6526), .op(
        n6530) );
  nand4_1 U7014 ( .ip1(n6721), .ip2(n6720), .ip3(n6719), .ip4(n6718), .op(
        n6722) );
  nor4_1 U7015 ( .ip1(n11797), .ip2(n7016), .ip3(n7015), .ip4(n7014), .op(
        n7524) );
  nor4_1 U7016 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n8424), .ip3(
        n10698), .ip4(n11682), .op(n7016) );
  nor4_1 U7017 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip3(n12623), .ip4(n11682), .op(
        n7014) );
  nand4_1 U7018 ( .ip1(n6678), .ip2(n6677), .ip3(n6676), .ip4(n6675), .op(
        n6679) );
  nand4_1 U7019 ( .ip1(n6768), .ip2(n6767), .ip3(n6766), .ip4(n6765), .op(
        n6769) );
  nand4_1 U7020 ( .ip1(n6515), .ip2(n6514), .ip3(n6513), .ip4(n6512), .op(
        n6516) );
  nor4_1 U7021 ( .ip1(n6810), .ip2(n6809), .ip3(n6808), .ip4(n6807), .op(n7106) );
  nand4_1 U7022 ( .ip1(n6611), .ip2(n6610), .ip3(n6609), .ip4(n6608), .op(
        n6612) );
  nand4_1 U7023 ( .ip1(n6568), .ip2(n6567), .ip3(n6566), .ip4(n6565), .op(
        n6569) );
  nand4_1 U7024 ( .ip1(n6595), .ip2(n6594), .ip3(n6593), .ip4(n6592), .op(
        n6596) );
  nand4_1 U7025 ( .ip1(n6735), .ip2(n6734), .ip3(n6733), .ip4(n6732), .op(
        n6736) );
  nand4_1 U7026 ( .ip1(n6629), .ip2(n6628), .ip3(n6627), .ip4(n6626), .op(
        n6630) );
  nand4_1 U7027 ( .ip1(n6620), .ip2(n6619), .ip3(n6618), .ip4(n6617), .op(
        n6621) );
  nand4_1 U7028 ( .ip1(n6638), .ip2(n6637), .ip3(n6636), .ip4(n6635), .op(
        n6639) );
  nand4_1 U7029 ( .ip1(n6651), .ip2(n6650), .ip3(n6649), .ip4(n6648), .op(
        n6652) );
  nand4_1 U7030 ( .ip1(n6488), .ip2(n6487), .ip3(n6486), .ip4(n6485), .op(
        n6489) );
  nand4_1 U7031 ( .ip1(n6817), .ip2(n6816), .ip3(n6815), .ip4(n6814), .op(
        n6818) );
  nand4_1 U7032 ( .ip1(n6702), .ip2(n6701), .ip3(n6700), .ip4(n6699), .op(
        n6703) );
  nand4_1 U7033 ( .ip1(n6873), .ip2(n6872), .ip3(n6871), .ip4(n6870), .op(
        n6877) );
  nand4_1 U7034 ( .ip1(n6391), .ip2(n6390), .ip3(n6389), .ip4(n6388), .op(
        n6392) );
  nor4_1 U7035 ( .ip1(n7021), .ip2(n7020), .ip3(n7019), .ip4(n7018), .op(n7022) );
  nor4_1 U7036 ( .ip1(n9740), .ip2(n6838), .ip3(n6837), .ip4(n6836), .op(n6839) );
  nand4_1 U7037 ( .ip1(n6452), .ip2(n6451), .ip3(n6450), .ip4(n6449), .op(
        n6453) );
  nand4_1 U7038 ( .ip1(n6447), .ip2(n6446), .ip3(n6445), .ip4(n6444), .op(
        n6454) );
  nand4_1 U7039 ( .ip1(n6915), .ip2(n6914), .ip3(n6913), .ip4(n6912), .op(
        n6916) );
  nand4_1 U7040 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip3(n12609), .ip4(n9807), .op(
        n6856) );
  nand4_1 U7041 ( .ip1(n6998), .ip2(n6997), .ip3(n6996), .ip4(n6995), .op(
        n6999) );
  nand4_1 U7042 ( .ip1(n7036), .ip2(n7035), .ip3(n7034), .ip4(n7033), .op(
        n7037) );
  nand4_1 U7043 ( .ip1(n7459), .ip2(n7458), .ip3(n7457), .ip4(n7456), .op(
        n7460) );
  nand4_1 U7044 ( .ip1(n7486), .ip2(n7485), .ip3(n7484), .ip4(n7483), .op(
        n7487) );
  nand4_1 U7045 ( .ip1(n7510), .ip2(n7509), .ip3(n7508), .ip4(n7507), .op(
        n7511) );
  nand4_1 U7046 ( .ip1(n7537), .ip2(n7536), .ip3(n7535), .ip4(n7534), .op(
        n7538) );
  nor4_1 U7047 ( .ip1(n10555), .ip2(n11794), .ip3(n6300), .ip4(n6299), .op(
        n6306) );
  nand4_1 U7048 ( .ip1(n6886), .ip2(n6885), .ip3(n6884), .ip4(n6883), .op(
        n6887) );
  nand4_1 U7049 ( .ip1(n7427), .ip2(n7426), .ip3(n7425), .ip4(n7424), .op(
        n7428) );
  nand4_1 U7050 ( .ip1(n7414), .ip2(n7413), .ip3(n7412), .ip4(n7411), .op(
        n7415) );
  nand4_1 U7051 ( .ip1(n7389), .ip2(n7388), .ip3(n7387), .ip4(n7386), .op(
        n7390) );
  nand4_1 U7052 ( .ip1(n7367), .ip2(n7366), .ip3(n7365), .ip4(n7364), .op(
        n7368) );
  nand4_1 U7053 ( .ip1(n7341), .ip2(n7340), .ip3(n7339), .ip4(n7338), .op(
        n7342) );
  nand4_1 U7054 ( .ip1(n7292), .ip2(n7291), .ip3(n7290), .ip4(n7289), .op(
        n7293) );
  nand4_1 U7055 ( .ip1(n7280), .ip2(n7279), .ip3(n7278), .ip4(n7277), .op(
        n7281) );
  nand4_1 U7056 ( .ip1(n7244), .ip2(n7243), .ip3(n7242), .ip4(n7241), .op(
        n7245) );
  nand4_1 U7057 ( .ip1(n7222), .ip2(n7221), .ip3(n7220), .ip4(n7219), .op(
        n7223) );
  nand4_1 U7058 ( .ip1(n7198), .ip2(n7197), .ip3(n7196), .ip4(n7195), .op(
        n7199) );
  nand4_1 U7059 ( .ip1(n7152), .ip2(n7151), .ip3(n7150), .ip4(n7149), .op(
        n7153) );
  nand4_1 U7060 ( .ip1(n7095), .ip2(n7094), .ip3(n7093), .ip4(n7092), .op(
        n7096) );
  nand4_1 U7061 ( .ip1(n8570), .ip2(n8569), .ip3(n8568), .ip4(n8567), .op(
        n8571) );
  nand4_1 U7062 ( .ip1(n6731), .ip2(n6730), .ip3(n6729), .ip4(n6728), .op(
        n6781) );
  nand4_1 U7063 ( .ip1(n6647), .ip2(n6646), .ip3(n6645), .ip4(n6644), .op(
        n6689) );
  nand4_1 U7064 ( .ip1(n7528), .ip2(n7527), .ip3(n7526), .ip4(n7525), .op(
        n7529) );
  nor4_1 U7065 ( .ip1(n11228), .ip2(n10945), .ip3(n8494), .ip4(n10865), .op(
        n11797) );
  nand4_1 U7066 ( .ip1(n7555), .ip2(n7554), .ip3(n7553), .ip4(n7552), .op(
        n7556) );
  nand4_1 U7067 ( .ip1(n7609), .ip2(n7608), .ip3(n7607), .ip4(n7606), .op(
        n7610) );
  nand4_1 U7068 ( .ip1(n7580), .ip2(n7579), .ip3(n7578), .ip4(n7577), .op(
        n7581) );
  nand4_1 U7069 ( .ip1(n7028), .ip2(n7027), .ip3(n7026), .ip4(n7025), .op(
        n7029) );
  nand4_1 U7070 ( .ip1(n7053), .ip2(n7052), .ip3(n7051), .ip4(n7050), .op(
        n7054) );
  nand4_1 U7071 ( .ip1(n7232), .ip2(n7231), .ip3(n7230), .ip4(n7229), .op(
        n7233) );
  nand4_1 U7072 ( .ip1(n7476), .ip2(n7475), .ip3(n7474), .ip4(n7473), .op(
        n7477) );
  nand4_1 U7073 ( .ip1(n7503), .ip2(n7502), .ip3(n7501), .ip4(n7500), .op(
        n7504) );
  nand4_1 U7074 ( .ip1(n6335), .ip2(n6334), .ip3(n6435), .ip4(n10810), .op(
        n6336) );
  nand4_1 U7075 ( .ip1(n11693), .ip2(n11692), .ip3(n10698), .ip4(n11793), .op(
        n6321) );
  nand4_1 U7076 ( .ip1(n7978), .ip2(n7977), .ip3(n7976), .ip4(n7975), .op(
        n7983) );
  nand4_1 U7077 ( .ip1(n6374), .ip2(n6373), .ip3(n6372), .ip4(n6371), .op(
        n8934) );
  nand4_1 U7078 ( .ip1(n7763), .ip2(n7762), .ip3(n7761), .ip4(n7760), .op(
        n7764) );
  nand4_1 U7079 ( .ip1(n7759), .ip2(n7758), .ip3(n7757), .ip4(n7756), .op(
        n7765) );
  nand4_1 U7080 ( .ip1(n7830), .ip2(n7829), .ip3(n7828), .ip4(n7827), .op(
        n7831) );
  nand4_1 U7081 ( .ip1(n7826), .ip2(n7825), .ip3(n7824), .ip4(n7823), .op(
        n7832) );
  nand4_1 U7082 ( .ip1(n7877), .ip2(n7876), .ip3(n7875), .ip4(n7874), .op(
        n7878) );
  nand4_1 U7083 ( .ip1(n7873), .ip2(n7872), .ip3(n7871), .ip4(n7870), .op(
        n7879) );
  nand4_1 U7084 ( .ip1(n7621), .ip2(n7620), .ip3(n7619), .ip4(n7618), .op(
        n7622) );
  nand4_1 U7085 ( .ip1(n7617), .ip2(n7616), .ip3(n7615), .ip4(n7614), .op(
        n7623) );
  nand4_1 U7086 ( .ip1(n7117), .ip2(n7116), .ip3(n7115), .ip4(n7114), .op(
        n7118) );
  nand4_1 U7087 ( .ip1(n7113), .ip2(n7112), .ip3(n7111), .ip4(n7110), .op(
        n7119) );
  nand4_1 U7088 ( .ip1(n7671), .ip2(n7670), .ip3(n7669), .ip4(n7668), .op(
        n7672) );
  nand4_1 U7089 ( .ip1(n7667), .ip2(n7666), .ip3(n7665), .ip4(n7664), .op(
        n7673) );
  nand4_1 U7090 ( .ip1(n8550), .ip2(n8549), .ip3(n8548), .ip4(n8547), .op(
        n8555) );
  nand4_1 U7091 ( .ip1(n7716), .ip2(n7715), .ip3(n7714), .ip4(n7713), .op(
        n7717) );
  nand4_1 U7092 ( .ip1(n7712), .ip2(n7711), .ip3(n7710), .ip4(n7709), .op(
        n7718) );
  nand4_1 U7093 ( .ip1(n7738), .ip2(n7737), .ip3(n7736), .ip4(n7735), .op(
        n7739) );
  nand4_1 U7094 ( .ip1(n7734), .ip2(n7733), .ip3(n7732), .ip4(n7731), .op(
        n7740) );
  nand4_1 U7095 ( .ip1(n6307), .ip2(n6306), .ip3(n6305), .ip4(n6414), .op(
        n6308) );
  nand4_1 U7096 ( .ip1(n6960), .ip2(n6959), .ip3(n6958), .ip4(n6957), .op(
        n6961) );
  nand4_1 U7097 ( .ip1(n7442), .ip2(n7441), .ip3(n7440), .ip4(n7439), .op(
        n7443) );
  nand4_1 U7098 ( .ip1(n7433), .ip2(n7432), .ip3(n7431), .ip4(n7430), .op(
        n7434) );
  nand4_1 U7099 ( .ip1(n7420), .ip2(n7419), .ip3(n7418), .ip4(n7417), .op(
        n7421) );
  nand4_1 U7100 ( .ip1(n7404), .ip2(n7403), .ip3(n7402), .ip4(n7401), .op(
        n7405) );
  nand4_1 U7101 ( .ip1(n7395), .ip2(n7394), .ip3(n7393), .ip4(n7392), .op(
        n7396) );
  nand4_1 U7102 ( .ip1(n7377), .ip2(n7376), .ip3(n7375), .ip4(n7374), .op(
        n7378) );
  nand4_1 U7103 ( .ip1(n7373), .ip2(n7372), .ip3(n7371), .ip4(n7370), .op(
        n9498) );
  nand4_1 U7104 ( .ip1(n7355), .ip2(n7354), .ip3(n7353), .ip4(n7352), .op(
        n7356) );
  nand4_1 U7105 ( .ip1(n7347), .ip2(n7346), .ip3(n7345), .ip4(n7344), .op(
        n7348) );
  nand4_1 U7106 ( .ip1(n7329), .ip2(n7328), .ip3(n7327), .ip4(n7326), .op(
        n7330) );
  nand4_1 U7107 ( .ip1(n7304), .ip2(n7303), .ip3(n7302), .ip4(n7301), .op(
        n7305) );
  nand4_1 U7108 ( .ip1(n7298), .ip2(n7297), .ip3(n7296), .ip4(n7295), .op(
        n7299) );
  nand4_1 U7109 ( .ip1(n7286), .ip2(n7285), .ip3(n7284), .ip4(n7283), .op(
        n7287) );
  nand4_1 U7110 ( .ip1(n7270), .ip2(n7269), .ip3(n7268), .ip4(n7267), .op(
        n7271) );
  nand4_1 U7111 ( .ip1(n7256), .ip2(n7255), .ip3(n7254), .ip4(n7253), .op(
        n7257) );
  nand4_1 U7112 ( .ip1(n7250), .ip2(n7249), .ip3(n7248), .ip4(n7247), .op(
        n7251) );
  nand4_1 U7113 ( .ip1(n7228), .ip2(n7227), .ip3(n7226), .ip4(n7225), .op(
        n9598) );
  nand4_1 U7114 ( .ip1(n7208), .ip2(n7207), .ip3(n7206), .ip4(n7205), .op(
        n7209) );
  nand4_1 U7115 ( .ip1(n7204), .ip2(n7203), .ip3(n7202), .ip4(n7201), .op(
        n9624) );
  nand4_1 U7116 ( .ip1(n7164), .ip2(n7163), .ip3(n7162), .ip4(n7161), .op(
        n7165) );
  nand4_1 U7117 ( .ip1(n7158), .ip2(n7157), .ip3(n7156), .ip4(n7155), .op(
        n7159) );
  nand4_1 U7118 ( .ip1(n7101), .ip2(n7100), .ip3(n7099), .ip4(n7098), .op(
        n7102) );
  nand4_1 U7119 ( .ip1(n7085), .ip2(n7084), .ip3(n7083), .ip4(n7082), .op(
        n7086) );
  nand4_1 U7120 ( .ip1(n8576), .ip2(n8575), .ip3(n8574), .ip4(n8573), .op(
        n9524) );
  nand4_1 U7121 ( .ip1(n9294), .ip2(n9293), .ip3(n9292), .ip4(n9291), .op(
        n9295) );
  nand4_1 U7122 ( .ip1(n9360), .ip2(n9359), .ip3(n9358), .ip4(n9357), .op(
        n9361) );
  nor4_1 U7123 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n12623), .ip3(
        n5639), .ip4(n11693), .op(n6419) );
  nor4_1 U7124 ( .ip1(n6402), .ip2(n11884), .ip3(n11892), .ip4(n12049), .op(
        n8937) );
  nand4_1 U7125 ( .ip1(n7238), .ip2(n7237), .ip3(n7236), .ip4(n7235), .op(
        n7239) );
  nand4_1 U7126 ( .ip1(n6977), .ip2(n6976), .ip3(n6975), .ip4(n6974), .op(
        n6978) );
  nand4_1 U7127 ( .ip1(n6340), .ip2(n6339), .ip3(n6338), .ip4(n6337), .op(
        n2139) );
  nand4_1 U7128 ( .ip1(n7987), .ip2(n7986), .ip3(n7985), .ip4(n7984), .op(
        n7988) );
  nor4_1 U7129 ( .ip1(n11796), .ip2(n12117), .ip3(n12623), .ip4(n11223), .op(
        n10556) );
  nand4_1 U7130 ( .ip1(n6831), .ip2(n6830), .ip3(n6829), .ip4(n6828), .op(
        n6832) );
  nand4_1 U7131 ( .ip1(n7769), .ip2(n7768), .ip3(n7767), .ip4(n7766), .op(
        n7770) );
  nand4_1 U7132 ( .ip1(n7784), .ip2(n7783), .ip3(n7782), .ip4(n7781), .op(
        n7785) );
  nand4_1 U7133 ( .ip1(n7780), .ip2(n7779), .ip3(n7778), .ip4(n7777), .op(
        n7786) );
  nand4_1 U7134 ( .ip1(n7806), .ip2(n7805), .ip3(n7804), .ip4(n7803), .op(
        n7811) );
  nand4_1 U7135 ( .ip1(n7849), .ip2(n7848), .ip3(n7847), .ip4(n7846), .op(
        n7855) );
  nand4_1 U7136 ( .ip1(n7853), .ip2(n7852), .ip3(n7851), .ip4(n7850), .op(
        n7854) );
  nand4_1 U7137 ( .ip1(n7904), .ip2(n7903), .ip3(n7902), .ip4(n7901), .op(
        n7905) );
  nand4_1 U7138 ( .ip1(n7900), .ip2(n7899), .ip3(n7898), .ip4(n7897), .op(
        n7906) );
  nand4_1 U7139 ( .ip1(n7923), .ip2(n7922), .ip3(n7921), .ip4(n7920), .op(
        n7929) );
  nand4_1 U7140 ( .ip1(n7927), .ip2(n7926), .ip3(n7925), .ip4(n7924), .op(
        n7928) );
  nand4_1 U7141 ( .ip1(n7952), .ip2(n7951), .ip3(n7950), .ip4(n7949), .op(
        n7953) );
  nand4_1 U7142 ( .ip1(n7948), .ip2(n7947), .ip3(n7946), .ip4(n7945), .op(
        n7954) );
  nand4_1 U7143 ( .ip1(n7566), .ip2(n7565), .ip3(n7564), .ip4(n7563), .op(
        n7572) );
  nand4_1 U7144 ( .ip1(n7570), .ip2(n7569), .ip3(n7568), .ip4(n7567), .op(
        n7571) );
  nand4_1 U7145 ( .ip1(n7179), .ip2(n7178), .ip3(n7177), .ip4(n7176), .op(
        n7185) );
  nand4_1 U7146 ( .ip1(n7183), .ip2(n7182), .ip3(n7181), .ip4(n7180), .op(
        n7184) );
  nand4_1 U7147 ( .ip1(n7595), .ip2(n7594), .ip3(n7593), .ip4(n7592), .op(
        n7601) );
  nand4_1 U7148 ( .ip1(n7599), .ip2(n7598), .ip3(n7597), .ip4(n7596), .op(
        n7600) );
  nand4_1 U7149 ( .ip1(n7137), .ip2(n7136), .ip3(n7135), .ip4(n7134), .op(
        n7142) );
  nand4_1 U7150 ( .ip1(n7646), .ip2(n7645), .ip3(n7644), .ip4(n7643), .op(
        n7647) );
  nand4_1 U7151 ( .ip1(n7642), .ip2(n7641), .ip3(n7640), .ip4(n7639), .op(
        n7648) );
  nand4_1 U7152 ( .ip1(n7677), .ip2(n7676), .ip3(n7675), .ip4(n7674), .op(
        n7678) );
  nand4_1 U7153 ( .ip1(n7692), .ip2(n7691), .ip3(n7690), .ip4(n7689), .op(
        n7693) );
  nand4_1 U7154 ( .ip1(n7688), .ip2(n7687), .ip3(n7686), .ip4(n7685), .op(
        n7694) );
  nand4_1 U7155 ( .ip1(n8559), .ip2(n8558), .ip3(n8557), .ip4(n8556), .op(
        n8560) );
  nand4_1 U7156 ( .ip1(n9276), .ip2(n9275), .ip3(n9274), .ip4(n9273), .op(
        n9277) );
  nand4_1 U7157 ( .ip1(n9272), .ip2(n9271), .ip3(n9270), .ip4(n9269), .op(
        n9278) );
  nand4_1 U7158 ( .ip1(n9330), .ip2(n9329), .ip3(n9328), .ip4(n9327), .op(
        n9331) );
  nand4_1 U7159 ( .ip1(n9322), .ip2(n9321), .ip3(n9320), .ip4(n9319), .op(
        n9332) );
  nand4_1 U7160 ( .ip1(n6945), .ip2(n12606), .ip3(n11242), .ip4(n12343), .op(
        n2208) );
  nand4_1 U7161 ( .ip1(n6907), .ip2(n6906), .ip3(n6905), .ip4(n6904), .op(
        n6908) );
  nand4_1 U7162 ( .ip1(n6967), .ip2(n6966), .ip3(n6965), .ip4(n6964), .op(
        n6968) );
  nand4_1 U7163 ( .ip1(n7448), .ip2(n7447), .ip3(n7446), .ip4(n7445), .op(
        n7449) );
  nand4_1 U7164 ( .ip1(n7383), .ip2(n7382), .ip3(n7381), .ip4(n7380), .op(
        n7384) );
  nand4_1 U7165 ( .ip1(n7361), .ip2(n7360), .ip3(n7359), .ip4(n7358), .op(
        n12191) );
  nand4_1 U7166 ( .ip1(n7335), .ip2(n7334), .ip3(n7333), .ip4(n7332), .op(
        n7336) );
  nand4_1 U7167 ( .ip1(n7318), .ip2(n7317), .ip3(n7316), .ip4(n7315), .op(
        n7319) );
  nand4_1 U7168 ( .ip1(n7310), .ip2(n7309), .ip3(n7308), .ip4(n7307), .op(
        n7311) );
  nor4_1 U7169 ( .ip1(n10193), .ip2(n10197), .ip3(n10329), .ip4(n8064), .op(
        n8533) );
  nand4_1 U7170 ( .ip1(n7276), .ip2(n7275), .ip3(n7274), .ip4(n7273), .op(
        n12235) );
  nand4_1 U7171 ( .ip1(n7262), .ip2(n7261), .ip3(n7260), .ip4(n7259), .op(
        n7263) );
  nand4_1 U7172 ( .ip1(n7214), .ip2(n7213), .ip3(n7212), .ip4(n7211), .op(
        n7215) );
  nand4_1 U7173 ( .ip1(n7170), .ip2(n7169), .ip3(n7168), .ip4(n7167), .op(
        n7171) );
  nand4_1 U7174 ( .ip1(n7091), .ip2(n7090), .ip3(n7089), .ip4(n7088), .op(
        n9513) );
  nand4_1 U7175 ( .ip1(n9300), .ip2(n9299), .ip3(n9298), .ip4(n9297), .op(
        n9471) );
  nand4_1 U7176 ( .ip1(n9370), .ip2(n9369), .ip3(n9368), .ip4(n9367), .op(
        n9990) );
  nand4_1 U7177 ( .ip1(n6983), .ip2(n6982), .ip3(n6981), .ip4(n6980), .op(
        n6984) );
  nand4_1 U7178 ( .ip1(n6925), .ip2(n6924), .ip3(n6923), .ip4(n6922), .op(
        n6926) );
  nand4_1 U7179 ( .ip1(n6212), .ip2(n12079), .ip3(n10224), .ip4(n10204), .op(
        n10955) );
  nor4_1 U7180 ( .ip1(n12108), .ip2(n12397), .ip3(n12381), .ip4(n12370), .op(
        n6212) );
  nand4_1 U7181 ( .ip1(n7012), .ip2(n7011), .ip3(n7010), .ip4(n7009), .op(
        n12671) );
  nand4_1 U7182 ( .ip1(n7815), .ip2(n7814), .ip3(n7813), .ip4(n7812), .op(
        n7816) );
  nand4_1 U7183 ( .ip1(n7049), .ip2(n7048), .ip3(n7047), .ip4(n7046), .op(
        n12677) );
  nand4_1 U7184 ( .ip1(n7472), .ip2(n7471), .ip3(n7470), .ip4(n7469), .op(
        n12675) );
  nand4_1 U7185 ( .ip1(n7499), .ip2(n7498), .ip3(n7497), .ip4(n7496), .op(
        n12679) );
  nand4_1 U7186 ( .ip1(n7910), .ip2(n7909), .ip3(n7908), .ip4(n7907), .op(
        n12680) );
  nand4_1 U7187 ( .ip1(n7523), .ip2(n7522), .ip3(n7521), .ip4(n7520), .op(
        n12681) );
  nand4_1 U7188 ( .ip1(n7933), .ip2(n7932), .ip3(n7931), .ip4(n7930), .op(
        n12682) );
  nand4_1 U7189 ( .ip1(n7550), .ip2(n7549), .ip3(n7548), .ip4(n7547), .op(
        n12685) );
  nand4_1 U7190 ( .ip1(n7576), .ip2(n7575), .ip3(n7574), .ip4(n7573), .op(
        n12661) );
  nand4_1 U7191 ( .ip1(n7605), .ip2(n7604), .ip3(n7603), .ip4(n7602), .op(
        n12662) );
  nand4_1 U7192 ( .ip1(n7146), .ip2(n7145), .ip3(n7144), .ip4(n7143), .op(
        n7147) );
  nand4_1 U7193 ( .ip1(n7324), .ip2(n7323), .ip3(n7322), .ip4(n7321), .op(
        n10027) );
  nand4_1 U7194 ( .ip1(n6892), .ip2(n9379), .ip3(n10971), .ip4(n6891), .op(
        n6893) );
  nand4_1 U7195 ( .ip1(n6440), .ip2(n6439), .ip3(n6438), .ip4(n6437), .op(
        n12343) );
  nor4_1 U7196 ( .ip1(n6434), .ip2(n10555), .ip3(n6433), .ip4(n10052), .op(
        n6439) );
  nor4_1 U7197 ( .ip1(n10054), .ip2(n6428), .ip3(n6427), .ip4(n6426), .op(
        n6440) );
  nor4_1 U7198 ( .ip1(n10054), .ip2(n10053), .ip3(n10052), .ip4(n10427), .op(
        n10055) );
  nor4_1 U7199 ( .ip1(n6867), .ip2(n6866), .ip3(n6865), .ip4(n6864), .op(n9371) );
  buf_1 U7200 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12722) );
  buf_1 U7201 ( .ip(n12722), .op(n12715) );
  buf_1 U7202 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12717) );
  buf_1 U7203 ( .ip(n12717), .op(n12716) );
  buf_1 U7204 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12725) );
  buf_1 U7205 ( .ip(n12725), .op(n12718) );
  buf_1 U7206 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12713) );
  buf_1 U7207 ( .ip(n12713), .op(n12703) );
  buf_1 U7208 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12706) );
  buf_1 U7209 ( .ip(n12709), .op(n12704) );
  buf_1 U7210 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12721) );
  buf_1 U7211 ( .ip(n12721), .op(n12705) );
  buf_1 U7212 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12712) );
  buf_1 U7213 ( .ip(n12712), .op(n12708) );
  buf_1 U7214 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12719) );
  buf_1 U7215 ( .ip(n12719), .op(n12710) );
  buf_1 U7216 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12728) );
  buf_1 U7217 ( .ip(n12728), .op(n12730) );
  buf_1 U7218 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12702) );
  buf_1 U7219 ( .ip(n12702), .op(n12726) );
  buf_1 U7220 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12735) );
  buf_1 U7221 ( .ip(n12735), .op(n12736) );
  buf_1 U7222 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12727) );
  buf_1 U7223 ( .ip(n12727), .op(n12720) );
  buf_1 U7224 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12729) );
  buf_1 U7225 ( .ip(n12729), .op(n12723) );
  buf_1 U7226 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12731) );
  buf_1 U7227 ( .ip(n12731), .op(n12724) );
  buf_1 U7228 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12733) );
  buf_1 U7229 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12707) );
  buf_1 U7230 ( .ip(n12707), .op(n12701) );
  buf_1 U7231 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12714) );
  buf_1 U7232 ( .ip(n12714), .op(n12697) );
  buf_1 U7233 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12700) );
  buf_1 U7234 ( .ip(n12707), .op(n12699) );
  buf_1 U7235 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12709) );
  buf_1 U7236 ( .ip(n12709), .op(n12698) );
  buf_1 U7237 ( .ip(n12710), .op(n12711) );
  buf_1 U7238 ( .ip(n12710), .op(n12696) );
  buf_1 U7239 ( .ip(n12732), .op(n12695) );
  inv_1 U7240 ( .ip(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .op(n12118) );
  nand2_1 U7241 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Fjgvx4 ), .op(n7079) );
  inv_1 U7242 ( .ip(n7079), .op(n10200) );
  inv_1 U7243 ( .ip(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(n11786) );
  inv_1 U7244 ( .ip(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .op(n12117) );
  inv_1 U7245 ( .ip(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .op(n8424) );
  nand2_1 U7246 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n8424), .op(
        n12126) );
  inv_1 U7247 ( .ip(n12126), .op(n12619) );
  nand2_1 U7248 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Z6gvx4 ), .op(n10722) );
  inv_1 U7249 ( .ip(n10722), .op(n10764) );
  inv_1 U7250 ( .ip(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .op(n11228) );
  nand2_1 U7251 ( .ip1(n10764), .ip2(n11228), .op(n11010) );
  inv_1 U7252 ( .ip(n11010), .op(n10888) );
  nand2_1 U7253 ( .ip1(n12619), .ip2(n10888), .op(n6270) );
  nor2_1 U7254 ( .ip1(n11786), .ip2(n6270), .op(n6191) );
  inv_1 U7255 ( .ip(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .op(n11693) );
  nor2_1 U7256 ( .ip1(n12126), .ip2(n11693), .op(n11267) );
  inv_1 U7257 ( .ip(n11267), .op(n6225) );
  nand2_1 U7258 ( .ip1(n12118), .ip2(n9807), .op(n10851) );
  nor2_1 U7259 ( .ip1(n6225), .ip2(n10851), .op(n6252) );
  nor3_1 U7260 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip3(n10722), .op(n9789) );
  inv_1 U7261 ( .ip(n9789), .op(n6190) );
  inv_1 U7262 ( .ip(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .op(n12588) );
  nor2_1 U7263 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(n12588), .op(
        n10932) );
  inv_1 U7264 ( .ip(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .op(n11100) );
  nor2_1 U7265 ( .ip1(n9807), .ip2(n11100), .op(n9955) );
  inv_1 U7266 ( .ip(n9955), .op(n10833) );
  nor2_1 U7267 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n10833), .op(
        n10651) );
  nand2_1 U7268 ( .ip1(n10932), .ip2(n10651), .op(n10486) );
  nand2_1 U7269 ( .ip1(n6190), .ip2(n10486), .op(n6274) );
  nor4_1 U7270 ( .ip1(n10200), .ip2(n6191), .ip3(n6252), .ip4(n6274), .op(
        n6216) );
  nand2_1 U7271 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Mcgvx4 ), .op(n11015) );
  inv_1 U7272 ( .ip(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .op(n12623) );
  nand2_1 U7273 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n12623), .op(
        n6859) );
  inv_1 U7274 ( .ip(n6859), .op(n12132) );
  nand2_1 U7275 ( .ip1(n12132), .ip2(\CORTEXM0DS_INST/u_logic/Q5gvx4 ), .op(
        n9927) );
  nor2_1 U7276 ( .ip1(n11015), .ip2(n9927), .op(n6208) );
  nand2_1 U7277 ( .ip1(n11228), .ip2(n11786), .op(n10971) );
  inv_1 U7278 ( .ip(n10971), .op(n11132) );
  nand2_1 U7279 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n11132), .op(
        n6271) );
  nor2_1 U7280 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n6271), .op(
        n6207) );
  inv_1 U7281 ( .ip(\CORTEXM0DS_INST/vis_pc [2]), .op(n8587) );
  inv_1 U7282 ( .ip(\CORTEXM0DS_INST/u_logic/Eg8vx4 ), .op(n6192) );
  nor3_1 U7283 ( .ip1(\CORTEXM0DS_INST/u_logic/Ki8vx4 ), .ip2(n8587), .ip3(
        n6192), .op(n11131) );
  nor2_1 U7284 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(n11051) );
  nand2_1 U7285 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n11051), .op(
        n10988) );
  inv_1 U7286 ( .ip(n10988), .op(n12121) );
  nand2_1 U7287 ( .ip1(n12121), .ip2(n11796), .op(n11216) );
  nor2_1 U7288 ( .ip1(n11131), .ip2(n11216), .op(n6221) );
  nand2_1 U7289 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n8424), .op(
        n11253) );
  nor2_1 U7290 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n10851), .op(
        n9962) );
  inv_1 U7291 ( .ip(n9962), .op(n6349) );
  nor2_1 U7292 ( .ip1(n11253), .ip2(n6349), .op(n6193) );
  or2_1 U7293 ( .ip1(n6221), .ip2(n6193), .op(n6254) );
  inv_1 U7294 ( .ip(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .op(n12599) );
  nand2_1 U7295 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n12599), .op(
        n10842) );
  inv_1 U7296 ( .ip(n10842), .op(n10551) );
  nand2_1 U7297 ( .ip1(n10551), .ip2(n10492), .op(n6195) );
  nor2_1 U7298 ( .ip1(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip2(n9807), .op(
        n10647) );
  nand2_1 U7299 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Fb9vx4 ), .op(n10820) );
  nand2_1 U7300 ( .ip1(n10647), .ip2(n10820), .op(n6194) );
  nand2_1 U7301 ( .ip1(n6195), .ip2(n6194), .op(n6237) );
  nand2_1 U7302 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n12117), .op(
        n9377) );
  nor2_1 U7303 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Cn8vx4 ), .op(n10873) );
  inv_1 U7304 ( .ip(n10873), .op(n10795) );
  nor3_1 U7305 ( .ip1(n11228), .ip2(n9377), .ip3(n10795), .op(n6281) );
  nor2_1 U7306 ( .ip1(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip2(n11100), .op(
        n9082) );
  inv_1 U7307 ( .ip(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .op(n10492) );
  nand2_1 U7308 ( .ip1(n9082), .ip2(n10492), .op(n9771) );
  inv_1 U7309 ( .ip(n9771), .op(n6409) );
  nand3_1 U7310 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n6409), .ip3(
        n10873), .op(n10779) );
  nor2_1 U7311 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n10779), .op(
        n11803) );
  and2_1 U7312 ( .ip1(n11228), .ip2(n11803), .op(n6196) );
  not_ab_or_c_or_d U7313 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(n6237), 
        .ip3(n6281), .ip4(n6196), .op(n6266) );
  inv_1 U7314 ( .ip(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .op(n12538) );
  nor2_1 U7315 ( .ip1(n9807), .ip2(n12538), .op(n11090) );
  inv_1 U7316 ( .ip(\CORTEXM0DS_INST/u_logic/Ho8vx4 ), .op(n12122) );
  nand2_1 U7317 ( .ip1(n11100), .ip2(n12122), .op(n10539) );
  inv_1 U7318 ( .ip(n10539), .op(n10869) );
  inv_1 U7319 ( .ip(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .op(n12592) );
  nand2_1 U7320 ( .ip1(n9955), .ip2(n12592), .op(n11088) );
  nor3_1 U7321 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip3(n11088), .op(n6197) );
  or2_1 U7322 ( .ip1(n10869), .ip2(n6197), .op(n6198) );
  nand2_1 U7323 ( .ip1(n11090), .ip2(n6198), .op(n6206) );
  inv_1 U7324 ( .ip(\CORTEXM0DS_INST/u_logic/P39vx4 ), .op(n12558) );
  nor2_1 U7325 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n9807), .op(
        n10933) );
  nor2_1 U7326 ( .ip1(n12592), .ip2(n10842), .op(n11107) );
  nor2_1 U7327 ( .ip1(n10933), .ip2(n11107), .op(n8581) );
  inv_1 U7328 ( .ip(n10647), .op(n6267) );
  nor2_1 U7329 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n6267), .op(
        n12320) );
  inv_1 U7330 ( .ip(n12320), .op(n6219) );
  nand2_1 U7331 ( .ip1(n10551), .ip2(n12538), .op(n9886) );
  nand2_1 U7332 ( .ip1(n6219), .ip2(n9886), .op(n10990) );
  inv_1 U7333 ( .ip(n10990), .op(n6199) );
  nor2_1 U7334 ( .ip1(n8581), .ip2(n6199), .op(n9868) );
  nand3_1 U7335 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/R89vx4 ), .op(n6200) );
  nor2_1 U7336 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Mc9vx4 ), .op(n9667) );
  inv_1 U7337 ( .ip(\CORTEXM0DS_INST/u_logic/K79vx4 ), .op(n12567) );
  nor2_1 U7338 ( .ip1(\CORTEXM0DS_INST/u_logic/R89vx4 ), .ip2(n12567), .op(
        n9828) );
  nand3_1 U7339 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip3(n9828), .op(n9937) );
  and2_1 U7340 ( .ip1(n9667), .ip2(n9937), .op(n6287) );
  nor2_1 U7341 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n10842), .op(
        n10803) );
  inv_1 U7342 ( .ip(n10803), .op(n10491) );
  not_ab_or_c_or_d U7343 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n6200), 
        .ip3(n6287), .ip4(n10491), .op(n6201) );
  nor2_1 U7344 ( .ip1(n9868), .ip2(n6201), .op(n6202) );
  nor2_1 U7345 ( .ip1(\CORTEXM0DS_INST/u_logic/Ho8vx4 ), .ip2(n6202), .op(
        n6204) );
  nand3_1 U7346 ( .ip1(\CORTEXM0DS_INST/vis_pc [27]), .ip2(
        \CORTEXM0DS_INST/vis_pc [28]), .ip3(\CORTEXM0DS_INST/vis_pc [29]), 
        .op(n10457) );
  inv_1 U7347 ( .ip(n10457), .op(n6203) );
  nor3_1 U7348 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [5]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [4]), .ip3(\CORTEXM0DS_INST/vis_ipsr [3]), 
        .op(n12403) );
  nor3_1 U7349 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [2]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [1]), .ip3(\CORTEXM0DS_INST/vis_ipsr [0]), 
        .op(n6377) );
  nand2_1 U7350 ( .ip1(n12403), .ip2(n6377), .op(n11811) );
  nand4_1 U7351 ( .ip1(\CORTEXM0DS_INST/u_logic/Hx8vx4 ), .ip2(
        \CORTEXM0DS_INST/vis_pc [30]), .ip3(n6203), .ip4(n11811), .op(n10770)
         );
  inv_1 U7352 ( .ip(n10770), .op(n12138) );
  nand2_1 U7353 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n12118), .op(
        n12128) );
  nor2_1 U7354 ( .ip1(n12138), .ip2(n12128), .op(n11802) );
  not_ab_or_c_or_d U7355 ( .ip1(n11803), .ip2(n12558), .ip3(n6204), .ip4(
        n11802), .op(n6205) );
  inv_1 U7356 ( .ip(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .op(n11796) );
  nand2_1 U7357 ( .ip1(n11796), .ip2(n9807), .op(n9943) );
  inv_1 U7358 ( .ip(n9943), .op(n10632) );
  nor2_1 U7359 ( .ip1(n11693), .ip2(n11786), .op(n11248) );
  nand4_1 U7360 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10632), .ip3(
        n11248), .ip4(n11228), .op(n9779) );
  nand4_1 U7361 ( .ip1(n6266), .ip2(n6206), .ip3(n6205), .ip4(n9779), .op(
        n6273) );
  nor4_1 U7362 ( .ip1(n6208), .ip2(n6207), .ip3(n6254), .ip4(n6273), .op(n6215) );
  nor4_1 U7363 ( .ip1(\CORTEXM0DS_INST/u_logic/Bx9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Wv9vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Su9vx4 ), .ip4(
        \CORTEXM0DS_INST/u_logic/Ot9vx4 ), .op(n9044) );
  inv_1 U7364 ( .ip(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .op(n12104) );
  nor2_1 U7365 ( .ip1(n9044), .ip2(n12104), .op(n12108) );
  nor3_1 U7366 ( .ip1(\CORTEXM0DS_INST/u_logic/Wv9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Su9vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Ot9vx4 ), .op(n6209) );
  inv_1 U7367 ( .ip(\CORTEXM0DS_INST/u_logic/Bx9vx4 ), .op(n12384) );
  nor2_1 U7368 ( .ip1(n6209), .ip2(n12384), .op(n12397) );
  inv_1 U7369 ( .ip(\CORTEXM0DS_INST/u_logic/Su9vx4 ), .op(n12373) );
  inv_1 U7370 ( .ip(\CORTEXM0DS_INST/u_logic/Ot9vx4 ), .op(n11206) );
  nor2_1 U7371 ( .ip1(n12373), .ip2(n11206), .op(n12381) );
  nor2_1 U7372 ( .ip1(\CORTEXM0DS_INST/u_logic/Su9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Ot9vx4 ), .op(n6210) );
  inv_1 U7373 ( .ip(\CORTEXM0DS_INST/u_logic/Wv9vx4 ), .op(n12362) );
  nor2_1 U7374 ( .ip1(n6210), .ip2(n12362), .op(n12370) );
  nand2_1 U7375 ( .ip1(n9044), .ip2(n12104), .op(n9014) );
  nand2_1 U7376 ( .ip1(\CORTEXM0DS_INST/u_logic/Cq9vx4 ), .ip2(n9014), .op(
        n12079) );
  inv_1 U7377 ( .ip(\CORTEXM0DS_INST/u_logic/Gr9vx4 ), .op(n6211) );
  nor2_1 U7378 ( .ip1(n9014), .ip2(\CORTEXM0DS_INST/u_logic/Cq9vx4 ), .op(
        n9000) );
  or2_1 U7379 ( .ip1(n6211), .ip2(n9000), .op(n10224) );
  nand2_1 U7380 ( .ip1(n9000), .ip2(n6211), .op(n9043) );
  nand2_1 U7381 ( .ip1(\CORTEXM0DS_INST/u_logic/Ks9vx4 ), .ip2(n9043), .op(
        n10204) );
  inv_1 U7382 ( .ip(n10955), .op(n10892) );
  nand2_1 U7383 ( .ip1(n10892), .ip2(n12121), .op(n6277) );
  or2_1 U7384 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n6277), .op(n6214) );
  nor2_1 U7385 ( .ip1(n12592), .ip2(n10492), .op(n10512) );
  inv_1 U7386 ( .ip(n10512), .op(n9952) );
  nand2_1 U7387 ( .ip1(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip2(n10492), .op(
        n9948) );
  nand3_1 U7388 ( .ip1(n9955), .ip2(n9952), .ip3(n9948), .op(n6213) );
  nand4_1 U7389 ( .ip1(n6216), .ip2(n6215), .ip3(n6214), .ip4(n6213), .op(
        n2167) );
  nand2_1 U7390 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n12623), .op(
        n10852) );
  inv_1 U7391 ( .ip(n10852), .op(n10421) );
  or2_1 U7392 ( .ip1(n10421), .ip2(n10200), .op(n6218) );
  inv_1 U7393 ( .ip(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .op(n12125) );
  nand2_1 U7394 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n12125), .op(
        n10673) );
  nor2_1 U7395 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n10673), .op(
        n10922) );
  inv_1 U7396 ( .ip(n10922), .op(n10949) );
  nor2_1 U7397 ( .ip1(n11796), .ip2(n10949), .op(n10983) );
  or2_1 U7398 ( .ip1(n10983), .ip2(n10200), .op(n6217) );
  nand2_1 U7399 ( .ip1(n6218), .ip2(n6217), .op(n10425) );
  nor2_1 U7400 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n11228), .op(
        n9853) );
  nand2_1 U7401 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Mcgvx4 ), .op(n12072) );
  nor3_1 U7402 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n11786), .ip3(
        n12072), .op(n9773) );
  nor2_1 U7403 ( .ip1(n12126), .ip2(n6859), .op(n10762) );
  inv_1 U7404 ( .ip(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .op(n12609) );
  nand2_1 U7405 ( .ip1(n10762), .ip2(n12609), .op(n10201) );
  nor2_1 U7406 ( .ip1(n11796), .ip2(n10201), .op(n6261) );
  not_ab_or_c_or_d U7407 ( .ip1(n9853), .ip2(n12132), .ip3(n9773), .ip4(n6261), 
        .op(n6236) );
  nand2_1 U7408 ( .ip1(n10873), .ip2(n12623), .op(n10739) );
  nand2_1 U7409 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n11796), .op(
        n10479) );
  nor3_1 U7410 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10739), .ip3(
        n10479), .op(n6220) );
  nand2_1 U7411 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n10869), .op(
        n10542) );
  nor2_1 U7412 ( .ip1(n10542), .ip2(n6219), .op(n10490) );
  or2_1 U7413 ( .ip1(n6220), .ip2(n10490), .op(n6223) );
  nand2_1 U7414 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n12588), .op(
        n9963) );
  nand2_1 U7415 ( .ip1(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip2(n10647), .op(
        n11089) );
  nor3_1 U7416 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Ho8vx4 ), .op(n9870) );
  inv_1 U7417 ( .ip(n9870), .op(n9884) );
  not_ab_or_c_or_d U7418 ( .ip1(n9963), .ip2(n10492), .ip3(n11089), .ip4(n9884), .op(n6222) );
  not_ab_or_c_or_d U7419 ( .ip1(n12125), .ip2(n6223), .ip3(n6222), .ip4(n6221), 
        .op(n6235) );
  nand3_1 U7420 ( .ip1(n11803), .ip2(n11228), .ip3(n12125), .op(n9905) );
  inv_1 U7421 ( .ip(n9905), .op(n6233) );
  nand2_1 U7422 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n11796), .op(
        n11240) );
  nor3_1 U7423 ( .ip1(n10955), .ip2(n6859), .ip3(n11240), .op(n6262) );
  inv_1 U7424 ( .ip(\CORTEXM0DS_INST/u_logic/D69vx4 ), .op(n12562) );
  inv_1 U7425 ( .ip(n9828), .op(n10837) );
  nor2_1 U7426 ( .ip1(n12562), .ip2(n10837), .op(n6258) );
  inv_1 U7427 ( .ip(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .op(n11190) );
  nand3_1 U7428 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(n6258), .ip3(
        n11190), .op(n10715) );
  nor2_1 U7429 ( .ip1(n11100), .ip2(n12599), .op(n10206) );
  nor2_1 U7430 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Sh9vx4 ), .op(n10818) );
  nand4_1 U7431 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n10206), .ip3(
        n10818), .ip4(n11090), .op(n11110) );
  nor3_1 U7432 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n10715), .ip3(
        n11110), .op(n6231) );
  nand2_1 U7433 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/R89vx4 ), .op(n10623) );
  nor2_1 U7434 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n10492), .op(
        n11101) );
  inv_1 U7435 ( .ip(n11101), .op(n10794) );
  nor2_1 U7436 ( .ip1(n11100), .ip2(n10794), .op(n11108) );
  nand2_1 U7437 ( .ip1(n11108), .ip2(n11090), .op(n10572) );
  inv_1 U7438 ( .ip(n10572), .op(n12389) );
  nand2_1 U7439 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n12389), .op(
        n12378) );
  nand4_1 U7440 ( .ip1(n9667), .ip2(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip3(
        n12567), .ip4(n12562), .op(n6224) );
  nor3_1 U7441 ( .ip1(n10623), .ip2(n12378), .ip3(n6224), .op(n6230) );
  nor2_1 U7442 ( .ip1(n12125), .ip2(n11216), .op(n6229) );
  nand2_1 U7443 ( .ip1(n12118), .ip2(n12125), .op(n10782) );
  nor2_1 U7444 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n10782), .op(
        n11099) );
  inv_1 U7445 ( .ip(n11099), .op(n10796) );
  or2_1 U7446 ( .ip1(n6225), .ip2(n10796), .op(n6227) );
  nand2_1 U7447 ( .ip1(n11693), .ip2(n11228), .op(n6842) );
  or2_1 U7448 ( .ip1(n6842), .ip2(n10796), .op(n6226) );
  nand2_1 U7449 ( .ip1(n6227), .ip2(n6226), .op(n6228) );
  or4_1 U7450 ( .ip1(n6231), .ip2(n6230), .ip3(n6229), .ip4(n6228), .op(n6232)
         );
  not_ab_or_c_or_d U7451 ( .ip1(n6233), .ip2(\CORTEXM0DS_INST/u_logic/P39vx4 ), 
        .ip3(n6262), .ip4(n6232), .op(n6234) );
  nand4_1 U7452 ( .ip1(n10425), .ip2(n6236), .ip3(n6235), .ip4(n6234), .op(
        n3317) );
  nor2_1 U7453 ( .ip1(n11100), .ip2(n10491), .op(n10862) );
  nand2_1 U7454 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Cf9vx4 ), .op(n12321) );
  nor3_1 U7455 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n10492), .ip3(
        n12321), .op(n6251) );
  not_ab_or_c_or_d U7456 ( .ip1(n10803), .ip2(n11190), .ip3(n6251), .ip4(n6237), .op(n6238) );
  nor2_1 U7457 ( .ip1(\CORTEXM0DS_INST/u_logic/Ho8vx4 ), .ip2(n6238), .op(
        n6244) );
  nand2_1 U7458 ( .ip1(n12592), .ip2(n12538), .op(n10835) );
  inv_1 U7459 ( .ip(n10835), .op(n10635) );
  inv_1 U7460 ( .ip(\CORTEXM0DS_INST/u_logic/R89vx4 ), .op(n12571) );
  not_ab_or_c_or_d U7461 ( .ip1(n10635), .ip2(n12571), .ip3(n9807), .ip4(
        n10539), .op(n6243) );
  nor2_1 U7462 ( .ip1(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Cf9vx4 ), .op(n9834) );
  nand2_1 U7463 ( .ip1(n10492), .ip2(n12122), .op(n10664) );
  nor2_1 U7464 ( .ip1(n6267), .ip2(n10664), .op(n6239) );
  not_ab_or_c_or_d U7465 ( .ip1(n9834), .ip2(n9955), .ip3(n11802), .ip4(n6239), 
        .op(n6242) );
  nand2_1 U7466 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(n12588), .op(
        n10481) );
  nor2_1 U7467 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n10481), .op(
        n9933) );
  nor2_1 U7468 ( .ip1(\CORTEXM0DS_INST/u_logic/K79vx4 ), .ip2(n12571), .op(
        n10979) );
  inv_1 U7469 ( .ip(n10979), .op(n6240) );
  nand3_1 U7470 ( .ip1(n9933), .ip2(n10651), .ip3(n6240), .op(n6241) );
  nand3_1 U7471 ( .ip1(n6242), .ip2(n10486), .ip3(n6241), .op(n6253) );
  nor4_1 U7472 ( .ip1(n10862), .ip2(n6244), .ip3(n6243), .ip4(n6253), .op(
        n6247) );
  nand2_1 U7473 ( .ip1(n10764), .ip2(n11693), .op(n6246) );
  nor2_1 U7474 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Whgvx4 ), .op(n9388) );
  nand2_1 U7475 ( .ip1(n12132), .ip2(n9388), .op(n6269) );
  inv_1 U7476 ( .ip(n11088), .op(n9968) );
  nand3_1 U7477 ( .ip1(n9968), .ip2(n12588), .ip3(n11190), .op(n6245) );
  nand4_1 U7478 ( .ip1(n6247), .ip2(n6246), .ip3(n6269), .ip4(n6245), .op(
        n3369) );
  nand4_1 U7479 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip4(n12592), .op(n10848) );
  nor2_1 U7480 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n12118), .op(
        n9785) );
  nand2_1 U7481 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n9785), .op(
        n10523) );
  nand2_1 U7482 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Ho8vx4 ), .op(n5092) );
  inv_1 U7483 ( .ip(n5092), .op(n8982) );
  nand2_1 U7484 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n8982), .op(
        n6249) );
  nand3_1 U7485 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n10512), .ip3(
        n11100), .op(n6248) );
  nand4_1 U7486 ( .ip1(n10848), .ip2(n10523), .ip3(n6249), .ip4(n6248), .op(
        n6250) );
  nor3_1 U7487 ( .ip1(n6252), .ip2(n6251), .ip3(n6250), .op(n6265) );
  nor2_1 U7488 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n12623), .op(
        n12369) );
  nor3_1 U7489 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip3(n11786), .op(n11258) );
  nand2_1 U7490 ( .ip1(n12369), .ip2(n11258), .op(n12123) );
  nor2_1 U7491 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n12123), .op(
        n9776) );
  not_ab_or_c_or_d U7492 ( .ip1(\CORTEXM0DS_INST/u_logic/Ho8vx4 ), .ip2(n9776), 
        .ip3(n6254), .ip4(n6253), .op(n6264) );
  nand2_1 U7493 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n12132), .op(
        n10972) );
  inv_1 U7494 ( .ip(n11051), .op(n11763) );
  or2_1 U7495 ( .ip1(n10972), .ip2(n11763), .op(n6257) );
  nand2_1 U7496 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n11796), .op(
        n6255) );
  or2_1 U7497 ( .ip1(n6255), .ip2(n11763), .op(n6256) );
  nand2_1 U7498 ( .ip1(n6257), .ip2(n6256), .op(n6260) );
  nor2_1 U7499 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Fb9vx4 ), .op(n10500) );
  nor2_1 U7500 ( .ip1(n6258), .ip2(n12588), .op(n10931) );
  nor4_1 U7501 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n10500), .ip3(
        n10931), .ip4(n11088), .op(n6259) );
  nor4_1 U7502 ( .ip1(n6262), .ip2(n6261), .ip3(n6260), .ip4(n6259), .op(n6263) );
  nand4_1 U7503 ( .ip1(n6266), .ip2(n6265), .ip3(n6264), .ip4(n6263), .op(
        n1743) );
  nor2_1 U7504 ( .ip1(n10851), .ip2(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(
        n10652) );
  nand2_1 U7505 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(n8424), .op(
        n12628) );
  nor3_1 U7506 ( .ip1(n10852), .ip2(n10851), .ip3(n12628), .op(n9777) );
  nor3_1 U7507 ( .ip1(n12588), .ip2(n6267), .ip3(n10664), .op(n6268) );
  not_ab_or_c_or_d U7508 ( .ip1(n12619), .ip2(n10652), .ip3(n9777), .ip4(n6268), .op(n6279) );
  nor3_1 U7509 ( .ip1(n12118), .ip2(n12117), .ip3(n8424), .op(n11076) );
  nand2_1 U7510 ( .ip1(\CORTEXM0DS_INST/u_logic/Q5gvx4 ), .ip2(n11076), .op(
        n10679) );
  nor2_1 U7511 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n10679), .op(
        n6275) );
  nand4_1 U7512 ( .ip1(n7079), .ip2(n6271), .ip3(n6270), .ip4(n6269), .op(
        n6272) );
  nor4_1 U7513 ( .ip1(n6275), .ip2(n6274), .ip3(n6273), .ip4(n6272), .op(n6278) );
  nand2_1 U7514 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n9968), .op(
        n6276) );
  nand4_1 U7515 ( .ip1(n6279), .ip2(n6278), .ip3(n6277), .ip4(n6276), .op(
        n4619) );
  nand2_1 U7516 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(n11223) );
  nor2_1 U7517 ( .ip1(n12609), .ip2(n11223), .op(n11262) );
  inv_1 U7518 ( .ip(n11262), .op(n12071) );
  nand2_1 U7519 ( .ip1(n12071), .ip2(n10523), .op(n10798) );
  inv_1 U7520 ( .ip(n10798), .op(n6291) );
  inv_1 U7521 ( .ip(n11089), .op(n11146) );
  and2_1 U7522 ( .ip1(n11108), .ip2(n11146), .op(n10965) );
  nand2_1 U7523 ( .ip1(n11796), .ip2(n11228), .op(n11218) );
  nand2_1 U7524 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Efgvx4 ), .op(n10864) );
  inv_1 U7525 ( .ip(n10864), .op(n11773) );
  not_ab_or_c_or_d U7526 ( .ip1(n11218), .ip2(n10972), .ip3(n11773), .ip4(
        n12072), .op(n6286) );
  nand2_1 U7527 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n12609), .op(
        n12627) );
  inv_1 U7528 ( .ip(n12627), .op(n11275) );
  nand4_1 U7529 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n11275), .ip3(
        n11228), .ip4(n12623), .op(n11764) );
  nor2_1 U7530 ( .ip1(n11764), .ip2(n10988), .op(n6280) );
  nand3_1 U7531 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n10873), .ip3(
        n11786), .op(n9780) );
  nor2_1 U7532 ( .ip1(n9780), .ip2(n10673), .op(n9858) );
  not_ab_or_c_or_d U7533 ( .ip1(n6281), .ip2(n12125), .ip3(n6280), .ip4(n9858), 
        .op(n6284) );
  nor2_1 U7534 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n12117), .op(
        n11065) );
  nand2_1 U7535 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n11248), .op(
        n8157) );
  inv_1 U7536 ( .ip(n8157), .op(n9945) );
  and3_1 U7537 ( .ip1(n10632), .ip2(n11065), .ip3(n9945), .op(n10555) );
  nand2_1 U7538 ( .ip1(n10555), .ip2(n12125), .op(n6441) );
  nand3_1 U7539 ( .ip1(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip2(n11101), .ip3(
        n9968), .op(n6283) );
  nor2_1 U7540 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Mcgvx4 ), .op(n11066) );
  nand2_1 U7541 ( .ip1(n11066), .ip2(n10983), .op(n6282) );
  nand4_1 U7542 ( .ip1(n6284), .ip2(n6441), .ip3(n6283), .ip4(n6282), .op(
        n6285) );
  not_ab_or_c_or_d U7543 ( .ip1(n10965), .ip2(n10820), .ip3(n6286), .ip4(n6285), .op(n6290) );
  nor2_1 U7544 ( .ip1(n10794), .ip2(n9886), .op(n11181) );
  nand2_1 U7545 ( .ip1(n10869), .ip2(n11181), .op(n8986) );
  or2_1 U7546 ( .ip1(n6287), .ip2(n8986), .op(n6289) );
  nand2_1 U7547 ( .ip1(n11090), .ip2(n12599), .op(n10806) );
  or4_1 U7548 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip3(n11100), .ip4(n10806), .op(
        n6288) );
  nand4_1 U7549 ( .ip1(n6291), .ip2(n6290), .ip3(n6289), .ip4(n6288), .op(
        n1788) );
  nor2_1 U7550 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n11131), .op(
        n10043) );
  nand2_1 U7551 ( .ip1(n11796), .ip2(n10955), .op(n6431) );
  nor2_1 U7552 ( .ip1(n10043), .ip2(n6431), .op(n10989) );
  nand2_1 U7553 ( .ip1(n12609), .ip2(n8424), .op(n7017) );
  nor2_1 U7554 ( .ip1(n6859), .ip2(n7017), .op(n10758) );
  nor2_1 U7555 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n12609), .op(
        n8358) );
  nand2_1 U7556 ( .ip1(n12117), .ip2(n9807), .op(n11690) );
  inv_1 U7557 ( .ip(n11690), .op(n9946) );
  nor2_1 U7558 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n12609), .op(
        n9730) );
  inv_1 U7559 ( .ip(n9730), .op(n11692) );
  inv_1 U7560 ( .ip(n10851), .op(n9941) );
  nand2_1 U7561 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n9941), .op(
        n11277) );
  or2_1 U7562 ( .ip1(n11692), .ip2(n11277), .op(n6293) );
  nand2_1 U7563 ( .ip1(n11228), .ip2(n10770), .op(n10531) );
  or2_1 U7564 ( .ip1(n10531), .ip2(n11277), .op(n6292) );
  nand2_1 U7565 ( .ip1(n6293), .ip2(n6292), .op(n6294) );
  not_ab_or_c_or_d U7566 ( .ip1(n8358), .ip2(n9946), .ip3(n10556), .ip4(n6294), 
        .op(n6295) );
  or2_1 U7567 ( .ip1(n6295), .ip2(n12125), .op(n6298) );
  inv_1 U7568 ( .ip(n11240), .op(n10530) );
  nor2_1 U7569 ( .ip1(n12623), .ip2(n10530), .op(n10689) );
  or2_1 U7570 ( .ip1(n6349), .ip2(n10689), .op(n6296) );
  or2_1 U7571 ( .ip1(n6296), .ip2(n12125), .op(n6297) );
  nand2_1 U7572 ( .ip1(n6298), .ip2(n6297), .op(n6309) );
  nor2_1 U7573 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Mcgvx4 ), .op(n10478) );
  inv_1 U7574 ( .ip(n10478), .op(n11788) );
  nor2_1 U7575 ( .ip1(n9927), .ip2(n11788), .op(n10516) );
  nor2_1 U7576 ( .ip1(n11786), .ip2(n10679), .op(n11686) );
  nand2_1 U7577 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n11786), .op(
        n11243) );
  nor2_1 U7578 ( .ip1(n11243), .ip2(n11010), .op(n10515) );
  not_ab_or_c_or_d U7579 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n10516), .ip3(n11686), .ip4(n10515), .op(n6307) );
  nor2_1 U7580 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n11693), .op(
        n9374) );
  nand3_1 U7581 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n9374), .ip3(
        n10764), .op(n6430) );
  inv_1 U7582 ( .ip(n6430), .op(n11794) );
  nand2_1 U7583 ( .ip1(n12117), .ip2(n11228), .op(n10973) );
  inv_1 U7584 ( .ip(n9785), .op(n11789) );
  not_ab_or_c_or_d U7585 ( .ip1(n11786), .ip2(n10973), .ip3(
        \CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip4(n11789), .op(n6300) );
  nand2_1 U7586 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n12619), .op(
        n10671) );
  nor2_1 U7587 ( .ip1(n12128), .ip2(n10671), .op(n6299) );
  nor2_1 U7588 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n11228), .op(
        n11256) );
  nand2_1 U7589 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n11256), .op(
        n11765) );
  inv_1 U7590 ( .ip(n11765), .op(n10814) );
  inv_1 U7591 ( .ip(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .op(n5639) );
  inv_1 U7592 ( .ip(n10739), .op(n10203) );
  nor2_1 U7593 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n8424), .op(
        n9659) );
  nor2_1 U7594 ( .ip1(n12117), .ip2(n11228), .op(n9573) );
  nand2_1 U7595 ( .ip1(n9659), .ip2(n9573), .op(n6435) );
  nor2_1 U7596 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n6435), .op(
        n6786) );
  or2_1 U7597 ( .ip1(n10203), .ip2(n6786), .op(n6302) );
  inv_1 U7598 ( .ip(n12128), .op(n11779) );
  or2_1 U7599 ( .ip1(n11779), .ip2(n6786), .op(n6301) );
  nand2_1 U7600 ( .ip1(n6302), .ip2(n6301), .op(n6303) );
  nor2_1 U7601 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n11693), .op(
        n12641) );
  inv_1 U7602 ( .ip(n12641), .op(n11682) );
  nor2_1 U7603 ( .ip1(n6303), .ip2(n11682), .op(n6304) );
  not_ab_or_c_or_d U7604 ( .ip1(n10814), .ip2(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip3(n6419), .ip4(n6304), .op(n6305) );
  nand2_1 U7605 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .op(n11689) );
  nand2_1 U7606 ( .ip1(n11796), .ip2(n10421), .op(n11756) );
  nor2_1 U7607 ( .ip1(n11689), .ip2(n11756), .op(n6866) );
  nand3_1 U7608 ( .ip1(n12641), .ip2(n6866), .ip3(n12117), .op(n6414) );
  not_ab_or_c_or_d U7609 ( .ip1(n10989), .ip2(n10758), .ip3(n6309), .ip4(n6308), .op(n6945) );
  inv_1 U7610 ( .ip(n11248), .op(n9928) );
  nand2_1 U7611 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n9928), .op(
        n10631) );
  nand2_1 U7612 ( .ip1(n12609), .ip2(n11228), .op(n9815) );
  nand2_1 U7613 ( .ip1(n9815), .ip2(n10973), .op(n6311) );
  nand2_1 U7614 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(n10944) );
  nor3_1 U7615 ( .ip1(n12609), .ip2(n12117), .ip3(n10944), .op(n6310) );
  not_ab_or_c_or_d U7616 ( .ip1(n10631), .ip2(n6311), .ip3(n6310), .ip4(n10873), .op(n10028) );
  inv_1 U7617 ( .ip(n10028), .op(n8916) );
  nor3_1 U7618 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n9730), .ip3(
        n11228), .op(n8062) );
  nor2_1 U7619 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n12117), .op(
        n11230) );
  nor2_1 U7620 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(n11796), .op(
        n11209) );
  nand4_1 U7621 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip3(n11693), .ip4(n11786), .op(
        n9736) );
  inv_1 U7622 ( .ip(n9736), .op(n6316) );
  inv_1 U7623 ( .ip(n10782), .op(n11782) );
  nand3_1 U7624 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n11782), .ip3(
        n12609), .op(n10687) );
  or2_1 U7625 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10687), .op(
        n6314) );
  nor2_1 U7626 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n8424), .op(
        n11213) );
  inv_1 U7627 ( .ip(n11213), .op(n6312) );
  or2_1 U7628 ( .ip1(n6312), .ip2(n10687), .op(n6313) );
  nand2_1 U7629 ( .ip1(n6314), .ip2(n6313), .op(n6315) );
  not_ab_or_c_or_d U7630 ( .ip1(n11230), .ip2(n11209), .ip3(n6316), .ip4(n6315), .op(n6340) );
  nor2_1 U7631 ( .ip1(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip2(n9807), .op(
        n12618) );
  nand2_1 U7632 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n11228), .op(
        n10698) );
  inv_1 U7633 ( .ip(n11256), .op(n11793) );
  nor2_1 U7634 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(n11224) );
  inv_1 U7635 ( .ip(n11224), .op(n11239) );
  nor2_1 U7636 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Efgvx4 ), .op(n12633) );
  nand2_1 U7637 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n9807), .op(
        n10865) );
  inv_1 U7638 ( .ip(n10865), .op(n12653) );
  nand2_1 U7639 ( .ip1(n12633), .ip2(n12653), .op(n9402) );
  nor2_1 U7640 ( .ip1(n11239), .ip2(n9402), .op(n6320) );
  inv_1 U7641 ( .ip(n9388), .op(n9751) );
  or2_1 U7642 ( .ip1(n9751), .ip2(n10944), .op(n6318) );
  inv_1 U7643 ( .ip(n11689), .op(n11250) );
  nand2_1 U7644 ( .ip1(n11250), .ip2(n11786), .op(n11681) );
  or3_1 U7645 ( .ip1(n12609), .ip2(n12117), .ip3(n11681), .op(n6317) );
  not_ab_or_c_or_d U7646 ( .ip1(n6318), .ip2(n6317), .ip3(
        \CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip4(n12125), .op(n6319) );
  not_ab_or_c_or_d U7647 ( .ip1(n12618), .ip2(n6321), .ip3(n6320), .ip4(n6319), 
        .op(n6339) );
  nand2_1 U7648 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .op(n11252) );
  ab_or_c_or_d U7649 ( .ip1(n11682), .ip2(n11252), .ip3(
        \CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip4(n5639), .op(n6420) );
  nand4_1 U7650 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n11250), .ip3(
        n12641), .ip4(n12117), .op(n6322) );
  nand2_1 U7651 ( .ip1(n6420), .ip2(n6322), .op(n6323) );
  nand2_1 U7652 ( .ip1(\CORTEXM0DS_INST/u_logic/Rkgvx4 ), .ip2(n6323), .op(
        n6338) );
  nand2_1 U7653 ( .ip1(n11796), .ip2(n5639), .op(n11231) );
  nand2_1 U7654 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n12125), .op(
        n11680) );
  nor2_1 U7655 ( .ip1(n11231), .ip2(n11680), .op(n12654) );
  or2_1 U7656 ( .ip1(n9785), .ip2(n12654), .op(n6326) );
  nand2_1 U7657 ( .ip1(n5639), .ip2(n11786), .op(n6324) );
  or2_1 U7658 ( .ip1(n6324), .ip2(n12654), .op(n6325) );
  nand2_1 U7659 ( .ip1(n6326), .ip2(n6325), .op(n6335) );
  inv_1 U7660 ( .ip(n10673), .op(n12656) );
  inv_1 U7661 ( .ip(n9082), .op(n10696) );
  nand3_1 U7662 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n10539), .ip3(
        n10696), .op(n6410) );
  nand3_1 U7663 ( .ip1(n9771), .ip2(n11782), .ip3(n6410), .op(n6327) );
  nand2_1 U7664 ( .ip1(\CORTEXM0DS_INST/u_logic/W49vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/D69vx4 ), .op(n10683) );
  nand2_1 U7665 ( .ip1(n9828), .ip2(n10683), .op(n10697) );
  nand3_1 U7666 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n10818), .ip3(
        n10697), .op(n6407) );
  nand2_1 U7667 ( .ip1(n6327), .ip2(n6407), .op(n6329) );
  nor3_1 U7668 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n11689), .ip3(
        n10782), .op(n6328) );
  or2_1 U7669 ( .ip1(n6329), .ip2(n6328), .op(n6330) );
  nand2_1 U7670 ( .ip1(n11796), .ip2(n6330), .op(n6331) );
  inv_1 U7671 ( .ip(\CORTEXM0DS_INST/u_logic/Rkgvx4 ), .op(n10743) );
  nor2_1 U7672 ( .ip1(n6331), .ip2(n10743), .op(n6333) );
  nor3_1 U7673 ( .ip1(n12609), .ip2(n11693), .ip3(n11231), .op(n6332) );
  not_ab_or_c_or_d U7674 ( .ip1(n12656), .ip2(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip3(n6333), .ip4(n6332), .op(n6334) );
  inv_1 U7675 ( .ip(n11223), .op(n12624) );
  nand2_1 U7676 ( .ip1(n12624), .ip2(n10478), .op(n10810) );
  nand2_1 U7677 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n6336), .op(
        n6337) );
  nand2_1 U7678 ( .ip1(n8062), .ip2(n2139), .op(n6341) );
  nand2_1 U7679 ( .ip1(\CORTEXM0DS_INST/u_logic/A3gvx4 ), .ip2(n6341), .op(
        n12645) );
  nand2_1 U7680 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n11228), .op(
        n11232) );
  nor2_1 U7681 ( .ip1(n12118), .ip2(n11232), .op(n10813) );
  inv_1 U7682 ( .ip(n10813), .op(n10484) );
  inv_1 U7683 ( .ip(n11232), .op(n12655) );
  nand3_1 U7684 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n12655), .ip3(
        n9807), .op(n10487) );
  nand2_1 U7685 ( .ip1(n10484), .ip2(n10487), .op(n11061) );
  nand2_1 U7686 ( .ip1(n2139), .ip2(n11061), .op(n12111) );
  nand2_1 U7687 ( .ip1(n12645), .ip2(n12111), .op(n6346) );
  nand2_1 U7688 ( .ip1(\CORTEXM0DS_INST/u_logic/I4gvx4 ), .ip2(n6341), .op(
        n6971) );
  nor2_1 U7689 ( .ip1(\CORTEXM0DS_INST/u_logic/Xyfvx4 ), .ip2(n9807), .op(
        n6342) );
  or2_1 U7690 ( .ip1(n6971), .ip2(n6342), .op(n6344) );
  or2_1 U7691 ( .ip1(n12111), .ip2(n6342), .op(n6343) );
  nand2_1 U7692 ( .ip1(n6344), .ip2(n6343), .op(n6345) );
  mux2_1 U7693 ( .ip1(n6346), .ip2(n6345), .s(\CORTEXM0DS_INST/vis_pc [0]), 
        .op(n6421) );
  nor3_1 U7694 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip3(n10944), .op(n6834) );
  nand3_1 U7695 ( .ip1(n6834), .ip2(n10818), .ip3(
        \CORTEXM0DS_INST/u_logic/Rkgvx4 ), .op(n6348) );
  nand2_1 U7696 ( .ip1(n12609), .ip2(n12623), .op(n11683) );
  inv_1 U7697 ( .ip(n11683), .op(n12610) );
  nand2_1 U7698 ( .ip1(n12633), .ip2(n12610), .op(n6347) );
  not_ab_or_c_or_d U7699 ( .ip1(n6348), .ip2(n6347), .ip3(n9943), .ip4(n8424), 
        .op(n6418) );
  nor3_1 U7700 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n11239), .ip3(
        n6349), .op(n11684) );
  inv_1 U7701 ( .ip(\CORTEXM0DS_INST/vis_ipsr [2]), .op(n6359) );
  nand3_1 U7702 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [1]), .ip2(n12403), .ip3(
        n6359), .op(n8942) );
  inv_1 U7703 ( .ip(\CORTEXM0DS_INST/vis_ipsr [5]), .op(n9604) );
  nand3_1 U7704 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [4]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [3]), .ip3(n9604), .op(n11897) );
  nand3_1 U7705 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [2]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [1]), .ip3(\CORTEXM0DS_INST/vis_ipsr [0]), 
        .op(n11896) );
  nor2_1 U7706 ( .ip1(n11897), .ip2(n11896), .op(n6394) );
  inv_1 U7707 ( .ip(\CORTEXM0DS_INST/vis_ipsr [4]), .op(n11023) );
  nor3_1 U7708 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [5]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [3]), .ip3(n11023), .op(n6376) );
  inv_1 U7709 ( .ip(n6376), .op(n11880) );
  nor2_1 U7710 ( .ip1(n11880), .ip2(n11896), .op(n9113) );
  and2_1 U7711 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [15]), .ip2(n9113), .op(
        n6351) );
  inv_1 U7712 ( .ip(\CORTEXM0DS_INST/vis_ipsr [0]), .op(n11048) );
  nand3_1 U7713 ( .ip1(n11048), .ip2(\CORTEXM0DS_INST/vis_ipsr [1]), .ip3(
        \CORTEXM0DS_INST/vis_ipsr [2]), .op(n6360) );
  nand3_1 U7714 ( .ip1(n9604), .ip2(n11023), .ip3(
        \CORTEXM0DS_INST/vis_ipsr [3]), .op(n6370) );
  nor2_1 U7715 ( .ip1(n6360), .ip2(n6370), .op(n11892) );
  and2_1 U7716 ( .ip1(\CORTEXM0DS_INST/u_logic/Psh2z4 [1]), .ip2(n11892), .op(
        n6350) );
  not_ab_or_c_or_d U7717 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [31]), .ip2(
        n6394), .ip3(n6351), .ip4(n6350), .op(n6374) );
  nor2_1 U7718 ( .ip1(n6360), .ip2(n11897), .op(n9125) );
  inv_1 U7719 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [9]), .op(n8242) );
  inv_1 U7720 ( .ip(\CORTEXM0DS_INST/vis_ipsr [1]), .op(n11032) );
  nand4_1 U7721 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [2]), .ip2(n6376), .ip3(
        n11048), .ip4(n11032), .op(n10001) );
  nor2_1 U7722 ( .ip1(n8242), .ip2(n10001), .op(n6358) );
  nor4_1 U7723 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [2]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [0]), .ip3(n11032), .ip4(n11897), .op(n11890) );
  nand2_1 U7724 ( .ip1(n11890), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [21]), 
        .op(n6356) );
  nor4_1 U7725 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [2]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [0]), .ip3(n11032), .ip4(n11880), .op(n9119)
         );
  nand2_1 U7726 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [5]), .ip2(n9119), .op(
        n6355) );
  nor2_1 U7727 ( .ip1(n6370), .ip2(n11896), .op(n12049) );
  inv_1 U7728 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [11]), .op(n8243) );
  nand4_1 U7729 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [2]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [0]), .ip3(n6376), .ip4(n11032), .op(n9996)
         );
  nor2_1 U7730 ( .ip1(n8243), .ip2(n9996), .op(n6353) );
  nor3_1 U7731 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [2]), .ip2(n11032), .ip3(
        n11048), .op(n12402) );
  inv_1 U7732 ( .ip(n12402), .op(n11879) );
  nor2_1 U7733 ( .ip1(n11897), .ip2(n11879), .op(n6949) );
  and2_1 U7734 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [23]), .ip2(n6949), .op(
        n6352) );
  not_ab_or_c_or_d U7735 ( .ip1(\CORTEXM0DS_INST/u_logic/Txh2z4 [1]), .ip2(
        n12049), .ip3(n6353), .ip4(n6352), .op(n6354) );
  nand3_1 U7736 ( .ip1(n6356), .ip2(n6355), .ip3(n6354), .op(n6357) );
  not_ab_or_c_or_d U7737 ( .ip1(n9125), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [29]), .ip3(n6358), .ip4(n6357), .op(
        n6373) );
  nor4_1 U7738 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [0]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [1]), .ip3(n6359), .ip4(n11897), .op(n6383)
         );
  inv_1 U7739 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [27]), .op(n8336) );
  inv_1 U7740 ( .ip(n11897), .op(n6363) );
  nand4_1 U7741 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [2]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [0]), .ip3(n6363), .ip4(n11032), .op(n6952)
         );
  nor2_1 U7742 ( .ip1(n8336), .ip2(n6952), .op(n6362) );
  inv_1 U7743 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [13]), .op(n8232) );
  nor2_1 U7744 ( .ip1(n11880), .ip2(n6360), .op(n6398) );
  inv_1 U7745 ( .ip(n6398), .op(n11877) );
  nor2_1 U7746 ( .ip1(n8232), .ip2(n11877), .op(n6361) );
  not_ab_or_c_or_d U7747 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [25]), .ip2(
        n6383), .ip3(n6362), .ip4(n6361), .op(n6369) );
  nor4_1 U7748 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [2]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [1]), .ip3(n11048), .ip4(n11880), .op(n9131)
         );
  inv_1 U7749 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [1]), .op(n11858) );
  nand2_1 U7750 ( .ip1(n6377), .ip2(n6376), .op(n11876) );
  nor2_1 U7751 ( .ip1(n11858), .ip2(n11876), .op(n6365) );
  inv_1 U7752 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [17]), .op(n8197) );
  nand2_1 U7753 ( .ip1(n6377), .ip2(n6363), .op(n11891) );
  nor2_1 U7754 ( .ip1(n8197), .ip2(n11891), .op(n6364) );
  not_ab_or_c_or_d U7755 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [3]), .ip2(
        n9131), .ip3(n6365), .ip4(n6364), .op(n6368) );
  nor4_1 U7756 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [2]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [1]), .ip3(n11048), .ip4(n11897), .op(n6946)
         );
  nand2_1 U7757 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [19]), .ip2(n6946), 
        .op(n6367) );
  nor2_1 U7758 ( .ip1(n11880), .ip2(n11879), .op(n6375) );
  nand2_1 U7759 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [7]), .ip2(n6375), .op(
        n6366) );
  and4_1 U7760 ( .ip1(n6369), .ip2(n6368), .ip3(n6367), .ip4(n6366), .op(n6372) );
  nor2_1 U7761 ( .ip1(n6370), .ip2(n11879), .op(n11884) );
  nand2_1 U7762 ( .ip1(\CORTEXM0DS_INST/u_logic/Uth2z4 [1]), .ip2(n11884), 
        .op(n6371) );
  inv_1 U7763 ( .ip(\CORTEXM0DS_INST/u_logic/Uth2z4 [0]), .op(n8315) );
  nand2_1 U7764 ( .ip1(n6946), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [18]), 
        .op(n6401) );
  nand2_1 U7765 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [14]), .ip2(n9113), 
        .op(n6380) );
  nand2_1 U7766 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [6]), .ip2(n6375), .op(
        n6379) );
  nand3_1 U7767 ( .ip1(n6377), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [0]), 
        .ip3(n6376), .op(n6378) );
  nand3_1 U7768 ( .ip1(n6380), .ip2(n6379), .ip3(n6378), .op(n6393) );
  inv_1 U7769 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [16]), .op(n8196) );
  nor2_1 U7770 ( .ip1(n8196), .ip2(n11891), .op(n6382) );
  inv_1 U7771 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [8]), .op(n8237) );
  nor2_1 U7772 ( .ip1(n8237), .ip2(n10001), .op(n6381) );
  not_ab_or_c_or_d U7773 ( .ip1(n6949), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [22]), .ip3(n6382), .ip4(n6381), .op(
        n6391) );
  and2_1 U7774 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [4]), .ip2(n9119), .op(
        n6385) );
  inv_1 U7775 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [24]), .op(n8181) );
  inv_1 U7776 ( .ip(n6383), .op(n11878) );
  nor2_1 U7777 ( .ip1(n8181), .ip2(n11878), .op(n6384) );
  not_ab_or_c_or_d U7778 ( .ip1(n11890), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [20]), .ip3(n6385), .ip4(n6384), .op(
        n6390) );
  and2_1 U7779 ( .ip1(\CORTEXM0DS_INST/u_logic/Txh2z4 [0]), .ip2(n12049), .op(
        n6387) );
  and2_1 U7780 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [2]), .ip2(n9131), .op(
        n6386) );
  not_ab_or_c_or_d U7781 ( .ip1(n11892), .ip2(
        \CORTEXM0DS_INST/u_logic/Psh2z4 [0]), .ip3(n6387), .ip4(n6386), .op(
        n6389) );
  nand2_1 U7782 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [28]), .ip2(n9125), 
        .op(n6388) );
  not_ab_or_c_or_d U7783 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [30]), .ip2(
        n6394), .ip3(n6393), .ip4(n6392), .op(n6400) );
  inv_1 U7784 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [26]), .op(n8739) );
  nor2_1 U7785 ( .ip1(n8739), .ip2(n6952), .op(n6397) );
  inv_1 U7786 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [10]), .op(n6395) );
  nor2_1 U7787 ( .ip1(n6395), .ip2(n9996), .op(n6396) );
  not_ab_or_c_or_d U7788 ( .ip1(n6398), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [12]), .ip3(n6397), .ip4(n6396), .op(
        n6399) );
  nand3_1 U7789 ( .ip1(n6401), .ip2(n6400), .ip3(n6399), .op(n8924) );
  nand2_1 U7790 ( .ip1(n8315), .ip2(n8924), .op(n6403) );
  nand2_1 U7791 ( .ip1(\CORTEXM0DS_INST/u_logic/Uth2z4 [1]), .ip2(n6403), .op(
        n6405) );
  nor2_1 U7792 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [5]), .ip2(n11023), .op(n6402)
         );
  nor2_1 U7793 ( .ip1(\CORTEXM0DS_INST/u_logic/Uth2z4 [1]), .ip2(n6403), .op(
        n6404) );
  ab_or_c_or_d U7794 ( .ip1(n8934), .ip2(n6405), .ip3(n8937), .ip4(n6404), 
        .op(n6406) );
  inv_1 U7795 ( .ip(\CORTEXM0DS_INST/cm0_primask[0] ), .op(n11515) );
  nand3_1 U7796 ( .ip1(n8942), .ip2(n6406), .ip3(n11515), .op(n11703) );
  nand2_1 U7797 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n11796), .op(
        n10737) );
  nor2_1 U7798 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n10737), .op(
        n10662) );
  inv_1 U7799 ( .ip(n10662), .op(n11080) );
  nor3_1 U7800 ( .ip1(n11232), .ip2(n11080), .ip3(n6407), .op(n6413) );
  nor2_1 U7801 ( .ip1(n10492), .ip2(n12122), .op(n6408) );
  nor2_1 U7802 ( .ip1(n6409), .ip2(n6408), .op(n10777) );
  nor2_1 U7803 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Efgvx4 ), .op(n11249) );
  and4_1 U7804 ( .ip1(n11248), .ip2(n12369), .ip3(n11249), .ip4(n12125), .op(
        n11697) );
  nand3_1 U7805 ( .ip1(n6410), .ip2(n10777), .ip3(n11697), .op(n6411) );
  nand2_1 U7806 ( .ip1(n6420), .ip2(n6411), .op(n6412) );
  not_ab_or_c_or_d U7807 ( .ip1(n11684), .ip2(n11703), .ip3(n6413), .ip4(n6412), .op(n11688) );
  or2_1 U7808 ( .ip1(n11688), .ip2(n10743), .op(n6416) );
  or2_1 U7809 ( .ip1(n6414), .ip2(n10743), .op(n6415) );
  nand2_1 U7810 ( .ip1(n6416), .ip2(n6415), .op(n6417) );
  not_ab_or_c_or_d U7811 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n6419), 
        .ip3(n6418), .ip4(n6417), .op(n8065) );
  nand3_1 U7812 ( .ip1(n6420), .ip2(n8065), .ip3(n6945), .op(n7063) );
  nor2_1 U7813 ( .ip1(n6421), .ip2(n7063), .op(n10041) );
  or2_1 U7814 ( .ip1(n8916), .ip2(n10041), .op(n9140) );
  or2_1 U7815 ( .ip1(n11256), .ip2(n10530), .op(n6423) );
  or2_1 U7816 ( .ip1(n10737), .ip2(n10530), .op(n6422) );
  nand2_1 U7817 ( .ip1(n6423), .ip2(n6422), .op(n8917) );
  nor2_1 U7818 ( .ip1(n8917), .ip2(n9140), .op(n10017) );
  or2_1 U7819 ( .ip1(n11253), .ip2(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(
        n6425) );
  nand2_1 U7820 ( .ip1(n9946), .ip2(n12656), .op(n9892) );
  or2_1 U7821 ( .ip1(n9892), .ip2(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(n6424) );
  nand2_1 U7822 ( .ip1(n6425), .ip2(n6424), .op(n10054) );
  nor3_1 U7823 ( .ip1(n11228), .ip2(n11239), .ip3(n9402), .op(n6428) );
  nand2_1 U7824 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Vdgvx4 ), .op(n12070) );
  nor3_1 U7825 ( .ip1(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip3(n12070), .op(n6427) );
  nand2_1 U7826 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Vdgvx4 ), .op(n11241) );
  nor2_1 U7827 ( .ip1(n9943), .ip2(n11241), .op(n6426) );
  nor2_1 U7828 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .op(n11208) );
  inv_1 U7829 ( .ip(n11208), .op(n6429) );
  nand2_1 U7830 ( .ip1(n5639), .ip2(n12125), .op(n10740) );
  not_ab_or_c_or_d U7831 ( .ip1(n6429), .ip2(n11252), .ip3(n10851), .ip4(
        n10740), .op(n6434) );
  nor2_1 U7832 ( .ip1(n10852), .ip2(n6430), .op(n6433) );
  nand2_1 U7833 ( .ip1(n10762), .ip2(n6431), .op(n6432) );
  nand2_1 U7834 ( .ip1(n7079), .ip2(n6432), .op(n10052) );
  inv_1 U7835 ( .ip(n6435), .op(n11792) );
  nor3_1 U7836 ( .ip1(\CORTEXM0DS_INST/u_logic/Q5gvx4 ), .ip2(n11786), .ip3(
        n10972), .op(n9865) );
  nor3_1 U7837 ( .ip1(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip2(n10782), .ip3(
        n10739), .op(n10953) );
  not_ab_or_c_or_d U7838 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n11792), .ip3(n9865), .ip4(n10953), .op(n6436) );
  or2_1 U7839 ( .ip1(n6436), .ip2(n11693), .op(n6438) );
  nand2_1 U7840 ( .ip1(n10762), .ip2(n12125), .op(n6437) );
  inv_1 U7841 ( .ip(n12343), .op(n12605) );
  nor2_1 U7842 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n11796), .op(
        n6860) );
  nor2_1 U7843 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n12072), .op(
        n6789) );
  nand3_1 U7844 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n11065), .ip3(
        n9730), .op(n6442) );
  nand2_1 U7845 ( .ip1(n6442), .ip2(n6441), .op(n7438) );
  inv_1 U7846 ( .ip(n7438), .op(n12088) );
  inv_1 U7847 ( .ip(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .op(n11517) );
  nor2_1 U7848 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n11517), .op(
        n11160) );
  inv_1 U7849 ( .ip(\CORTEXM0DS_INST/u_logic/Tjh2z4 [1]), .op(n9091) );
  nand2_1 U7850 ( .ip1(n9091), .ip2(\CORTEXM0DS_INST/u_logic/Tjh2z4 [0]), .op(
        n6956) );
  nor3_1 U7851 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [2]), .ip2(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [3]), .ip3(n6956), .op(n6759) );
  nand2_1 U7852 ( .ip1(n6759), .ip2(\CORTEXM0DS_INST/cm0_r01 [31]), .op(n6447)
         );
  nor2_1 U7853 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [2]), .ip2(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [3]), .op(n6443) );
  and3_1 U7854 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [0]), .ip2(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [1]), .ip3(n6443), .op(n6762) );
  nand2_1 U7855 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [31]), .op(n6446)
         );
  inv_1 U7856 ( .ip(\CORTEXM0DS_INST/u_logic/Tjh2z4 [0]), .op(n11207) );
  nand2_1 U7857 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [1]), .ip2(n11207), 
        .op(n6880) );
  nor3_1 U7858 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [2]), .ip2(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [3]), .ip3(n6880), .op(n6771) );
  nand2_1 U7859 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [31]), .op(n6445)
         );
  inv_1 U7860 ( .ip(\CORTEXM0DS_INST/u_logic/Tjh2z4 [3]), .op(n9065) );
  nand2_1 U7861 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [2]), .ip2(n9065), .op(
        n6448) );
  nand2_1 U7862 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [0]), .ip2(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [1]), .op(n6882) );
  nor2_1 U7863 ( .ip1(n6448), .ip2(n6882), .op(n6764) );
  nand2_1 U7864 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [31]), .op(n6444)
         );
  or4_1 U7865 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [0]), .ip2(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [1]), .ip3(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [2]), .ip4(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [3]), .op(n6717) );
  inv_1 U7866 ( .ip(n6717), .op(n6760) );
  nand2_1 U7867 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [31]), .op(n6452)
         );
  nor2_1 U7868 ( .ip1(n6448), .ip2(n6956), .op(n6761) );
  nand2_1 U7869 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [31]), .op(n6451)
         );
  nor3_1 U7870 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [0]), .ip2(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [1]), .ip3(n6448), .op(n6772) );
  nand2_1 U7871 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [31]), .op(n6450)
         );
  nor2_1 U7872 ( .ip1(n6880), .ip2(n6448), .op(n6763) );
  nand2_1 U7873 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [31]), .op(n6449)
         );
  nor2_1 U7874 ( .ip1(n6454), .ip2(n6453), .op(n9349) );
  inv_1 U7875 ( .ip(n9349), .op(n8776) );
  and2_1 U7876 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [29]), .op(n6463)
         );
  nand2_1 U7877 ( .ip1(n6759), .ip2(\CORTEXM0DS_INST/cm0_r01 [29]), .op(n6461)
         );
  nand2_1 U7878 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [29]), .op(n6458)
         );
  nand2_1 U7879 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [29]), .op(n6457)
         );
  nand2_1 U7880 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [29]), .op(n6456)
         );
  nand2_1 U7881 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [29]), .op(n6455)
         );
  and4_1 U7882 ( .ip1(n6458), .ip2(n6457), .ip3(n6456), .ip4(n6455), .op(n6460) );
  nand2_1 U7883 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [29]), .op(n6459)
         );
  nand3_1 U7884 ( .ip1(n6461), .ip2(n6460), .ip3(n6459), .op(n6462) );
  not_ab_or_c_or_d U7885 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [29]), 
        .ip3(n6463), .ip4(n6462), .op(n8673) );
  nand2_1 U7886 ( .ip1(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Ml9vx4 ), .op(n11154) );
  nor2_1 U7887 ( .ip1(n8673), .ip2(n11154), .op(n6484) );
  and2_1 U7888 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [30]), .op(n6472)
         );
  nand2_1 U7889 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [30]), .ip2(n6759), .op(n6470)
         );
  nand2_1 U7890 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [30]), .op(n6467)
         );
  nand2_1 U7891 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [30]), .op(n6466)
         );
  nand2_1 U7892 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [30]), .op(n6465)
         );
  nand2_1 U7893 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [30]), .op(n6464)
         );
  and4_1 U7894 ( .ip1(n6467), .ip2(n6466), .ip3(n6465), .ip4(n6464), .op(n6469) );
  nand2_1 U7895 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [30]), .op(n6468)
         );
  nand3_1 U7896 ( .ip1(n6470), .ip2(n6469), .ip3(n6468), .op(n6471) );
  not_ab_or_c_or_d U7897 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [30]), .ip2(n6762), 
        .ip3(n6472), .ip4(n6471), .op(n9287) );
  and2_1 U7898 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [0]), .ip2(n6763), .op(n6481)
         );
  nand2_1 U7899 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [0]), .ip2(n6771), .op(n6479)
         );
  nand2_1 U7900 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [0]), .ip2(n6762), .op(n6476)
         );
  nand2_1 U7901 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [0]), .ip2(n6772), .op(n6475)
         );
  nand2_1 U7902 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [0]), .ip2(n6759), .op(n6474)
         );
  nand2_1 U7903 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [0]), .ip2(n6764), .op(n6473)
         );
  and4_1 U7904 ( .ip1(n6476), .ip2(n6475), .ip3(n6474), .ip4(n6473), .op(n6478) );
  nand2_1 U7905 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [0]), .ip2(n6761), .op(n6477)
         );
  nand3_1 U7906 ( .ip1(n6479), .ip2(n6478), .ip3(n6477), .op(n6480) );
  not_ab_or_c_or_d U7907 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [0]), 
        .ip3(n6481), .ip4(n6480), .op(n8797) );
  inv_1 U7908 ( .ip(n8797), .op(n8637) );
  nor2_1 U7909 ( .ip1(n8637), .ip2(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .op(
        n6482) );
  not_ab_or_c_or_d U7910 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n9287), 
        .ip3(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip4(n6482), .op(n6483) );
  not_ab_or_c_or_d U7911 ( .ip1(n11160), .ip2(n8776), .ip3(n6484), .ip4(n6483), 
        .op(n6525) );
  nand2_1 U7912 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [23]), .ip2(n6761), .op(n6493)
         );
  and2_1 U7913 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [23]), .op(n6490)
         );
  nand2_1 U7914 ( .ip1(n6759), .ip2(\CORTEXM0DS_INST/cm0_r01 [23]), .op(n6488)
         );
  nand2_1 U7915 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [23]), .op(n6487)
         );
  nand2_1 U7916 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [23]), .op(n6486)
         );
  nand2_1 U7917 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [23]), .op(n6485)
         );
  not_ab_or_c_or_d U7918 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [23]), .ip2(n6763), 
        .ip3(n6490), .ip4(n6489), .op(n6492) );
  nand2_1 U7919 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [23]), .op(n6491)
         );
  nand3_1 U7920 ( .ip1(n6493), .ip2(n6492), .ip3(n6491), .op(n9180) );
  and2_1 U7921 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [21]), .op(n6502)
         );
  nand2_1 U7922 ( .ip1(n6759), .ip2(\CORTEXM0DS_INST/cm0_r01 [21]), .op(n6500)
         );
  nand2_1 U7923 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [21]), .op(n6497)
         );
  nand2_1 U7924 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [21]), .op(n6496)
         );
  nand2_1 U7925 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [21]), .op(n6495)
         );
  nand2_1 U7926 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [21]), .op(n6494)
         );
  and4_1 U7927 ( .ip1(n6497), .ip2(n6496), .ip3(n6495), .ip4(n6494), .op(n6499) );
  nand2_1 U7928 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [21]), .op(n6498)
         );
  nand3_1 U7929 ( .ip1(n6500), .ip2(n6499), .ip3(n6498), .op(n6501) );
  not_ab_or_c_or_d U7930 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [21]), 
        .ip3(n6502), .ip4(n6501), .op(n8726) );
  nor2_1 U7931 ( .ip1(n8726), .ip2(n11154), .op(n6523) );
  and2_1 U7932 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [22]), .op(n6511)
         );
  nand2_1 U7933 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [22]), .op(n6509)
         );
  nand2_1 U7934 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [22]), .op(n6506)
         );
  nand2_1 U7935 ( .ip1(n6759), .ip2(\CORTEXM0DS_INST/cm0_r01 [22]), .op(n6505)
         );
  nand2_1 U7936 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [22]), .op(n6504)
         );
  nand2_1 U7937 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [22]), .op(n6503)
         );
  and4_1 U7938 ( .ip1(n6506), .ip2(n6505), .ip3(n6504), .ip4(n6503), .op(n6508) );
  nand2_1 U7939 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [22]), .op(n6507)
         );
  nand3_1 U7940 ( .ip1(n6509), .ip2(n6508), .ip3(n6507), .op(n6510) );
  not_ab_or_c_or_d U7941 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [22]), .ip2(n6772), 
        .ip3(n6511), .ip4(n6510), .op(n8129) );
  nand2_1 U7942 ( .ip1(n6759), .ip2(\CORTEXM0DS_INST/cm0_r01 [24]), .op(n6520)
         );
  and2_1 U7943 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [24]), .op(n6517)
         );
  nand2_1 U7944 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [24]), .op(n6515)
         );
  nand2_1 U7945 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [24]), .op(n6514)
         );
  nand2_1 U7946 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [24]), .op(n6513)
         );
  nand2_1 U7947 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [24]), .op(n6512)
         );
  not_ab_or_c_or_d U7948 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [24]), .ip2(n6764), 
        .ip3(n6517), .ip4(n6516), .op(n6519) );
  nand2_1 U7949 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [24]), .op(n6518)
         );
  nand3_1 U7950 ( .ip1(n6520), .ip2(n6519), .ip3(n6518), .op(n9178) );
  nor2_1 U7951 ( .ip1(n9178), .ip2(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .op(
        n6521) );
  not_ab_or_c_or_d U7952 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n8129), 
        .ip3(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip4(n6521), .op(n6522) );
  not_ab_or_c_or_d U7953 ( .ip1(n11160), .ip2(n9180), .ip3(n6523), .ip4(n6522), 
        .op(n6524) );
  mux2_1 U7954 ( .ip1(n6525), .ip2(n6524), .s(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .op(n6607) );
  nand2_1 U7955 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [27]), .ip2(n6759), .op(n6534)
         );
  and2_1 U7956 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [27]), .op(n6531)
         );
  nand2_1 U7957 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [27]), .op(n6529)
         );
  nand2_1 U7958 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [27]), .op(n6528)
         );
  nand2_1 U7959 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [27]), .op(n6527)
         );
  nand2_1 U7960 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [27]), .op(n6526)
         );
  not_ab_or_c_or_d U7961 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [27]), .ip2(n6764), 
        .ip3(n6531), .ip4(n6530), .op(n6533) );
  nand2_1 U7962 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [27]), .op(n6532)
         );
  nand3_1 U7963 ( .ip1(n6534), .ip2(n6533), .ip3(n6532), .op(n8768) );
  and2_1 U7964 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [25]), .op(n6543)
         );
  nand2_1 U7965 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [25]), .ip2(n6763), .op(n6541)
         );
  nand2_1 U7966 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [25]), .op(n6538)
         );
  nand2_1 U7967 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [25]), .op(n6537)
         );
  nand2_1 U7968 ( .ip1(n6759), .ip2(\CORTEXM0DS_INST/cm0_r01 [25]), .op(n6536)
         );
  nand2_1 U7969 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [25]), .op(n6535)
         );
  and4_1 U7970 ( .ip1(n6538), .ip2(n6537), .ip3(n6536), .ip4(n6535), .op(n6540) );
  nand2_1 U7971 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [25]), .op(n6539)
         );
  nand3_1 U7972 ( .ip1(n6541), .ip2(n6540), .ip3(n6539), .op(n6542) );
  not_ab_or_c_or_d U7973 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [25]), .ip2(n6772), 
        .ip3(n6543), .ip4(n6542), .op(n8426) );
  nor2_1 U7974 ( .ip1(n8426), .ip2(n11154), .op(n6564) );
  nand2_1 U7975 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [26]), .op(n6552)
         );
  and2_1 U7976 ( .ip1(n6759), .ip2(\CORTEXM0DS_INST/cm0_r01 [26]), .op(n6549)
         );
  nand2_1 U7977 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [26]), .op(n6547)
         );
  nand2_1 U7978 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [26]), .op(n6546)
         );
  nand2_1 U7979 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [26]), .op(n6545)
         );
  nand2_1 U7980 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [26]), .op(n6544)
         );
  not_ab_or_c_or_d U7981 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [26]), .ip2(n6760), 
        .ip3(n6549), .ip4(n6548), .op(n6551) );
  nand2_1 U7982 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [26]), .op(n6550)
         );
  nand3_1 U7983 ( .ip1(n6552), .ip2(n6551), .ip3(n6550), .op(n9184) );
  inv_1 U7984 ( .ip(n9184), .op(n8672) );
  and2_1 U7985 ( .ip1(n6759), .ip2(\CORTEXM0DS_INST/cm0_r01 [28]), .op(n6561)
         );
  nand2_1 U7986 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [28]), .ip2(n6764), .op(n6559)
         );
  nand2_1 U7987 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [28]), .op(n6556)
         );
  nand2_1 U7988 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [28]), .op(n6555)
         );
  nand2_1 U7989 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [28]), .op(n6554)
         );
  nand2_1 U7990 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [28]), .op(n6553)
         );
  and4_1 U7991 ( .ip1(n6556), .ip2(n6555), .ip3(n6554), .ip4(n6553), .op(n6558) );
  nand2_1 U7992 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [28]), .op(n6557)
         );
  nand3_1 U7993 ( .ip1(n6559), .ip2(n6558), .ip3(n6557), .op(n6560) );
  not_ab_or_c_or_d U7994 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [28]), .ip2(n6760), 
        .ip3(n6561), .ip4(n6560), .op(n8671) );
  inv_1 U7995 ( .ip(n8671), .op(n8774) );
  nor2_1 U7996 ( .ip1(n8774), .ip2(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .op(
        n6562) );
  not_ab_or_c_or_d U7997 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n8672), 
        .ip3(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip4(n6562), .op(n6563) );
  not_ab_or_c_or_d U7998 ( .ip1(n11160), .ip2(n8768), .ip3(n6564), .ip4(n6563), 
        .op(n6605) );
  nand2_1 U7999 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [19]), .ip2(n6761), .op(n6573)
         );
  and2_1 U8000 ( .ip1(n6759), .ip2(\CORTEXM0DS_INST/cm0_r01 [19]), .op(n6570)
         );
  nand2_1 U8001 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [19]), .op(n6568)
         );
  nand2_1 U8002 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [19]), .op(n6567)
         );
  nand2_1 U8003 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [19]), .op(n6566)
         );
  nand2_1 U8004 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [19]), .op(n6565)
         );
  not_ab_or_c_or_d U8005 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [19]), .ip2(n6760), 
        .ip3(n6570), .ip4(n6569), .op(n6572) );
  nand2_1 U8006 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [19]), .op(n6571)
         );
  nand3_1 U8007 ( .ip1(n6573), .ip2(n6572), .ip3(n6571), .op(n8824) );
  inv_1 U8008 ( .ip(\CORTEXM0DS_INST/cm0_r00 [17]), .op(n7787) );
  nor2_1 U8009 ( .ip1(n6717), .ip2(n7787), .op(n6582) );
  nand2_1 U8010 ( .ip1(n6759), .ip2(\CORTEXM0DS_INST/cm0_r01 [17]), .op(n6580)
         );
  nand2_1 U8011 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [17]), .op(n6577)
         );
  nand2_1 U8012 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [17]), .op(n6576)
         );
  nand2_1 U8013 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [17]), .op(n6575)
         );
  nand2_1 U8014 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [17]), .op(n6574)
         );
  and4_1 U8015 ( .ip1(n6577), .ip2(n6576), .ip3(n6575), .ip4(n6574), .op(n6579) );
  nand2_1 U8016 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [17]), .op(n6578)
         );
  nand3_1 U8017 ( .ip1(n6580), .ip2(n6579), .ip3(n6578), .op(n6581) );
  not_ab_or_c_or_d U8018 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [17]), 
        .ip3(n6582), .ip4(n6581), .op(n8408) );
  nor2_1 U8019 ( .ip1(n8408), .ip2(n11154), .op(n6603) );
  and2_1 U8020 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [18]), .ip2(n6760), .op(n6591)
         );
  nand2_1 U8021 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [18]), .ip2(n6764), .op(n6589)
         );
  nand2_1 U8022 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [18]), .ip2(n6771), .op(n6586)
         );
  nand2_1 U8023 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [18]), .ip2(n6761), .op(n6585)
         );
  nand2_1 U8024 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [18]), .ip2(n6762), .op(n6584)
         );
  nand2_1 U8025 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [18]), .ip2(n6772), .op(n6583)
         );
  and4_1 U8026 ( .ip1(n6586), .ip2(n6585), .ip3(n6584), .ip4(n6583), .op(n6588) );
  nand2_1 U8027 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [18]), .ip2(n6759), .op(n6587)
         );
  nand3_1 U8028 ( .ip1(n6589), .ip2(n6588), .ip3(n6587), .op(n6590) );
  not_ab_or_c_or_d U8029 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [18]), 
        .ip3(n6591), .ip4(n6590), .op(n8821) );
  nand2_1 U8030 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [20]), .ip2(n6759), .op(n6600)
         );
  and2_1 U8031 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [20]), .op(n6597)
         );
  nand2_1 U8032 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [20]), .op(n6595)
         );
  nand2_1 U8033 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [20]), .op(n6594)
         );
  nand2_1 U8034 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [20]), .op(n6593)
         );
  nand2_1 U8035 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [20]), .op(n6592)
         );
  not_ab_or_c_or_d U8036 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [20]), 
        .ip3(n6597), .ip4(n6596), .op(n6599) );
  nand2_1 U8037 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [20]), .op(n6598)
         );
  nand3_1 U8038 ( .ip1(n6600), .ip2(n6599), .ip3(n6598), .op(n8815) );
  nor2_1 U8039 ( .ip1(n8815), .ip2(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .op(
        n6601) );
  not_ab_or_c_or_d U8040 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n8821), 
        .ip3(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip4(n6601), .op(n6602) );
  not_ab_or_c_or_d U8041 ( .ip1(n11160), .ip2(n8824), .ip3(n6603), .ip4(n6602), 
        .op(n6604) );
  mux2_1 U8042 ( .ip1(n6605), .ip2(n6604), .s(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .op(n6606) );
  mux2_1 U8043 ( .ip1(n6607), .ip2(n6606), .s(\CORTEXM0DS_INST/u_logic/Qm9vx4 ), .op(n6784) );
  nor2_1 U8044 ( .ip1(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Ml9vx4 ), .op(n8112) );
  nand2_1 U8045 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [8]), .op(n6616)
         );
  and2_1 U8046 ( .ip1(n6759), .ip2(\CORTEXM0DS_INST/cm0_r01 [8]), .op(n6613)
         );
  nand2_1 U8047 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [8]), .op(n6611)
         );
  nand2_1 U8048 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [8]), .op(n6610)
         );
  nand2_1 U8049 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [8]), .op(n6609)
         );
  nand2_1 U8050 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [8]), .op(n6608)
         );
  not_ab_or_c_or_d U8051 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [8]), 
        .ip3(n6613), .ip4(n6612), .op(n6615) );
  nand2_1 U8052 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [8]), .op(n6614)
         );
  nand3_1 U8053 ( .ip1(n6616), .ip2(n6615), .ip3(n6614), .op(n9155) );
  nand2_1 U8054 ( .ip1(n8112), .ip2(n9155), .op(n6647) );
  inv_1 U8055 ( .ip(n11154), .op(n11079) );
  nand2_1 U8056 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [5]), .ip2(n6763), .op(n6625)
         );
  inv_1 U8057 ( .ip(\CORTEXM0DS_INST/cm0_r00 [5]), .op(n7482) );
  nor2_1 U8058 ( .ip1(n7482), .ip2(n6717), .op(n6622) );
  nand2_1 U8059 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [5]), .ip2(n6761), .op(n6620)
         );
  nand2_1 U8060 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [5]), .ip2(n6772), .op(n6619)
         );
  nand2_1 U8061 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [5]), .ip2(n6759), .op(n6618)
         );
  nand2_1 U8062 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [5]), .ip2(n6762), .op(n6617)
         );
  not_ab_or_c_or_d U8063 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [5]), 
        .ip3(n6622), .ip4(n6621), .op(n6624) );
  nand2_1 U8064 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [5]), .ip2(n6764), .op(n6623)
         );
  nand3_1 U8065 ( .ip1(n6625), .ip2(n6624), .ip3(n6623), .op(n8643) );
  nand2_1 U8066 ( .ip1(n11079), .ip2(n8643), .op(n6646) );
  nand2_1 U8067 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [7]), .ip2(n6764), .op(n6634)
         );
  inv_1 U8068 ( .ip(\CORTEXM0DS_INST/cm0_r00 [7]), .op(n7533) );
  nor2_1 U8069 ( .ip1(n7533), .ip2(n6717), .op(n6631) );
  nand2_1 U8070 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [7]), .ip2(n6771), .op(n6629)
         );
  nand2_1 U8071 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [7]), .ip2(n6759), .op(n6628)
         );
  nand2_1 U8072 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [7]), .ip2(n6761), .op(n6627)
         );
  nand2_1 U8073 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [7]), .ip2(n6762), .op(n6626)
         );
  not_ab_or_c_or_d U8074 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [7]), 
        .ip3(n6631), .ip4(n6630), .op(n6633) );
  nand2_1 U8075 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [7]), .ip2(n6763), .op(n6632)
         );
  nand3_1 U8076 ( .ip1(n6634), .ip2(n6633), .ip3(n6632), .op(n8698) );
  nand2_1 U8077 ( .ip1(n11160), .ip2(n8698), .op(n6645) );
  inv_1 U8078 ( .ip(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .op(n8069) );
  nor2_1 U8079 ( .ip1(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip2(n8069), .op(
        n6727) );
  nand2_1 U8080 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [6]), .ip2(n6760), .op(n6643)
         );
  and2_1 U8081 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [6]), .ip2(n6771), .op(n6640)
         );
  nand2_1 U8082 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [6]), .ip2(n6762), .op(n6638)
         );
  nand2_1 U8083 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [6]), .ip2(n6763), .op(n6637)
         );
  nand2_1 U8084 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [6]), .ip2(n6761), .op(n6636)
         );
  nand2_1 U8085 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [6]), .ip2(n6759), .op(n6635)
         );
  not_ab_or_c_or_d U8086 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [6]), 
        .ip3(n6640), .ip4(n6639), .op(n6642) );
  nand2_1 U8087 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [6]), .ip2(n6772), .op(n6641)
         );
  nand3_1 U8088 ( .ip1(n6643), .ip2(n6642), .ip3(n6641), .op(n8790) );
  nand2_1 U8089 ( .ip1(n6727), .ip2(n8790), .op(n6644) );
  nand2_1 U8090 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [15]), .ip2(n6760), .op(n6656)
         );
  and2_1 U8091 ( .ip1(n6759), .ip2(\CORTEXM0DS_INST/cm0_r01 [15]), .op(n6653)
         );
  nand2_1 U8092 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [15]), .op(n6651)
         );
  nand2_1 U8093 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [15]), .op(n6650)
         );
  nand2_1 U8094 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [15]), .op(n6649)
         );
  nand2_1 U8095 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [15]), .op(n6648)
         );
  not_ab_or_c_or_d U8096 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [15]), .ip2(n6761), 
        .ip3(n6653), .ip4(n6652), .op(n6655) );
  nand2_1 U8097 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [15]), .op(n6654)
         );
  nand3_1 U8098 ( .ip1(n6656), .ip2(n6655), .ip3(n6654), .op(n8718) );
  and2_1 U8099 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [13]), .op(n6665)
         );
  nand2_1 U8100 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [13]), .op(n6663)
         );
  nand2_1 U8101 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [13]), .op(n6660)
         );
  nand2_1 U8102 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [13]), .op(n6659)
         );
  nand2_1 U8103 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [13]), .op(n6658)
         );
  nand2_1 U8104 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [13]), .op(n6657)
         );
  and4_1 U8105 ( .ip1(n6660), .ip2(n6659), .ip3(n6658), .ip4(n6657), .op(n6662) );
  nand2_1 U8106 ( .ip1(n6759), .ip2(\CORTEXM0DS_INST/cm0_r01 [13]), .op(n6661)
         );
  nand3_1 U8107 ( .ip1(n6663), .ip2(n6662), .ip3(n6661), .op(n6664) );
  not_ab_or_c_or_d U8108 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [13]), 
        .ip3(n6665), .ip4(n6664), .op(n9149) );
  nor2_1 U8109 ( .ip1(n9149), .ip2(n11154), .op(n6686) );
  and2_1 U8110 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [14]), .op(n6674)
         );
  nand2_1 U8111 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [14]), .ip2(n6759), .op(n6672)
         );
  nand2_1 U8112 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [14]), .op(n6669)
         );
  nand2_1 U8113 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [14]), .op(n6668)
         );
  nand2_1 U8114 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [14]), .op(n6667)
         );
  nand2_1 U8115 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [14]), .op(n6666)
         );
  and4_1 U8116 ( .ip1(n6669), .ip2(n6668), .ip3(n6667), .ip4(n6666), .op(n6671) );
  nand2_1 U8117 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [14]), .op(n6670)
         );
  nand3_1 U8118 ( .ip1(n6672), .ip2(n6671), .ip3(n6670), .op(n6673) );
  not_ab_or_c_or_d U8119 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [14]), .ip2(n6762), 
        .ip3(n6674), .ip4(n6673), .op(n9147) );
  nand2_1 U8120 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [16]), .ip2(n6759), .op(n6683)
         );
  and2_1 U8121 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [16]), .op(n6680)
         );
  nand2_1 U8122 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [16]), .op(n6678)
         );
  nand2_1 U8123 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [16]), .op(n6677)
         );
  nand2_1 U8124 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [16]), .op(n6676)
         );
  nand2_1 U8125 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [16]), .op(n6675)
         );
  not_ab_or_c_or_d U8126 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [16]), 
        .ip3(n6680), .ip4(n6679), .op(n6682) );
  nand2_1 U8127 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [16]), .op(n6681)
         );
  nand3_1 U8128 ( .ip1(n6683), .ip2(n6682), .ip3(n6681), .op(n8822) );
  nor2_1 U8129 ( .ip1(n8822), .ip2(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .op(
        n6684) );
  not_ab_or_c_or_d U8130 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n9147), 
        .ip3(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip4(n6684), .op(n6685) );
  not_ab_or_c_or_d U8131 ( .ip1(n11160), .ip2(n8718), .ip3(n6686), .ip4(n6685), 
        .op(n6687) );
  nor2_1 U8132 ( .ip1(n6687), .ip2(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .op(
        n6688) );
  inv_1 U8133 ( .ip(\CORTEXM0DS_INST/u_logic/Qm9vx4 ), .op(n10942) );
  nand2_1 U8134 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(n10942), .op(
        n11516) );
  not_ab_or_c_or_d U8135 ( .ip1(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .ip2(n6689), 
        .ip3(n6688), .ip4(n11516), .op(n6783) );
  nand2_1 U8136 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [3]), .ip2(n6772), .op(n6698)
         );
  inv_1 U8137 ( .ip(\CORTEXM0DS_INST/cm0_r00 [3]), .op(n7032) );
  nor2_1 U8138 ( .ip1(n7032), .ip2(n6717), .op(n6695) );
  nand2_1 U8139 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [3]), .ip2(n6761), .op(n6693)
         );
  nand2_1 U8140 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [3]), .ip2(n6764), .op(n6692)
         );
  nand2_1 U8141 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [3]), .ip2(n6763), .op(n6691)
         );
  nand2_1 U8142 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [3]), .ip2(n6759), .op(n6690)
         );
  not_ab_or_c_or_d U8143 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [3]), 
        .ip3(n6695), .ip4(n6694), .op(n6697) );
  nand2_1 U8144 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [3]), .ip2(n6771), .op(n6696)
         );
  nand3_1 U8145 ( .ip1(n6698), .ip2(n6697), .ip3(n6696), .op(n8461) );
  nand2_1 U8146 ( .ip1(n11160), .ip2(n8461), .op(n6731) );
  nand2_1 U8147 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [1]), .ip2(n6761), .op(n6707)
         );
  inv_1 U8148 ( .ip(\CORTEXM0DS_INST/cm0_r00 [1]), .op(n6911) );
  nor2_1 U8149 ( .ip1(n6911), .ip2(n6717), .op(n6704) );
  nand2_1 U8150 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [1]), .ip2(n6762), .op(n6702)
         );
  nand2_1 U8151 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [1]), .ip2(n6759), .op(n6701)
         );
  nand2_1 U8152 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [1]), .ip2(n6763), .op(n6700)
         );
  nand2_1 U8153 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [1]), .ip2(n6771), .op(n6699)
         );
  not_ab_or_c_or_d U8154 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [1]), 
        .ip3(n6704), .ip4(n6703), .op(n6706) );
  nand2_1 U8155 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [1]), .ip2(n6772), .op(n6705)
         );
  nand3_1 U8156 ( .ip1(n6707), .ip2(n6706), .ip3(n6705), .op(n8638) );
  nand2_1 U8157 ( .ip1(n11079), .ip2(n8638), .op(n6730) );
  nand2_1 U8158 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [4]), .ip2(n6759), .op(n6716)
         );
  and2_1 U8159 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [4]), .ip2(n6761), .op(n6713)
         );
  nand2_1 U8160 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [4]), .ip2(n6771), .op(n6711)
         );
  nand2_1 U8161 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [4]), .ip2(n6760), .op(n6710)
         );
  nand2_1 U8162 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [4]), .ip2(n6762), .op(n6709)
         );
  nand2_1 U8163 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [4]), .ip2(n6772), .op(n6708)
         );
  not_ab_or_c_or_d U8164 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [4]), 
        .ip3(n6713), .ip4(n6712), .op(n6715) );
  nand2_1 U8165 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [4]), .ip2(n6763), .op(n6714)
         );
  nand3_1 U8166 ( .ip1(n6716), .ip2(n6715), .ip3(n6714), .op(n8462) );
  nand2_1 U8167 ( .ip1(n8112), .ip2(n8462), .op(n6729) );
  nand2_1 U8168 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [2]), .ip2(n6772), .op(n6726)
         );
  inv_1 U8169 ( .ip(\CORTEXM0DS_INST/cm0_r00 [2]), .op(n6994) );
  nor2_1 U8170 ( .ip1(n6994), .ip2(n6717), .op(n6723) );
  nand2_1 U8171 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [2]), .ip2(n6763), .op(n6721)
         );
  nand2_1 U8172 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [2]), .ip2(n6761), .op(n6720)
         );
  nand2_1 U8173 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [2]), .ip2(n6762), .op(n6719)
         );
  nand2_1 U8174 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [2]), .ip2(n6764), .op(n6718)
         );
  not_ab_or_c_or_d U8175 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [2]), 
        .ip3(n6723), .ip4(n6722), .op(n6725) );
  nand2_1 U8176 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [2]), .ip2(n6759), .op(n6724)
         );
  nand3_1 U8177 ( .ip1(n6726), .ip2(n6725), .ip3(n6724), .op(n8384) );
  nand2_1 U8178 ( .ip1(n6727), .ip2(n8384), .op(n6728) );
  nand2_1 U8179 ( .ip1(n6759), .ip2(\CORTEXM0DS_INST/cm0_r01 [11]), .op(n6740)
         );
  and2_1 U8180 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [11]), .op(n6737)
         );
  nand2_1 U8181 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [11]), .op(n6735)
         );
  nand2_1 U8182 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [11]), .op(n6734)
         );
  nand2_1 U8183 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [11]), .op(n6733)
         );
  nand2_1 U8184 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [11]), .op(n6732)
         );
  not_ab_or_c_or_d U8185 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [11]), .ip2(n6764), 
        .ip3(n6737), .ip4(n6736), .op(n6739) );
  nand2_1 U8186 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [11]), .op(n6738)
         );
  nand3_1 U8187 ( .ip1(n6740), .ip2(n6739), .ip3(n6738), .op(n8692) );
  and2_1 U8188 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [9]), .op(n6749)
         );
  nand2_1 U8189 ( .ip1(n6759), .ip2(\CORTEXM0DS_INST/cm0_r01 [9]), .op(n6747)
         );
  nand2_1 U8190 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [9]), .op(n6744)
         );
  nand2_1 U8191 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [9]), .op(n6743)
         );
  nand2_1 U8192 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [9]), .op(n6742)
         );
  nand2_1 U8193 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [9]), .op(n6741)
         );
  and4_1 U8194 ( .ip1(n6744), .ip2(n6743), .ip3(n6742), .ip4(n6741), .op(n6746) );
  nand2_1 U8195 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [9]), .op(n6745)
         );
  nand3_1 U8196 ( .ip1(n6747), .ip2(n6746), .ip3(n6745), .op(n6748) );
  not_ab_or_c_or_d U8197 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [9]), 
        .ip3(n6749), .ip4(n6748), .op(n9159) );
  nor2_1 U8198 ( .ip1(n9159), .ip2(n11154), .op(n6778) );
  nand2_1 U8199 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [10]), .op(n6756)
         );
  nand2_1 U8200 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [10]), .op(n6753)
         );
  nand2_1 U8201 ( .ip1(n6759), .ip2(\CORTEXM0DS_INST/cm0_r01 [10]), .op(n6752)
         );
  nand2_1 U8202 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [10]), .op(n6751)
         );
  nand2_1 U8203 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [10]), .op(n6750)
         );
  and4_1 U8204 ( .ip1(n6753), .ip2(n6752), .ip3(n6751), .ip4(n6750), .op(n6755) );
  nand2_1 U8205 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [10]), .op(n6754)
         );
  nand3_1 U8206 ( .ip1(n6756), .ip2(n6755), .ip3(n6754), .op(n6758) );
  and2_1 U8207 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [10]), .op(n6757)
         );
  not_ab_or_c_or_d U8208 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [10]), 
        .ip3(n6758), .ip4(n6757), .op(n9157) );
  nand2_1 U8209 ( .ip1(n6759), .ip2(\CORTEXM0DS_INST/cm0_r01 [12]), .op(n6775)
         );
  and2_1 U8210 ( .ip1(n6760), .ip2(\CORTEXM0DS_INST/cm0_r00 [12]), .op(n6770)
         );
  nand2_1 U8211 ( .ip1(n6761), .ip2(\CORTEXM0DS_INST/cm0_r05 [12]), .op(n6768)
         );
  nand2_1 U8212 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r03 [12]), .op(n6767)
         );
  nand2_1 U8213 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r06 [12]), .op(n6766)
         );
  nand2_1 U8214 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r07 [12]), .op(n6765)
         );
  not_ab_or_c_or_d U8215 ( .ip1(n6771), .ip2(\CORTEXM0DS_INST/cm0_r02 [12]), 
        .ip3(n6770), .ip4(n6769), .op(n6774) );
  nand2_1 U8216 ( .ip1(n6772), .ip2(\CORTEXM0DS_INST/cm0_r04 [12]), .op(n6773)
         );
  nand3_1 U8217 ( .ip1(n6775), .ip2(n6774), .ip3(n6773), .op(n8690) );
  nor2_1 U8218 ( .ip1(n8690), .ip2(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .op(
        n6776) );
  not_ab_or_c_or_d U8219 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n9157), 
        .ip3(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip4(n6776), .op(n6777) );
  not_ab_or_c_or_d U8220 ( .ip1(n11160), .ip2(n8692), .ip3(n6778), .ip4(n6777), 
        .op(n6779) );
  nor2_1 U8221 ( .ip1(n6779), .ip2(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .op(
        n6780) );
  nand2_1 U8222 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Qm9vx4 ), .op(n11810) );
  not_ab_or_c_or_d U8223 ( .ip1(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .ip2(n6781), 
        .ip3(n6780), .ip4(n11810), .op(n6782) );
  not_ab_or_c_or_d U8224 ( .ip1(n6784), .ip2(n12104), .ip3(n6783), .ip4(n6782), 
        .op(n6890) );
  nor2_1 U8225 ( .ip1(n12088), .ip2(n6890), .op(n9393) );
  nor3_1 U8226 ( .ip1(n12609), .ip2(n11228), .ip3(n11763), .op(n6787) );
  inv_1 U8227 ( .ip(n7017), .op(n9799) );
  nor2_1 U8228 ( .ip1(n9659), .ip2(n10478), .op(n10533) );
  nor3_1 U8229 ( .ip1(n9799), .ip2(n10533), .ip3(n10479), .op(n6785) );
  or4_1 U8230 ( .ip1(n9393), .ip2(n6787), .ip3(n6786), .ip4(n6785), .op(n6788)
         );
  not_ab_or_c_or_d U8231 ( .ip1(n11066), .ip2(n6860), .ip3(n6789), .ip4(n6788), 
        .op(n6790) );
  nor2_1 U8232 ( .ip1(n12605), .ip2(n6790), .op(n12316) );
  inv_1 U8233 ( .ip(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .op(n9807) );
  nor3_1 U8234 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip3(n9807), .op(n9754) );
  nand2_1 U8235 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .op(n11755) );
  nand2_1 U8236 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n11693), .op(
        n12131) );
  nor2_1 U8237 ( .ip1(n11755), .ip2(n12131), .op(n11257) );
  not_ab_or_c_or_d U8238 ( .ip1(n10813), .ip2(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip3(n9754), .ip4(n11257), .op(n6806) );
  inv_1 U8239 ( .ip(\CORTEXM0DS_INST/u_logic/O8gvx4 ), .op(n9797) );
  or2_1 U8240 ( .ip1(n6806), .ip2(n9797), .op(n6804) );
  nor2_1 U8241 ( .ip1(n9928), .ip2(n10479), .op(n10642) );
  or2_1 U8242 ( .ip1(\CORTEXM0DS_INST/vis_apsr [1]), .ip2(n10642), .op(n6794)
         );
  nand4_1 U8243 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip4(n11693), .op(n6791) );
  nand2_1 U8244 ( .ip1(n11253), .ip2(n6791), .op(n6792) );
  or2_1 U8245 ( .ip1(n6792), .ip2(n10642), .op(n6793) );
  nand2_1 U8246 ( .ip1(n6794), .ip2(n6793), .op(n6795) );
  nor2_1 U8247 ( .ip1(n6795), .ip2(n9807), .op(n6801) );
  nand2_1 U8248 ( .ip1(n9730), .ip2(n9853), .op(n6796) );
  or2_1 U8249 ( .ip1(n6796), .ip2(n11796), .op(n6799) );
  nand4_1 U8250 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip3(n11256), .ip4(n10421), .op(
        n6797) );
  or2_1 U8251 ( .ip1(n6797), .ip2(n11796), .op(n6798) );
  nand2_1 U8252 ( .ip1(n6799), .ip2(n6798), .op(n6800) );
  not_ab_or_c_or_d U8253 ( .ip1(n11256), .ip2(n12132), .ip3(n6801), .ip4(n6800), .op(n6802) );
  or2_1 U8254 ( .ip1(n6802), .ip2(n9797), .op(n6803) );
  nand2_1 U8255 ( .ip1(n6804), .ip2(n6803), .op(n6936) );
  nand2_1 U8256 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n11248), .op(
        n6805) );
  not_ab_or_c_or_d U8257 ( .ip1(n11253), .ip2(n6805), .ip3(n11228), .ip4(
        n12609), .op(n6810) );
  nor2_1 U8258 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n11765), .op(
        n6809) );
  nor2_1 U8259 ( .ip1(n12609), .ip2(n11786), .op(n9657) );
  nand2_1 U8260 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n11693), .op(
        n9382) );
  nor3_1 U8261 ( .ip1(n9657), .ip2(n11224), .ip3(n9382), .op(n6808) );
  inv_1 U8262 ( .ip(n6806), .op(n6807) );
  nor2_1 U8263 ( .ip1(n7106), .ip2(n9797), .op(n7940) );
  inv_1 U8264 ( .ip(n7940), .op(n7941) );
  nand2_1 U8265 ( .ip1(\CORTEXM0DS_INST/u_logic/Xq8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Fs8vx4 ), .op(n6825) );
  inv_1 U8266 ( .ip(\CORTEXM0DS_INST/u_logic/Nt8vx4 ), .op(n9037) );
  nand2_1 U8267 ( .ip1(n9037), .ip2(\CORTEXM0DS_INST/u_logic/Vu8vx4 ), .op(
        n6827) );
  nor2_1 U8268 ( .ip1(n6825), .ip2(n6827), .op(n9326) );
  inv_1 U8269 ( .ip(\CORTEXM0DS_INST/u_logic/Xq8vx4 ), .op(n11205) );
  nand2_1 U8270 ( .ip1(n11205), .ip2(\CORTEXM0DS_INST/u_logic/Fs8vx4 ), .op(
        n6826) );
  nor2_1 U8271 ( .ip1(n6826), .ip2(n6827), .op(n9335) );
  and2_1 U8272 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [0]), .op(n6833)
         );
  nand2_1 U8273 ( .ip1(\CORTEXM0DS_INST/u_logic/Vu8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nt8vx4 ), .op(n6824) );
  nor3_1 U8274 ( .ip1(\CORTEXM0DS_INST/u_logic/Xq8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Fs8vx4 ), .ip3(n6824), .op(n9317) );
  inv_1 U8275 ( .ip(\CORTEXM0DS_INST/u_logic/Fs8vx4 ), .op(n9010) );
  nand2_1 U8276 ( .ip1(n11205), .ip2(n9010), .op(n6811) );
  nor2_1 U8277 ( .ip1(n6811), .ip2(n6827), .op(n9334) );
  inv_1 U8278 ( .ip(n9334), .op(n7956) );
  inv_1 U8279 ( .ip(\CORTEXM0DS_INST/cm0_r08 [0]), .op(n6876) );
  nor2_1 U8280 ( .ip1(n7956), .ip2(n6876), .op(n6823) );
  inv_1 U8281 ( .ip(\CORTEXM0DS_INST/u_logic/Vu8vx4 ), .op(n9050) );
  nand2_1 U8282 ( .ip1(\CORTEXM0DS_INST/u_logic/Nt8vx4 ), .ip2(n9050), .op(
        n6813) );
  nor3_1 U8283 ( .ip1(\CORTEXM0DS_INST/u_logic/Xq8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Fs8vx4 ), .ip3(n6813), .op(n9318) );
  nand2_1 U8284 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [0]), .op(n6822)
         );
  nor2_1 U8285 ( .ip1(n6825), .ip2(n6813), .op(n9315) );
  nand2_1 U8286 ( .ip1(n9050), .ip2(n9037), .op(n6812) );
  or2_1 U8287 ( .ip1(n6812), .ip2(n6811), .op(n7788) );
  inv_1 U8288 ( .ip(n7788), .op(n9338) );
  and2_1 U8289 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [0]), .op(n6819)
         );
  nor3_1 U8290 ( .ip1(\CORTEXM0DS_INST/u_logic/Vu8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nt8vx4 ), .ip3(n6825), .op(n9344) );
  nand2_1 U8291 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [0]), .op(n6817)
         );
  nor3_1 U8292 ( .ip1(\CORTEXM0DS_INST/u_logic/Vu8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nt8vx4 ), .ip3(n6826), .op(n9316) );
  nand2_1 U8293 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [0]), .op(n6816)
         );
  nor2_1 U8294 ( .ip1(n6813), .ip2(n6826), .op(n9314) );
  nand2_1 U8295 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [0]), .op(n6815)
         );
  nand2_1 U8296 ( .ip1(n9010), .ip2(\CORTEXM0DS_INST/u_logic/Xq8vx4 ), .op(
        n6990) );
  nor2_1 U8297 ( .ip1(n6813), .ip2(n6990), .op(n9310) );
  nand2_1 U8298 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [0]), .op(n6814)
         );
  not_ab_or_c_or_d U8299 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [0]), .ip2(n9315), 
        .ip3(n6819), .ip4(n6818), .op(n6821) );
  nor3_1 U8300 ( .ip1(\CORTEXM0DS_INST/u_logic/Vu8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nt8vx4 ), .ip3(n6990), .op(n9308) );
  nand2_1 U8301 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [0]), .op(n6820)
         );
  nand3_1 U8302 ( .ip1(n6822), .ip2(n6821), .ip3(n6820), .op(n8075) );
  not_ab_or_c_or_d U8303 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [0]), 
        .ip3(n6823), .ip4(n8075), .op(n6831) );
  nor2_1 U8304 ( .ip1(n6825), .ip2(n6824), .op(n9325) );
  nand2_1 U8305 ( .ip1(n9325), .ip2(\CORTEXM0DS_INST/u_logic/Kycvx4 ), .op(
        n6830) );
  or3_1 U8306 ( .ip1(n9050), .ip2(n9037), .ip3(n6826), .op(n7857) );
  inv_1 U8307 ( .ip(n7857), .op(n9324) );
  nand2_1 U8308 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [0]), .op(n6829)
         );
  nor2_1 U8309 ( .ip1(n6990), .ip2(n6827), .op(n9309) );
  nand2_1 U8310 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [0]), .op(n6828)
         );
  not_ab_or_c_or_d U8311 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [0]), .ip2(n9326), 
        .ip3(n6833), .ip4(n6832), .op(n10058) );
  inv_1 U8312 ( .ip(n9382), .op(n9740) );
  nand2_1 U8313 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n12623), .op(
        n10945) );
  not_ab_or_c_or_d U8314 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n10945), .ip3(n12369), .ip4(n6834), .op(n6835) );
  nor2_1 U8315 ( .ip1(n6835), .ip2(n11796), .op(n6838) );
  nand2_1 U8316 ( .ip1(n12609), .ip2(n11796), .op(n10612) );
  nand2_1 U8317 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n12641), .op(
        n9772) );
  not_ab_or_c_or_d U8318 ( .ip1(n10612), .ip2(n9772), .ip3(n10698), .ip4(n8424), .op(n6837) );
  nor2_1 U8319 ( .ip1(n9377), .ip2(n10971), .op(n6836) );
  or2_1 U8320 ( .ip1(n6839), .ip2(n9797), .op(n6841) );
  nand2_1 U8321 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n9388), .op(
        n11754) );
  or2_1 U8322 ( .ip1(n11754), .ip2(n9797), .op(n6840) );
  nand2_1 U8323 ( .ip1(n6841), .ip2(n6840), .op(n7938) );
  inv_1 U8324 ( .ip(n7938), .op(n7887) );
  nor2_1 U8325 ( .ip1(n10058), .ip2(n7887), .op(n6851) );
  or2_1 U8326 ( .ip1(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip2(n6851), .op(n6853) );
  not_ab_or_c_or_d U8327 ( .ip1(n6842), .ip2(n11243), .ip3(n12117), .ip4(
        n12609), .op(n6847) );
  nor2_1 U8328 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Whgvx4 ), .op(n12133) );
  nor2_1 U8329 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n12117), .op(
        n9798) );
  nand2_1 U8330 ( .ip1(n9853), .ip2(n12609), .op(n6868) );
  or2_1 U8331 ( .ip1(n6868), .ip2(n9807), .op(n6843) );
  or2_1 U8332 ( .ip1(n10864), .ip2(n9807), .op(n9727) );
  nand2_1 U8333 ( .ip1(n6843), .ip2(n9727), .op(n6845) );
  nor2_1 U8334 ( .ip1(n11690), .ip2(n11241), .op(n6844) );
  ab_or_c_or_d U8335 ( .ip1(n12133), .ip2(n9798), .ip3(n6845), .ip4(n6844), 
        .op(n6846) );
  not_ab_or_c_or_d U8336 ( .ip1(n6860), .ip2(n11230), .ip3(n6847), .ip4(n6846), 
        .op(n6848) );
  nor2_1 U8337 ( .ip1(n6848), .ip2(n9797), .op(n7551) );
  inv_1 U8338 ( .ip(n7551), .op(n6850) );
  or4_1 U8339 ( .ip1(n9797), .ip2(n11755), .ip3(n11756), .ip4(
        \CORTEXM0DS_INST/u_logic/Whgvx4 ), .op(n6849) );
  nand2_1 U8340 ( .ip1(n6850), .ip2(n6849), .op(n7013) );
  or2_1 U8341 ( .ip1(n7013), .ip2(n6851), .op(n6852) );
  nand2_1 U8342 ( .ip1(n6853), .ip2(n6852), .op(n6854) );
  mux2_1 U8343 ( .ip1(n7941), .ip2(n7940), .s(n6854), .op(n9489) );
  nor3_1 U8344 ( .ip1(n11230), .ip2(n11267), .ip3(n11683), .op(n6855) );
  or2_1 U8345 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n6855), .op(n6858) );
  or2_1 U8346 ( .ip1(n6856), .ip2(n6855), .op(n6857) );
  nand2_1 U8347 ( .ip1(n6858), .ip2(n6857), .op(n6867) );
  or2_1 U8348 ( .ip1(n6859), .ip2(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(n6862) );
  inv_1 U8349 ( .ip(n6860), .op(n8961) );
  or2_1 U8350 ( .ip1(n8961), .ip2(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(n6861) );
  nand2_1 U8351 ( .ip1(n6862), .ip2(n6861), .op(n6865) );
  nand3_1 U8352 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip3(n8424), .op(n6863) );
  nand2_1 U8353 ( .ip1(n12641), .ip2(n12118), .op(n10919) );
  nand2_1 U8354 ( .ip1(n9657), .ip2(n12117), .op(n9724) );
  nand4_1 U8355 ( .ip1(\CORTEXM0DS_INST/u_logic/O8gvx4 ), .ip2(n6863), .ip3(
        n10919), .ip4(n9724), .op(n6864) );
  nand2_1 U8356 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [2]), .ip2(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [3]), .op(n6874) );
  inv_1 U8357 ( .ip(n6868), .op(n11217) );
  inv_1 U8358 ( .ip(n10945), .op(n9658) );
  nor3_1 U8359 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip3(n11756), .op(n12632) );
  nor3_1 U8360 ( .ip1(n9853), .ip2(n11208), .ip3(n12118), .op(n6869) );
  not_ab_or_c_or_d U8361 ( .ip1(n11217), .ip2(n9658), .ip3(n12632), .ip4(n6869), .op(n6873) );
  nand2_1 U8362 ( .ip1(n12619), .ip2(n10662), .op(n6872) );
  nand4_1 U8363 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [0]), .ip2(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [1]), .ip3(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [2]), .ip4(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [3]), .op(n6871) );
  or2_1 U8364 ( .ip1(n10612), .ip2(n12133), .op(n6870) );
  nor2_1 U8365 ( .ip1(n7438), .ip2(n6877), .op(n7437) );
  inv_1 U8366 ( .ip(n7437), .op(n9348) );
  or2_1 U8367 ( .ip1(n6874), .ip2(n9348), .op(n6955) );
  nor3_1 U8368 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [0]), .ip2(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [1]), .ip3(n6955), .op(n9365) );
  nand2_1 U8369 ( .ip1(n11207), .ip2(n9091), .op(n6875) );
  inv_1 U8370 ( .ip(\CORTEXM0DS_INST/u_logic/Tjh2z4 [2]), .op(n9102) );
  nand3_1 U8371 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [3]), .ip2(n7437), 
        .ip3(n9102), .op(n6881) );
  nor2_1 U8372 ( .ip1(n6875), .ip2(n6881), .op(n9354) );
  inv_1 U8373 ( .ip(n9354), .op(n7325) );
  nor2_1 U8374 ( .ip1(n7325), .ip2(n6876), .op(n6888) );
  nor2_1 U8375 ( .ip1(n6880), .ip2(n6881), .op(n9355) );
  nor2_1 U8376 ( .ip1(n8797), .ip2(n9348), .op(n6879) );
  nand2_1 U8377 ( .ip1(n6877), .ip2(n12088), .op(n7398) );
  inv_1 U8378 ( .ip(\CORTEXM0DS_INST/u_logic/Kycvx4 ), .op(n12328) );
  nor2_1 U8379 ( .ip1(n7398), .ip2(n12328), .op(n6878) );
  not_ab_or_c_or_d U8380 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [0]), .ip2(n9355), 
        .ip3(n6879), .ip4(n6878), .op(n6886) );
  or2_1 U8381 ( .ip1(n6880), .ip2(n6955), .op(n7423) );
  inv_1 U8382 ( .ip(n7423), .op(n9347) );
  nand2_1 U8383 ( .ip1(n9347), .ip2(\CORTEXM0DS_INST/cm0_r14 [0]), .op(n6885)
         );
  nor2_1 U8384 ( .ip1(n6956), .ip2(n6881), .op(n9364) );
  nand2_1 U8385 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [0]), .op(n6884)
         );
  nor2_1 U8386 ( .ip1(n6882), .ip2(n6881), .op(n9363) );
  nand2_1 U8387 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [0]), .op(n6883)
         );
  not_ab_or_c_or_d U8388 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [0]), .ip2(n9365), 
        .ip3(n6888), .ip4(n6887), .op(n9487) );
  nor2_1 U8389 ( .ip1(n9371), .ip2(n9487), .op(n6889) );
  xor2_1 U8390 ( .ip1(n9489), .ip2(n6889), .op(n6937) );
  xor2_1 U8391 ( .ip1(n6936), .ip2(n6937), .op(n11528) );
  inv_1 U8392 ( .ip(n11528), .op(n11060) );
  nand2_1 U8393 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n8424), .op(
        n11016) );
  nand2_1 U8394 ( .ip1(n11016), .ip2(n8961), .op(n6895) );
  nor3_1 U8395 ( .ip1(n12610), .ip2(n11208), .ip3(n11796), .op(n6894) );
  not_ab_or_c_or_d U8396 ( .ip1(n12633), .ip2(n11213), .ip3(n9799), .ip4(
        n11693), .op(n6892) );
  nand2_1 U8397 ( .ip1(n6890), .ip2(n7438), .op(n9379) );
  nand2_1 U8398 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n11250), .op(
        n6891) );
  not_ab_or_c_or_d U8399 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n6895), 
        .ip3(n6894), .ip4(n6893), .op(n6896) );
  nor2_1 U8400 ( .ip1(n12605), .ip2(n6896), .op(n12352) );
  inv_1 U8401 ( .ip(n12352), .op(n12311) );
  nor2_1 U8402 ( .ip1(n11060), .ip2(n12311), .op(n6897) );
  or2_1 U8403 ( .ip1(n12316), .ip2(n6897), .op(n6899) );
  inv_1 U8404 ( .ip(n9487), .op(n6931) );
  or2_1 U8405 ( .ip1(n6931), .ip2(n6897), .op(n6898) );
  nand2_1 U8406 ( .ip1(n6899), .ip2(n6898), .op(n10016) );
  nor2_1 U8407 ( .ip1(n10017), .ip2(n10016), .op(n6942) );
  or2_1 U8408 ( .ip1(n9140), .ip2(n6942), .op(n6944) );
  inv_1 U8409 ( .ip(\CORTEXM0DS_INST/cm0_r14 [1]), .op(n6910) );
  nor2_1 U8410 ( .ip1(n7423), .ip2(n6910), .op(n6909) );
  nand2_1 U8411 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [1]), .op(n6903)
         );
  nand2_1 U8412 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [1]), .op(n6902)
         );
  nand2_1 U8413 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [1]), .op(n6901)
         );
  nand2_1 U8414 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [1]), .op(n6900)
         );
  and4_1 U8415 ( .ip1(n6903), .ip2(n6902), .ip3(n6901), .ip4(n6900), .op(n6907) );
  nand2_1 U8416 ( .ip1(n7437), .ip2(n8638), .op(n6906) );
  nand2_1 U8417 ( .ip1(\CORTEXM0DS_INST/u_logic/Kycvx4 ), .ip2(n7438), .op(
        n6905) );
  inv_1 U8418 ( .ip(n7398), .op(n9353) );
  nand2_1 U8419 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/Uzcvx4 ), .op(
        n6904) );
  ab_or_c_or_d U8420 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [1]), .ip2(n9363), .ip3(
        n6909), .ip4(n6908), .op(n9505) );
  nand2_1 U8421 ( .ip1(n9505), .ip2(n12316), .op(n6941) );
  nor2_1 U8422 ( .ip1(n7857), .ip2(n6910), .op(n6927) );
  and2_1 U8423 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [1]), .op(n6921)
         );
  nand2_1 U8424 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [1]), .op(n6920)
         );
  nor2_1 U8425 ( .ip1(n7788), .ip2(n6911), .op(n6917) );
  nand2_1 U8426 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [1]), .op(n6915)
         );
  nand2_1 U8427 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [1]), .op(n6914)
         );
  nand2_1 U8428 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [1]), .op(n6913)
         );
  nand2_1 U8429 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [1]), .op(n6912)
         );
  not_ab_or_c_or_d U8430 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [1]), 
        .ip3(n6917), .ip4(n6916), .op(n6919) );
  nand2_1 U8431 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [1]), .op(n6918)
         );
  nand3_1 U8432 ( .ip1(n6920), .ip2(n6919), .ip3(n6918), .op(n8071) );
  not_ab_or_c_or_d U8433 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [1]), 
        .ip3(n6921), .ip4(n8071), .op(n6925) );
  nand2_1 U8434 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [1]), .op(n6924)
         );
  nand2_1 U8435 ( .ip1(n9325), .ip2(\CORTEXM0DS_INST/u_logic/Uzcvx4 ), .op(
        n6923) );
  nand2_1 U8436 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [1]), .op(n6922)
         );
  not_ab_or_c_or_d U8437 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [1]), .ip2(n9317), 
        .ip3(n6927), .ip4(n6926), .op(n11807) );
  nor2_1 U8438 ( .ip1(n11807), .ip2(n7887), .op(n6929) );
  nor3_1 U8439 ( .ip1(n9797), .ip2(n11241), .ip3(n11240), .op(n7889) );
  inv_1 U8440 ( .ip(n7889), .op(n7935) );
  inv_1 U8441 ( .ip(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), .op(n12542) );
  nor2_1 U8442 ( .ip1(n7935), .ip2(n12542), .op(n6928) );
  not_ab_or_c_or_d U8443 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n7013), 
        .ip3(n6929), .ip4(n6928), .op(n6930) );
  mux2_1 U8444 ( .ip1(n7941), .ip2(n7940), .s(n6930), .op(n9504) );
  nand2_1 U8445 ( .ip1(n9261), .ip2(n9505), .op(n6933) );
  and2_1 U8446 ( .ip1(n6931), .ip2(n9489), .op(n9493) );
  nand2_1 U8447 ( .ip1(n9493), .ip2(n9261), .op(n6932) );
  nand2_1 U8448 ( .ip1(n6933), .ip2(n6932), .op(n6987) );
  inv_1 U8449 ( .ip(n6933), .op(n6934) );
  nand2_1 U8450 ( .ip1(n9493), .ip2(n6934), .op(n6989) );
  nand2_1 U8451 ( .ip1(n6987), .ip2(n6989), .op(n6935) );
  xor2_1 U8452 ( .ip1(n9504), .ip2(n6935), .op(n7056) );
  nand2_1 U8453 ( .ip1(n6937), .ip2(n6936), .op(n7055) );
  xor2_1 U8454 ( .ip1(n7056), .ip2(n7055), .op(n10915) );
  nand2_1 U8455 ( .ip1(n10915), .ip2(n12352), .op(n6940) );
  inv_1 U8456 ( .ip(n12645), .op(n12112) );
  nand2_1 U8457 ( .ip1(n12112), .ip2(\CORTEXM0DS_INST/vis_pc [0]), .op(n6970)
         );
  inv_1 U8458 ( .ip(\CORTEXM0DS_INST/vis_pc [0]), .op(n8629) );
  nand2_1 U8459 ( .ip1(n12645), .ip2(n8629), .op(n6938) );
  nand3_1 U8460 ( .ip1(n12605), .ip2(n6970), .ip3(n6938), .op(n6939) );
  nand3_1 U8461 ( .ip1(n6941), .ip2(n6940), .ip3(n6939), .op(n11201) );
  or2_1 U8462 ( .ip1(n11201), .ip2(n6942), .op(n6943) );
  nand2_1 U8463 ( .ip1(n6944), .ip2(n6943), .op(n12606) );
  nor2_1 U8464 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n5639), .op(
        n9385) );
  inv_1 U8465 ( .ip(n9385), .op(n11242) );
  nand3_1 U8466 ( .ip1(n10556), .ip2(n11228), .ip3(n12125), .op(n11895) );
  inv_1 U8467 ( .ip(n11895), .op(n3276) );
  and2_1 U8468 ( .ip1(n6946), .ip2(n3276), .op(n6948) );
  inv_1 U8469 ( .ip(\CORTEXM0DS_INST/u_logic/Z7hvx4 ), .op(n9146) );
  nand2_1 U8470 ( .ip1(\CORTEXM0DS_INST/u_logic/B5hvx4 ), .ip2(n9146), .op(
        n8337) );
  nor2_1 U8471 ( .ip1(\CORTEXM0DS_INST/u_logic/L9hvx4 ), .ip2(n8337), .op(
        n11903) );
  inv_1 U8472 ( .ip(\CORTEXM0DS_INST/u_logic/Xahvx4 ), .op(n11898) );
  nand2_1 U8473 ( .ip1(\CORTEXM0DS_INST/u_logic/N6hvx4 ), .ip2(n11898), .op(
        n8659) );
  inv_1 U8474 ( .ip(n8659), .op(n8658) );
  nand3_1 U8475 ( .ip1(n11903), .ip2(n8658), .ip3(
        \CORTEXM0DS_INST/u_logic/Mf8vx4 ), .op(n11705) );
  inv_1 U8476 ( .ip(n11705), .op(n9919) );
  nor2_1 U8477 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [9]), .ip2(n9919), .op(
        n6947) );
  nor4_1 U8478 ( .ip1(n6948), .ip2(n2528), .ip3(n12738), .ip4(n6947), .op(
        \CORTEXM0DS_INST/u_logic/I0ivx4 ) );
  and2_1 U8479 ( .ip1(n6949), .ip2(n3276), .op(n6951) );
  nor2_1 U8480 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [11]), .ip2(n9919), .op(
        n6950) );
  nor4_1 U8481 ( .ip1(n6951), .ip2(n2531), .ip3(n12737), .ip4(n6950), .op(
        \CORTEXM0DS_INST/u_logic/Uzhvx4 ) );
  nor2_1 U8482 ( .ip1(n6952), .ip2(n11895), .op(n6954) );
  nor2_1 U8483 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [13]), .ip2(n9919), .op(
        n6953) );
  nor4_1 U8484 ( .ip1(n6954), .ip2(n2502), .ip3(n12740), .ip4(n6953), .op(
        \CORTEXM0DS_INST/u_logic/Gzhvx4 ) );
  and2_1 U8485 ( .ip1(n9347), .ip2(\CORTEXM0DS_INST/cm0_r14 [3]), .op(n6969)
         );
  and2_1 U8486 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [3]), .op(n6962)
         );
  inv_1 U8487 ( .ip(\CORTEXM0DS_INST/u_logic/O7evx4 ), .op(n11571) );
  or2_1 U8488 ( .ip1(n6956), .ip2(n6955), .op(n6963) );
  nor2_1 U8489 ( .ip1(n11571), .ip2(n6963), .op(n9356) );
  nand2_1 U8490 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [1]), .op(n6960)
         );
  nand2_1 U8491 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/O2dvx4 ), .op(
        n6959) );
  nand2_1 U8492 ( .ip1(\CORTEXM0DS_INST/u_logic/E1dvx4 ), .ip2(n7438), .op(
        n6958) );
  nand2_1 U8493 ( .ip1(n7437), .ip2(n8461), .op(n6957) );
  not_ab_or_c_or_d U8494 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [3]), .ip2(n9364), 
        .ip3(n6962), .ip4(n6961), .op(n6967) );
  nand2_1 U8495 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [3]), .op(n6966)
         );
  nand2_1 U8496 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [3]), .op(n6965)
         );
  nor2_1 U8497 ( .ip1(\CORTEXM0DS_INST/u_logic/O7evx4 ), .ip2(n6963), .op(
        n9366) );
  nand2_1 U8498 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [1]), .op(n6964)
         );
  not_ab_or_c_or_d U8499 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [3]), .ip2(n9355), 
        .ip3(n6969), .ip4(n6968), .op(n9486) );
  inv_1 U8500 ( .ip(n9486), .op(n7061) );
  inv_1 U8501 ( .ip(\CORTEXM0DS_INST/u_logic/I4gvx4 ), .op(n7062) );
  nor2_1 U8502 ( .ip1(n7062), .ip2(n6970), .op(n6972) );
  mux2_1 U8503 ( .ip1(\CORTEXM0DS_INST/u_logic/I4gvx4 ), .ip2(n6971), .s(n6970), .op(n8858) );
  inv_1 U8504 ( .ip(\CORTEXM0DS_INST/vis_pc [1]), .op(n12401) );
  nor2_1 U8505 ( .ip1(n8858), .ip2(n12401), .op(n8857) );
  nor2_1 U8506 ( .ip1(n6972), .ip2(n8857), .op(n6973) );
  nor2_1 U8507 ( .ip1(n6973), .ip2(n8587), .op(n8871) );
  not_ab_or_c_or_d U8508 ( .ip1(n6973), .ip2(n8587), .ip3(n8871), .ip4(n12343), 
        .op(n7060) );
  nor2_1 U8509 ( .ip1(n9371), .ip2(n9486), .op(n7452) );
  nor2_1 U8510 ( .ip1(n9797), .ip2(n12118), .op(n6986) );
  nor2_1 U8511 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n11793), .op(
        n9833) );
  and2_1 U8512 ( .ip1(n9347), .ip2(\CORTEXM0DS_INST/cm0_r14 [2]), .op(n6985)
         );
  inv_1 U8513 ( .ip(n9355), .op(n7436) );
  inv_1 U8514 ( .ip(\CORTEXM0DS_INST/cm0_r10 [2]), .op(n6991) );
  nor2_1 U8515 ( .ip1(n7436), .ip2(n6991), .op(n6979) );
  nand2_1 U8516 ( .ip1(n7437), .ip2(n8384), .op(n6977) );
  nand2_1 U8517 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/E1dvx4 ), .op(
        n6976) );
  nand2_1 U8518 ( .ip1(\CORTEXM0DS_INST/u_logic/Uzcvx4 ), .ip2(n7438), .op(
        n6975) );
  nand2_1 U8519 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [0]), .op(n6974)
         );
  not_ab_or_c_or_d U8520 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [2]), .ip2(n9365), 
        .ip3(n6979), .ip4(n6978), .op(n6983) );
  nand2_1 U8521 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [2]), .op(n6982)
         );
  nand2_1 U8522 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [2]), .op(n6981)
         );
  nand2_1 U8523 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [0]), .op(n6980)
         );
  not_ab_or_c_or_d U8524 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [2]), .ip2(n9364), 
        .ip3(n6985), .ip4(n6984), .op(n11760) );
  not_ab_or_c_or_d U8525 ( .ip1(n6986), .ip2(n9833), .ip3(n9371), .ip4(n11760), 
        .op(n7058) );
  nand2_1 U8526 ( .ip1(n6987), .ip2(n9504), .op(n6988) );
  nand2_1 U8527 ( .ip1(n6989), .ip2(n6988), .op(n7057) );
  or3_1 U8528 ( .ip1(n9050), .ip2(n9037), .ip3(n6990), .op(n7008) );
  nor2_1 U8529 ( .ip1(n7008), .ip2(n11571), .op(n9323) );
  inv_1 U8530 ( .ip(n9335), .op(n7585) );
  nor2_1 U8531 ( .ip1(n7585), .ip2(n6991), .op(n6993) );
  and2_1 U8532 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [2]), .op(n6992)
         );
  not_ab_or_c_or_d U8533 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [0]), 
        .ip3(n6993), .ip4(n6992), .op(n7012) );
  nand2_1 U8534 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [2]), .op(n7003)
         );
  nor2_1 U8535 ( .ip1(n7788), .ip2(n6994), .op(n7000) );
  nand2_1 U8536 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [2]), .op(n6998)
         );
  nand2_1 U8537 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [2]), .op(n6997)
         );
  nand2_1 U8538 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [2]), .op(n6996)
         );
  nand2_1 U8539 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [2]), .op(n6995)
         );
  not_ab_or_c_or_d U8540 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [2]), .ip2(n9308), 
        .ip3(n7000), .ip4(n6999), .op(n7002) );
  nand2_1 U8541 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [2]), .op(n7001)
         );
  nand3_1 U8542 ( .ip1(n7003), .ip2(n7002), .ip3(n7001), .op(n8090) );
  nand2_1 U8543 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [2]), .op(n7006)
         );
  nand2_1 U8544 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [2]), .op(n7005)
         );
  nand2_1 U8545 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [2]), .op(n7004)
         );
  nand3_1 U8546 ( .ip1(n7006), .ip2(n7005), .ip3(n7004), .op(n7007) );
  not_ab_or_c_or_d U8547 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [2]), .ip2(n9317), 
        .ip3(n8090), .ip4(n7007), .op(n7011) );
  nor2_1 U8548 ( .ip1(\CORTEXM0DS_INST/u_logic/O7evx4 ), .ip2(n7008), .op(
        n9333) );
  nand2_1 U8549 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [0]), .op(n7010)
         );
  nand2_1 U8550 ( .ip1(n9325), .ip2(\CORTEXM0DS_INST/u_logic/E1dvx4 ), .op(
        n7009) );
  nand2_1 U8551 ( .ip1(n7938), .ip2(n12671), .op(n7028) );
  nand2_1 U8552 ( .ip1(\CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip2(n7013), .op(
        n7027) );
  nand2_1 U8553 ( .ip1(n7889), .ip2(\CORTEXM0DS_INST/u_logic/B19vx4 ), .op(
        n7026) );
  inv_1 U8554 ( .ip(n9657), .op(n8494) );
  not_ab_or_c_or_d U8555 ( .ip1(n9658), .ip2(n8424), .ip3(n9853), .ip4(n11223), 
        .op(n7015) );
  or2_1 U8556 ( .ip1(n7524), .ip2(n9797), .op(n7024) );
  not_ab_or_c_or_d U8557 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n12627), .ip3(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip4(n11228), .op(n7021) );
  nand2_1 U8558 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n8424), .op(
        n9956) );
  nand2_1 U8559 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(n9807), .op(
        n9957) );
  not_ab_or_c_or_d U8560 ( .ip1(n9815), .ip2(n9956), .ip3(n8358), .ip4(n9957), 
        .op(n7020) );
  nor2_1 U8561 ( .ip1(n12118), .ip2(n10971), .op(n7019) );
  nor2_1 U8562 ( .ip1(n11682), .ip2(n7017), .op(n7018) );
  or2_1 U8563 ( .ip1(n7022), .ip2(n9797), .op(n7023) );
  nand2_1 U8564 ( .ip1(n7024), .ip2(n7023), .op(n7478) );
  nand2_1 U8565 ( .ip1(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip2(n7478), .op(
        n7025) );
  mux2_1 U8566 ( .ip1(n7940), .ip2(n7941), .s(n7029), .op(n9453) );
  and2_1 U8567 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [3]), .op(n7031)
         );
  and2_1 U8568 ( .ip1(n9325), .ip2(\CORTEXM0DS_INST/u_logic/O2dvx4 ), .op(
        n7030) );
  not_ab_or_c_or_d U8569 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [1]), 
        .ip3(n7031), .ip4(n7030), .op(n7049) );
  nand2_1 U8570 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [3]), .ip2(n9318), .op(n7041)
         );
  nor2_1 U8571 ( .ip1(n7788), .ip2(n7032), .op(n7038) );
  nand2_1 U8572 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [3]), .op(n7036)
         );
  nand2_1 U8573 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [3]), .op(n7035)
         );
  nand2_1 U8574 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [3]), .op(n7034)
         );
  nand2_1 U8575 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [3]), .op(n7033)
         );
  not_ab_or_c_or_d U8576 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [3]), 
        .ip3(n7038), .ip4(n7037), .op(n7040) );
  nand2_1 U8577 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [3]), .op(n7039)
         );
  nand3_1 U8578 ( .ip1(n7041), .ip2(n7040), .ip3(n7039), .op(n8108) );
  nand2_1 U8579 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [3]), .ip2(n9334), .op(n7044)
         );
  nand2_1 U8580 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [3]), .op(n7043)
         );
  nand2_1 U8581 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [3]), .op(n7042)
         );
  nand3_1 U8582 ( .ip1(n7044), .ip2(n7043), .ip3(n7042), .op(n7045) );
  not_ab_or_c_or_d U8583 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [3]), .ip2(n9317), 
        .ip3(n8108), .ip4(n7045), .op(n7048) );
  nand2_1 U8584 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [1]), .op(n7047)
         );
  nand2_1 U8585 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [3]), .op(n7046)
         );
  nand2_1 U8586 ( .ip1(n7938), .ip2(n12677), .op(n7053) );
  nand2_1 U8587 ( .ip1(n7889), .ip2(\CORTEXM0DS_INST/u_logic/I29vx4 ), .op(
        n7052) );
  nand2_1 U8588 ( .ip1(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .ip2(n7551), .op(
        n7051) );
  nand2_1 U8589 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n7478), .op(
        n7050) );
  mux2_1 U8590 ( .ip1(n7940), .ip2(n7941), .s(n7054), .op(n9481) );
  nor2_1 U8591 ( .ip1(n7056), .ip2(n7055), .op(n8856) );
  fulladder U8592 ( .a(n7058), .b(n7057), .ci(n9453), .co(n7451), .s(n8855) );
  nand2_1 U8593 ( .ip1(n8856), .ip2(n8855), .op(n8036) );
  xor2_1 U8594 ( .ip1(n8035), .ip2(n8036), .op(n9415) );
  nor2_1 U8595 ( .ip1(n9415), .ip2(n12311), .op(n7059) );
  not_ab_or_c_or_d U8596 ( .ip1(n12316), .ip2(n7061), .ip3(n7060), .ip4(n7059), 
        .op(\CORTEXM0DS_INST/u_logic/Ekovx4 ) );
  inv_1 U8597 ( .ip(n1185), .op(n12536) );
  nand3_1 U8598 ( .ip1(n12112), .ip2(n7062), .ip3(n12536), .op(n7064) );
  inv_1 U8599 ( .ip(n12111), .op(n12647) );
  not_ab_or_c_or_d U8600 ( .ip1(n1708), .ip2(n7064), .ip3(n12647), .ip4(n7063), 
        .op(n12600) );
  nand2_1 U8601 ( .ip1(n12600), .ip2(\CORTEXM0DS_INST/u_logic/V8evx4 ), .op(
        n12593) );
  inv_1 U8602 ( .ip(n12593), .op(n12598) );
  nor3_1 U8603 ( .ip1(\interconnect_ip_inst/i_ahb_U_mux_hsel_prev [4]), .ip2(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [3]), .ip3(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [2]), .op(n7065) );
  and2_1 U8604 ( .ip1(n7065), .ip2(n449), .op(n12608) );
  inv_1 U8605 ( .ip(\CORTEXM0DS_INST/cm0_xpsr[24] ), .op(n11071) );
  nor3_1 U8606 ( .ip1(n12608), .ip2(\CORTEXM0DS_INST/u_logic/H0gvx4 ), .ip3(
        n11071), .op(n9105) );
  inv_1 U8607 ( .ip(n9105), .op(n12660) );
  nand2_1 U8608 ( .ip1(n7065), .ip2(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [1]), .op(n9986) );
  nor2_1 U8609 ( .ip1(n12660), .ip2(n9986), .op(n4807) );
  inv_1 U8610 ( .ip(n4807), .op(n12535) );
  inv_1 U8611 ( .ip(n12600), .op(n12575) );
  nor4_1 U8612 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n8629), .ip3(
        n12535), .ip4(n12575), .op(n1143) );
  inv_1 U8613 ( .ip(n1143), .op(n12577) );
  nor2_1 U8614 ( .ip1(n1154), .ip2(n12577), .op(n7066) );
  or2_1 U8615 ( .ip1(n12598), .ip2(n7066), .op(n7068) );
  or2_1 U8616 ( .ip1(\CORTEXM0DS_INST/u_logic/G8fvx4 ), .ip2(n7066), .op(n7067) );
  nand2_1 U8617 ( .ip1(n7068), .ip2(n7067), .op(n7072) );
  or2_1 U8618 ( .ip1(\CORTEXM0DS_INST/u_logic/V8evx4 ), .ip2(n8629), .op(n7069) );
  not_ab_or_c_or_d U8619 ( .ip1(n12112), .ip2(n7069), .ip3(
        \CORTEXM0DS_INST/u_logic/Xyfvx4 ), .ip4(n12575), .op(n12603) );
  nand2_1 U8620 ( .ip1(n12603), .ip2(\CORTEXM0DS_INST/u_logic/Bwfvx4 ), .op(
        n7071) );
  nand2_1 U8621 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(n12575), .op(
        n7070) );
  nand4_1 U8622 ( .ip1(n1153), .ip2(n7072), .ip3(n7071), .ip4(n7070), .op(
        n6025) );
  inv_1 U8623 ( .ip(\CORTEXM0DS_INST/u_logic/W49vx4 ), .op(n9881) );
  nor2_1 U8624 ( .ip1(n12600), .ip2(n9881), .op(n7073) );
  or2_1 U8625 ( .ip1(n12598), .ip2(n7073), .op(n7075) );
  or2_1 U8626 ( .ip1(\CORTEXM0DS_INST/u_logic/Vsevx4 ), .ip2(n7073), .op(n7074) );
  nand2_1 U8627 ( .ip1(n7075), .ip2(n7074), .op(n7077) );
  nand2_1 U8628 ( .ip1(n12603), .ip2(\CORTEXM0DS_INST/u_logic/Qgfvx4 ), .op(
        n7076) );
  nand4_1 U8629 ( .ip1(n1120), .ip2(n1118), .ip3(n7077), .ip4(n7076), .op(
        n6019) );
  nand2_1 U8630 ( .ip1(\CORTEXM0DS_INST/u_logic/W1evx4 ), .ip2(n2119), .op(
        n8057) );
  nor2_1 U8631 ( .ip1(n2119), .ip2(n11789), .op(n12359) );
  nand2_1 U8632 ( .ip1(\CORTEXM0DS_INST/vis_pc [27]), .ip2(n12359), .op(n8056)
         );
  nor2_1 U8633 ( .ip1(n2119), .ip2(n12071), .op(n12358) );
  nand2_1 U8634 ( .ip1(\CORTEXM0DS_INST/vis_apsr [0]), .ip2(n12358), .op(n8055) );
  inv_1 U8635 ( .ip(n2119), .op(n12353) );
  nand4_1 U8636 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n9667), .ip3(
        n12118), .ip4(n11100), .op(n7078) );
  nand4_1 U8637 ( .ip1(n7079), .ip2(n11789), .ip3(n12353), .ip4(n7078), .op(
        n12355) );
  and2_1 U8638 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [28]), .op(n7087)
         );
  inv_1 U8639 ( .ip(\CORTEXM0DS_INST/u_logic/W1evx4 ), .op(n8564) );
  nor2_1 U8640 ( .ip1(n7398), .ip2(n8564), .op(n7081) );
  nor2_1 U8641 ( .ip1(n8671), .ip2(n9348), .op(n7080) );
  not_ab_or_c_or_d U8642 ( .ip1(\CORTEXM0DS_INST/u_logic/L0evx4 ), .ip2(n7438), 
        .ip3(n7081), .ip4(n7080), .op(n7085) );
  nand2_1 U8643 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [28]), .op(n7084)
         );
  nand2_1 U8644 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [28]), .op(n7083)
         );
  nand2_1 U8645 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [26]), .op(n7082)
         );
  not_ab_or_c_or_d U8646 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [28]), .ip2(n9354), 
        .ip3(n7087), .ip4(n7086), .op(n7091) );
  nand2_1 U8647 ( .ip1(n9347), .ip2(\CORTEXM0DS_INST/cm0_r14 [28]), .op(n7090)
         );
  nand2_1 U8648 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [28]), .op(n7089)
         );
  nand2_1 U8649 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [26]), .op(n7088)
         );
  inv_1 U8650 ( .ip(\CORTEXM0DS_INST/vis_pc [27]), .op(n10231) );
  nand2_1 U8651 ( .ip1(\CORTEXM0DS_INST/vis_pc [20]), .ip2(
        \CORTEXM0DS_INST/vis_pc [21]), .op(n8531) );
  nand3_1 U8652 ( .ip1(\CORTEXM0DS_INST/vis_pc [3]), .ip2(
        \CORTEXM0DS_INST/vis_pc [4]), .ip3(n8871), .op(n12281) );
  inv_1 U8653 ( .ip(\CORTEXM0DS_INST/vis_pc [5]), .op(n12280) );
  nor2_1 U8654 ( .ip1(n12281), .ip2(n12280), .op(n12332) );
  nand2_1 U8655 ( .ip1(n12332), .ip2(\CORTEXM0DS_INST/vis_pc [6]), .op(n12333)
         );
  inv_1 U8656 ( .ip(\CORTEXM0DS_INST/vis_pc [7]), .op(n12154) );
  nor2_1 U8657 ( .ip1(n12333), .ip2(n12154), .op(n12162) );
  nand2_1 U8658 ( .ip1(\CORTEXM0DS_INST/vis_pc [10]), .ip2(
        \CORTEXM0DS_INST/vis_pc [11]), .op(n10193) );
  inv_1 U8659 ( .ip(\CORTEXM0DS_INST/vis_pc [12]), .op(n10197) );
  inv_1 U8660 ( .ip(\CORTEXM0DS_INST/vis_pc [13]), .op(n10329) );
  nand2_1 U8661 ( .ip1(\CORTEXM0DS_INST/vis_pc [8]), .ip2(
        \CORTEXM0DS_INST/vis_pc [9]), .op(n8064) );
  nand2_1 U8662 ( .ip1(n12162), .ip2(n8533), .op(n11006) );
  inv_1 U8663 ( .ip(\CORTEXM0DS_INST/vis_pc [14]), .op(n11005) );
  nor2_1 U8664 ( .ip1(n11006), .ip2(n11005), .op(n12209) );
  nand2_1 U8665 ( .ip1(n12209), .ip2(\CORTEXM0DS_INST/vis_pc [15]), .op(n12221) );
  inv_1 U8666 ( .ip(\CORTEXM0DS_INST/vis_pc [16]), .op(n12220) );
  nor2_1 U8667 ( .ip1(n12221), .ip2(n12220), .op(n12240) );
  nand4_1 U8668 ( .ip1(\CORTEXM0DS_INST/vis_pc [17]), .ip2(
        \CORTEXM0DS_INST/vis_pc [18]), .ip3(\CORTEXM0DS_INST/vis_pc [19]), 
        .ip4(n12240), .op(n12261) );
  nor2_1 U8669 ( .ip1(n8531), .ip2(n12261), .op(n12270) );
  nand2_1 U8670 ( .ip1(n12270), .ip2(\CORTEXM0DS_INST/vis_pc [22]), .op(n12346) );
  inv_1 U8671 ( .ip(\CORTEXM0DS_INST/vis_pc [23]), .op(n12345) );
  nor2_1 U8672 ( .ip1(n12346), .ip2(n12345), .op(n12344) );
  nand3_1 U8673 ( .ip1(n12344), .ip2(\CORTEXM0DS_INST/vis_pc [24]), .ip3(
        \CORTEXM0DS_INST/vis_pc [25]), .op(n12310) );
  inv_1 U8674 ( .ip(\CORTEXM0DS_INST/vis_pc [26]), .op(n12309) );
  nor2_1 U8675 ( .ip1(n12310), .ip2(n12309), .op(n12308) );
  inv_1 U8676 ( .ip(n12308), .op(n9988) );
  nor2_1 U8677 ( .ip1(n10231), .ip2(n9988), .op(n10034) );
  not_ab_or_c_or_d U8678 ( .ip1(n10231), .ip2(n9988), .ip3(n10034), .ip4(
        n12343), .op(n8053) );
  and2_1 U8679 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [27]), .op(n7103)
         );
  and2_1 U8680 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [27]), .op(n7097)
         );
  nand2_1 U8681 ( .ip1(n7437), .ip2(n8768), .op(n7095) );
  nand2_1 U8682 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/L0evx4 ), .op(
        n7094) );
  nand2_1 U8683 ( .ip1(\CORTEXM0DS_INST/u_logic/Azdvx4 ), .ip2(n7438), .op(
        n7093) );
  nand2_1 U8684 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [25]), .op(n7092)
         );
  not_ab_or_c_or_d U8685 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [27]), .ip2(n9347), 
        .ip3(n7097), .ip4(n7096), .op(n7101) );
  nand2_1 U8686 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [27]), .op(n7100)
         );
  nand2_1 U8687 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [27]), .op(n7099)
         );
  nand2_1 U8688 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [25]), .op(n7098)
         );
  not_ab_or_c_or_d U8689 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [27]), 
        .ip3(n7103), .ip4(n7102), .op(n9543) );
  nand4_1 U8690 ( .ip1(\CORTEXM0DS_INST/u_logic/O8gvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip4(n9946), .op(n7632) );
  nor2_1 U8691 ( .ip1(n12384), .ip2(n7632), .op(n7937) );
  or2_1 U8692 ( .ip1(n7889), .ip2(n7937), .op(n7104) );
  nand2_1 U8693 ( .ip1(\CORTEXM0DS_INST/u_logic/Bx9vx4 ), .ip2(n7104), .op(
        n7105) );
  mux2_1 U8694 ( .ip1(n7941), .ip2(n7940), .s(n7105), .op(n9345) );
  mux2_1 U8695 ( .ip1(n7106), .ip2(n9345), .s(n7887), .op(n9346) );
  inv_1 U8696 ( .ip(n9346), .op(n8562) );
  inv_1 U8697 ( .ip(n9345), .op(n8563) );
  nand2_1 U8698 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [27]), .op(n7109)
         );
  nand2_1 U8699 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [27]), .op(n7108)
         );
  nand2_1 U8700 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [27]), .op(n7107)
         );
  nand3_1 U8701 ( .ip1(n7109), .ip2(n7108), .ip3(n7107), .op(n7126) );
  nand2_1 U8702 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [27]), .ip2(n9344), .op(n7124)
         );
  nand2_1 U8703 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [27]), .op(n7113)
         );
  nand2_1 U8704 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [27]), .op(n7112)
         );
  nand2_1 U8705 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [27]), .op(n7111)
         );
  nand2_1 U8706 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [27]), .op(n7110)
         );
  nand2_1 U8707 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [25]), .op(n7117)
         );
  nand2_1 U8708 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [25]), .op(n7116)
         );
  nand2_1 U8709 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [27]), .op(n7115)
         );
  nand2_1 U8710 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [27]), .op(n7114)
         );
  not_ab_or_c_or_d U8711 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [27]), 
        .ip3(n7119), .ip4(n7118), .op(n7123) );
  inv_1 U8712 ( .ip(n9325), .op(n9279) );
  inv_1 U8713 ( .ip(\CORTEXM0DS_INST/u_logic/L0evx4 ), .op(n12317) );
  nor2_1 U8714 ( .ip1(n9279), .ip2(n12317), .op(n7121) );
  and2_1 U8715 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [27]), .op(n7120)
         );
  not_ab_or_c_or_d U8716 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [27]), .ip2(n9317), 
        .ip3(n7121), .ip4(n7120), .op(n7122) );
  nand3_1 U8717 ( .ip1(n7124), .ip2(n7123), .ip3(n7122), .op(n7125) );
  not_ab_or_c_or_d U8718 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [27]), 
        .ip3(n7126), .ip4(n7125), .op(n10066) );
  mux2_1 U8719 ( .ip1(n8562), .ip2(n8563), .s(n10066), .op(n9546) );
  nor2_1 U8720 ( .ip1(n9543), .ip2(n9546), .op(n7127) );
  nand2_1 U8721 ( .ip1(n7127), .ip2(n9261), .op(n7969) );
  nor2_1 U8722 ( .ip1(n9371), .ip2(n9543), .op(n7128) );
  xnor2_1 U8723 ( .ip1(n9546), .ip2(n7128), .op(n7993) );
  nand2_1 U8724 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [26]), .op(n7131)
         );
  nand2_1 U8725 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [26]), .op(n7130)
         );
  nand2_1 U8726 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [26]), .op(n7129)
         );
  nand3_1 U8727 ( .ip1(n7131), .ip2(n7130), .ip3(n7129), .op(n7148) );
  and2_1 U8728 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [26]), .op(n7133)
         );
  inv_1 U8729 ( .ip(\CORTEXM0DS_INST/u_logic/Azdvx4 ), .op(n12305) );
  nor2_1 U8730 ( .ip1(n9279), .ip2(n12305), .op(n7132) );
  not_ab_or_c_or_d U8731 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [26]), 
        .ip3(n7133), .ip4(n7132), .op(n7146) );
  nand2_1 U8732 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [26]), .op(n7137)
         );
  nand2_1 U8733 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [26]), .op(n7136)
         );
  nand2_1 U8734 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [26]), .op(n7135)
         );
  nand2_1 U8735 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [26]), .op(n7134)
         );
  nand2_1 U8736 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [26]), .op(n7140)
         );
  nand2_1 U8737 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [26]), .op(n7139)
         );
  nand2_1 U8738 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [26]), .op(n7138)
         );
  nand3_1 U8739 ( .ip1(n7140), .ip2(n7139), .ip3(n7138), .op(n7141) );
  not_ab_or_c_or_d U8740 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [26]), 
        .ip3(n7142), .ip4(n7141), .op(n7145) );
  nand2_1 U8741 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [24]), .op(n7144)
         );
  nand2_1 U8742 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [24]), .op(n7143)
         );
  not_ab_or_c_or_d U8743 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [26]), 
        .ip3(n7148), .ip4(n7147), .op(n11477) );
  mux2_1 U8744 ( .ip1(n8562), .ip2(n8563), .s(n11477), .op(n11476) );
  inv_1 U8745 ( .ip(n11476), .op(n11471) );
  and2_1 U8746 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [26]), .op(n7160)
         );
  and2_1 U8747 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [26]), .op(n7154)
         );
  nand2_1 U8748 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [24]), .op(n7152)
         );
  nand2_1 U8749 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/Azdvx4 ), .op(
        n7151) );
  nand2_1 U8750 ( .ip1(n7437), .ip2(n9184), .op(n7150) );
  nand2_1 U8751 ( .ip1(\CORTEXM0DS_INST/u_logic/Pxdvx4 ), .ip2(n7438), .op(
        n7149) );
  not_ab_or_c_or_d U8752 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [26]), .ip2(n9347), 
        .ip3(n7154), .ip4(n7153), .op(n7158) );
  nand2_1 U8753 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [26]), .op(n7157)
         );
  nand2_1 U8754 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [26]), .op(n7156)
         );
  nand2_1 U8755 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [24]), .op(n7155)
         );
  not_ab_or_c_or_d U8756 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [26]), .ip2(n9354), 
        .ip3(n7160), .ip4(n7159), .op(n7964) );
  inv_1 U8757 ( .ip(n7964), .op(n12304) );
  nand2_1 U8758 ( .ip1(n11471), .ip2(n12304), .op(n11470) );
  or2_1 U8759 ( .ip1(n11470), .ip2(n9371), .op(n7967) );
  and2_1 U8760 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [25]), .op(n7172)
         );
  and2_1 U8761 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [25]), .op(n7166)
         );
  inv_1 U8762 ( .ip(n8426), .op(n9182) );
  nand2_1 U8763 ( .ip1(n7437), .ip2(n9182), .op(n7164) );
  nand2_1 U8764 ( .ip1(\CORTEXM0DS_INST/u_logic/Ewdvx4 ), .ip2(n7438), .op(
        n7163) );
  nand2_1 U8765 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/Pxdvx4 ), .op(
        n7162) );
  nand2_1 U8766 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [23]), .op(n7161)
         );
  not_ab_or_c_or_d U8767 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [25]), 
        .ip3(n7166), .ip4(n7165), .op(n7170) );
  nand2_1 U8768 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [25]), .op(n7169)
         );
  nand2_1 U8769 ( .ip1(n9347), .ip2(\CORTEXM0DS_INST/cm0_r14 [25]), .op(n7168)
         );
  nand2_1 U8770 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [23]), .op(n7167)
         );
  not_ab_or_c_or_d U8771 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [25]), .ip2(n9354), 
        .ip3(n7172), .ip4(n7171), .op(n12288) );
  nor2_1 U8772 ( .ip1(n9371), .ip2(n12288), .op(n7996) );
  nand2_1 U8773 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [25]), .op(n7175)
         );
  nand2_1 U8774 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [25]), .op(n7174)
         );
  nand2_1 U8775 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [25]), .op(n7173)
         );
  nand3_1 U8776 ( .ip1(n7175), .ip2(n7174), .ip3(n7173), .op(n7192) );
  nand2_1 U8777 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [25]), .ip2(n9316), .op(n7190)
         );
  nand2_1 U8778 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [25]), .op(n7179)
         );
  nand2_1 U8779 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [25]), .op(n7178)
         );
  nand2_1 U8780 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [25]), .op(n7177)
         );
  nand2_1 U8781 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [25]), .op(n7176)
         );
  nand2_1 U8782 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [23]), .op(n7183)
         );
  nand2_1 U8783 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [23]), .op(n7182)
         );
  nand2_1 U8784 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [25]), .op(n7181)
         );
  nand2_1 U8785 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [25]), .op(n7180)
         );
  not_ab_or_c_or_d U8786 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [25]), 
        .ip3(n7185), .ip4(n7184), .op(n7189) );
  inv_1 U8787 ( .ip(\CORTEXM0DS_INST/u_logic/Pxdvx4 ), .op(n12295) );
  nor2_1 U8788 ( .ip1(n9279), .ip2(n12295), .op(n7187) );
  and2_1 U8789 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [25]), .op(n7186)
         );
  not_ab_or_c_or_d U8790 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [25]), .ip2(n9314), 
        .ip3(n7187), .ip4(n7186), .op(n7188) );
  nand3_1 U8791 ( .ip1(n7190), .ip2(n7189), .ip3(n7188), .op(n7191) );
  not_ab_or_c_or_d U8792 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [25]), 
        .ip3(n7192), .ip4(n7191), .op(n11462) );
  mux2_1 U8793 ( .ip1(n9346), .ip2(n9345), .s(n11462), .op(n9542) );
  inv_1 U8794 ( .ip(\CORTEXM0DS_INST/cm0_r08 [24]), .op(n7955) );
  nor2_1 U8795 ( .ip1(n7325), .ip2(n7955), .op(n7200) );
  inv_1 U8796 ( .ip(\CORTEXM0DS_INST/u_logic/Ewdvx4 ), .op(n12354) );
  nor2_1 U8797 ( .ip1(n7398), .ip2(n12354), .op(n7194) );
  inv_1 U8798 ( .ip(\CORTEXM0DS_INST/u_logic/Tudvx4 ), .op(n12149) );
  nor2_1 U8799 ( .ip1(n12088), .ip2(n12149), .op(n7193) );
  not_ab_or_c_or_d U8800 ( .ip1(\CORTEXM0DS_INST/vis_msp [22]), .ip2(n9366), 
        .ip3(n7194), .ip4(n7193), .op(n7198) );
  nand2_1 U8801 ( .ip1(n9347), .ip2(\CORTEXM0DS_INST/cm0_r14 [24]), .op(n7197)
         );
  nand2_1 U8802 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [24]), .op(n7196)
         );
  nand2_1 U8803 ( .ip1(n7437), .ip2(n9178), .op(n7195) );
  not_ab_or_c_or_d U8804 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [24]), .ip2(n9364), 
        .ip3(n7200), .ip4(n7199), .op(n7204) );
  nand2_1 U8805 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [24]), .op(n7203)
         );
  nand2_1 U8806 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [24]), .op(n7202)
         );
  nand2_1 U8807 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [22]), .op(n7201)
         );
  inv_1 U8808 ( .ip(n9624), .op(n12348) );
  nor2_1 U8809 ( .ip1(n9371), .ip2(n12348), .op(n7998) );
  and2_1 U8810 ( .ip1(n9347), .ip2(\CORTEXM0DS_INST/cm0_r14 [23]), .op(n7216)
         );
  and2_1 U8811 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [23]), .op(n7210)
         );
  nand2_1 U8812 ( .ip1(\CORTEXM0DS_INST/u_logic/Itdvx4 ), .ip2(n7438), .op(
        n7208) );
  nand2_1 U8813 ( .ip1(n7437), .ip2(n9180), .op(n7207) );
  nand2_1 U8814 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/Tudvx4 ), .op(
        n7206) );
  nand2_1 U8815 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [21]), .op(n7205)
         );
  not_ab_or_c_or_d U8816 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [23]), .ip2(n9363), 
        .ip3(n7210), .ip4(n7209), .op(n7214) );
  nand2_1 U8817 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [23]), .op(n7213)
         );
  nand2_1 U8818 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [23]), .op(n7212)
         );
  nand2_1 U8819 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [21]), .op(n7211)
         );
  not_ab_or_c_or_d U8820 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [23]), .ip2(n9354), 
        .ip3(n7216), .ip4(n7215), .op(n12142) );
  nor2_1 U8821 ( .ip1(n9371), .ip2(n12142), .op(n8000) );
  and2_1 U8822 ( .ip1(n9347), .ip2(\CORTEXM0DS_INST/cm0_r14 [22]), .op(n7224)
         );
  nor2_1 U8823 ( .ip1(n8129), .ip2(n9348), .op(n7218) );
  inv_1 U8824 ( .ip(\CORTEXM0DS_INST/u_logic/Xrdvx4 ), .op(n12267) );
  nor2_1 U8825 ( .ip1(n12088), .ip2(n12267), .op(n7217) );
  not_ab_or_c_or_d U8826 ( .ip1(\CORTEXM0DS_INST/u_logic/Itdvx4 ), .ip2(n9353), 
        .ip3(n7218), .ip4(n7217), .op(n7222) );
  nand2_1 U8827 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [22]), .op(n7221)
         );
  nand2_1 U8828 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [22]), .op(n7220)
         );
  nand2_1 U8829 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [20]), .op(n7219)
         );
  not_ab_or_c_or_d U8830 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [22]), .ip2(n9363), 
        .ip3(n7224), .ip4(n7223), .op(n7228) );
  nand2_1 U8831 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [22]), .op(n7227)
         );
  nand2_1 U8832 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [22]), .op(n7226)
         );
  nand2_1 U8833 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [20]), .op(n7225)
         );
  inv_1 U8834 ( .ip(n9598), .op(n12273) );
  nor2_1 U8835 ( .ip1(n9371), .ip2(n12273), .op(n8002) );
  and2_1 U8836 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [21]), .op(n7240)
         );
  and2_1 U8837 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [21]), .op(n7234)
         );
  nand2_1 U8838 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [19]), .op(n7232)
         );
  inv_1 U8839 ( .ip(n8726), .op(n8814) );
  nand2_1 U8840 ( .ip1(n7437), .ip2(n8814), .op(n7231) );
  nand2_1 U8841 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/Xrdvx4 ), .op(
        n7230) );
  nand2_1 U8842 ( .ip1(\CORTEXM0DS_INST/u_logic/Mqdvx4 ), .ip2(n7438), .op(
        n7229) );
  not_ab_or_c_or_d U8843 ( .ip1(n9347), .ip2(\CORTEXM0DS_INST/cm0_r14 [21]), 
        .ip3(n7234), .ip4(n7233), .op(n7238) );
  nand2_1 U8844 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [21]), .op(n7237)
         );
  nand2_1 U8845 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [21]), .op(n7236)
         );
  nand2_1 U8846 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [19]), .op(n7235)
         );
  not_ab_or_c_or_d U8847 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [21]), 
        .ip3(n7240), .ip4(n7239), .op(n11410) );
  nor2_1 U8848 ( .ip1(n9371), .ip2(n11410), .op(n8004) );
  inv_1 U8849 ( .ip(\CORTEXM0DS_INST/cm0_r14 [20]), .op(n7856) );
  nor2_1 U8850 ( .ip1(n7423), .ip2(n7856), .op(n7252) );
  and2_1 U8851 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [20]), .op(n7246)
         );
  nand2_1 U8852 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [18]), .op(n7244)
         );
  nand2_1 U8853 ( .ip1(n7437), .ip2(n8815), .op(n7243) );
  nand2_1 U8854 ( .ip1(\CORTEXM0DS_INST/u_logic/Bpdvx4 ), .ip2(n7438), .op(
        n7242) );
  nand2_1 U8855 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/Mqdvx4 ), .op(
        n7241) );
  not_ab_or_c_or_d U8856 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [20]), 
        .ip3(n7246), .ip4(n7245), .op(n7250) );
  nand2_1 U8857 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [20]), .op(n7249)
         );
  nand2_1 U8858 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [20]), .op(n7248)
         );
  nand2_1 U8859 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [18]), .op(n7247)
         );
  not_ab_or_c_or_d U8860 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [20]), .ip2(n9364), 
        .ip3(n7252), .ip4(n7251), .op(n9590) );
  nor2_1 U8861 ( .ip1(n9371), .ip2(n9590), .op(n8006) );
  and2_1 U8862 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [19]), .op(n7264)
         );
  inv_1 U8863 ( .ip(\CORTEXM0DS_INST/cm0_r14 [19]), .op(n7833) );
  nor2_1 U8864 ( .ip1(n7423), .ip2(n7833), .op(n7258) );
  nand2_1 U8865 ( .ip1(\CORTEXM0DS_INST/u_logic/Qndvx4 ), .ip2(n7438), .op(
        n7256) );
  nand2_1 U8866 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/Bpdvx4 ), .op(
        n7255) );
  nand2_1 U8867 ( .ip1(n7437), .ip2(n8824), .op(n7254) );
  nand2_1 U8868 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [17]), .op(n7253)
         );
  not_ab_or_c_or_d U8869 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [19]), .ip2(n9363), 
        .ip3(n7258), .ip4(n7257), .op(n7262) );
  nand2_1 U8870 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [19]), .op(n7261)
         );
  nand2_1 U8871 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [19]), .op(n7260)
         );
  nand2_1 U8872 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [17]), .op(n7259)
         );
  not_ab_or_c_or_d U8873 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [19]), .ip2(n9365), 
        .ip3(n7264), .ip4(n7263), .op(n12239) );
  nor2_1 U8874 ( .ip1(n9371), .ip2(n12239), .op(n8008) );
  inv_1 U8875 ( .ip(n9371), .op(n9261) );
  and2_1 U8876 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [18]), .op(n7272)
         );
  inv_1 U8877 ( .ip(\CORTEXM0DS_INST/u_logic/Fmdvx4 ), .op(n12226) );
  nor2_1 U8878 ( .ip1(n12088), .ip2(n12226), .op(n7266) );
  nor2_1 U8879 ( .ip1(n8821), .ip2(n9348), .op(n7265) );
  not_ab_or_c_or_d U8880 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [16]), 
        .ip3(n7266), .ip4(n7265), .op(n7270) );
  nand2_1 U8881 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [18]), .op(n7269)
         );
  nand2_1 U8882 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [18]), .op(n7268)
         );
  nand2_1 U8883 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/Qndvx4 ), .op(
        n7267) );
  not_ab_or_c_or_d U8884 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [18]), .ip2(n9347), 
        .ip3(n7272), .ip4(n7271), .op(n7276) );
  nand2_1 U8885 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [18]), .op(n7275)
         );
  nand2_1 U8886 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [18]), .op(n7274)
         );
  nand2_1 U8887 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [16]), .op(n7273)
         );
  and2_1 U8888 ( .ip1(n9261), .ip2(n12235), .op(n8010) );
  and2_1 U8889 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [17]), .op(n7288)
         );
  and2_1 U8890 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [17]), .op(n7282)
         );
  nand2_1 U8891 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [15]), .op(n7280)
         );
  inv_1 U8892 ( .ip(n8408), .op(n8823) );
  nand2_1 U8893 ( .ip1(n7437), .ip2(n8823), .op(n7279) );
  nand2_1 U8894 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/Fmdvx4 ), .op(
        n7278) );
  nand2_1 U8895 ( .ip1(\CORTEXM0DS_INST/u_logic/Ukdvx4 ), .ip2(n7438), .op(
        n7277) );
  not_ab_or_c_or_d U8896 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [17]), .ip2(n9355), 
        .ip3(n7282), .ip4(n7281), .op(n7286) );
  nand2_1 U8897 ( .ip1(n9347), .ip2(\CORTEXM0DS_INST/cm0_r14 [17]), .op(n7285)
         );
  nand2_1 U8898 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [17]), .op(n7284)
         );
  nand2_1 U8899 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [15]), .op(n7283)
         );
  not_ab_or_c_or_d U8900 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [17]), 
        .ip3(n7288), .ip4(n7287), .op(n9557) );
  nor2_1 U8901 ( .ip1(n9371), .ip2(n9557), .op(n8012) );
  and2_1 U8902 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [16]), .op(n7300)
         );
  and2_1 U8903 ( .ip1(n9347), .ip2(\CORTEXM0DS_INST/cm0_r14 [16]), .op(n7294)
         );
  nand2_1 U8904 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [14]), .op(n7292)
         );
  nand2_1 U8905 ( .ip1(n7437), .ip2(n8822), .op(n7291) );
  nand2_1 U8906 ( .ip1(\CORTEXM0DS_INST/u_logic/Jjdvx4 ), .ip2(n7438), .op(
        n7290) );
  nand2_1 U8907 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/Ukdvx4 ), .op(
        n7289) );
  not_ab_or_c_or_d U8908 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [16]), 
        .ip3(n7294), .ip4(n7293), .op(n7298) );
  nand2_1 U8909 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [16]), .op(n7297)
         );
  nand2_1 U8910 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [16]), .op(n7296)
         );
  nand2_1 U8911 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [14]), .op(n7295)
         );
  not_ab_or_c_or_d U8912 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [16]), .ip2(n9364), 
        .ip3(n7300), .ip4(n7299), .op(n9595) );
  nor2_1 U8913 ( .ip1(n9371), .ip2(n9595), .op(n8014) );
  and2_1 U8914 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [15]), .op(n7312)
         );
  and2_1 U8915 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [15]), .op(n7306)
         );
  nand2_1 U8916 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [13]), .op(n7304)
         );
  nand2_1 U8917 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/Jjdvx4 ), .op(
        n7303) );
  nand2_1 U8918 ( .ip1(n7437), .ip2(n8718), .op(n7302) );
  nand2_1 U8919 ( .ip1(\CORTEXM0DS_INST/u_logic/Yhdvx4 ), .ip2(n7438), .op(
        n7301) );
  not_ab_or_c_or_d U8920 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [15]), 
        .ip3(n7306), .ip4(n7305), .op(n7310) );
  nand2_1 U8921 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [15]), .op(n7309)
         );
  nand2_1 U8922 ( .ip1(n9347), .ip2(\CORTEXM0DS_INST/cm0_r14 [15]), .op(n7308)
         );
  nand2_1 U8923 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [13]), .op(n7307)
         );
  not_ab_or_c_or_d U8924 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [15]), 
        .ip3(n7312), .ip4(n7311), .op(n11004) );
  nor2_1 U8925 ( .ip1(n9371), .ip2(n11004), .op(n8016) );
  and2_1 U8926 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [14]), .op(n7320)
         );
  nor2_1 U8927 ( .ip1(n9147), .ip2(n9348), .op(n7314) );
  inv_1 U8928 ( .ip(\CORTEXM0DS_INST/u_logic/Ngdvx4 ), .op(n7696) );
  nor2_1 U8929 ( .ip1(n12088), .ip2(n7696), .op(n7313) );
  not_ab_or_c_or_d U8930 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/Yhdvx4 ), 
        .ip3(n7314), .ip4(n7313), .op(n7318) );
  nand2_1 U8931 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [14]), .op(n7317)
         );
  nand2_1 U8932 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [14]), .op(n7316)
         );
  nand2_1 U8933 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [12]), .op(n7315)
         );
  not_ab_or_c_or_d U8934 ( .ip1(n9347), .ip2(\CORTEXM0DS_INST/cm0_r14 [14]), 
        .ip3(n7320), .ip4(n7319), .op(n7324) );
  nand2_1 U8935 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [14]), .op(n7323)
         );
  nand2_1 U8936 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [14]), .op(n7322)
         );
  nand2_1 U8937 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [12]), .op(n7321)
         );
  inv_1 U8938 ( .ip(n10027), .op(n9621) );
  nor2_1 U8939 ( .ip1(n9371), .ip2(n9621), .op(n8018) );
  inv_1 U8940 ( .ip(\CORTEXM0DS_INST/cm0_r08 [13]), .op(n7695) );
  nor2_1 U8941 ( .ip1(n7325), .ip2(n7695), .op(n7337) );
  and2_1 U8942 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [13]), .op(n7331)
         );
  nand2_1 U8943 ( .ip1(\CORTEXM0DS_INST/u_logic/Cfdvx4 ), .ip2(n7438), .op(
        n7329) );
  nand2_1 U8944 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/Ngdvx4 ), .op(
        n7328) );
  inv_1 U8945 ( .ip(n9149), .op(n8693) );
  nand2_1 U8946 ( .ip1(n7437), .ip2(n8693), .op(n7327) );
  nand2_1 U8947 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [11]), .op(n7326)
         );
  not_ab_or_c_or_d U8948 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [13]), .ip2(n9347), 
        .ip3(n7331), .ip4(n7330), .op(n7335) );
  nand2_1 U8949 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [13]), .op(n7334)
         );
  nand2_1 U8950 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [13]), .op(n7333)
         );
  nand2_1 U8951 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [11]), .op(n7332)
         );
  not_ab_or_c_or_d U8952 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [13]), 
        .ip3(n7337), .ip4(n7336), .op(n9617) );
  nor2_1 U8953 ( .ip1(n9371), .ip2(n9617), .op(n8020) );
  and2_1 U8954 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [12]), .op(n7349)
         );
  and2_1 U8955 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [12]), .op(n7343)
         );
  nand2_1 U8956 ( .ip1(n7437), .ip2(n8690), .op(n7341) );
  nand2_1 U8957 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [10]), .op(n7340)
         );
  nand2_1 U8958 ( .ip1(\CORTEXM0DS_INST/u_logic/Rddvx4 ), .ip2(n7438), .op(
        n7339) );
  nand2_1 U8959 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/Cfdvx4 ), .op(
        n7338) );
  not_ab_or_c_or_d U8960 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [12]), 
        .ip3(n7343), .ip4(n7342), .op(n7347) );
  nand2_1 U8961 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [12]), .op(n7346)
         );
  nand2_1 U8962 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [12]), .op(n7345)
         );
  nand2_1 U8963 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [10]), .op(n7344)
         );
  not_ab_or_c_or_d U8964 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [12]), .ip2(n9347), 
        .ip3(n7349), .ip4(n7348), .op(n11318) );
  nor2_1 U8965 ( .ip1(n9371), .ip2(n11318), .op(n8045) );
  and2_1 U8966 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [11]), .op(n7357)
         );
  inv_1 U8967 ( .ip(n8692), .op(n9161) );
  nor2_1 U8968 ( .ip1(n9161), .ip2(n9348), .op(n7351) );
  inv_1 U8969 ( .ip(\CORTEXM0DS_INST/u_logic/Gcdvx4 ), .op(n7624) );
  nor2_1 U8970 ( .ip1(n12088), .ip2(n7624), .op(n7350) );
  not_ab_or_c_or_d U8971 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [9]), 
        .ip3(n7351), .ip4(n7350), .op(n7355) );
  nand2_1 U8972 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [11]), .op(n7354)
         );
  nand2_1 U8973 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [11]), .op(n7353)
         );
  nand2_1 U8974 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/Rddvx4 ), .op(
        n7352) );
  not_ab_or_c_or_d U8975 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [11]), .ip2(n9347), 
        .ip3(n7357), .ip4(n7356), .op(n7361) );
  nand2_1 U8976 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [11]), .op(n7360)
         );
  nand2_1 U8977 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [11]), .op(n7359)
         );
  nand2_1 U8978 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [9]), .op(n7358)
         );
  inv_1 U8979 ( .ip(n12191), .op(n9619) );
  nor2_1 U8980 ( .ip1(n9371), .ip2(n9619), .op(n8042) );
  and2_1 U8981 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [10]), .op(n7369)
         );
  inv_1 U8982 ( .ip(\CORTEXM0DS_INST/u_logic/Wadvx4 ), .op(n12170) );
  nor2_1 U8983 ( .ip1(n12088), .ip2(n12170), .op(n7363) );
  nor2_1 U8984 ( .ip1(n9157), .ip2(n9348), .op(n7362) );
  not_ab_or_c_or_d U8985 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [8]), 
        .ip3(n7363), .ip4(n7362), .op(n7367) );
  nand2_1 U8986 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [10]), .op(n7366)
         );
  nand2_1 U8987 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [10]), .op(n7365)
         );
  nand2_1 U8988 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/Gcdvx4 ), .op(
        n7364) );
  not_ab_or_c_or_d U8989 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [10]), .ip2(n9347), 
        .ip3(n7369), .ip4(n7368), .op(n7373) );
  nand2_1 U8990 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [10]), .op(n7372)
         );
  nand2_1 U8991 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [10]), .op(n7371)
         );
  nand2_1 U8992 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [8]), .op(n7370)
         );
  inv_1 U8993 ( .ip(n9498), .op(n12177) );
  nor2_1 U8994 ( .ip1(n9371), .ip2(n12177), .op(n8022) );
  inv_1 U8995 ( .ip(\CORTEXM0DS_INST/cm0_r10 [9]), .op(n7584) );
  nor2_1 U8996 ( .ip1(n7436), .ip2(n7584), .op(n7385) );
  and2_1 U8997 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [9]), .op(n7379)
         );
  nand2_1 U8998 ( .ip1(\CORTEXM0DS_INST/u_logic/M9dvx4 ), .ip2(n7438), .op(
        n7377) );
  nand2_1 U8999 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/Wadvx4 ), .op(
        n7376) );
  inv_1 U9000 ( .ip(n9159), .op(n8699) );
  nand2_1 U9001 ( .ip1(n7437), .ip2(n8699), .op(n7375) );
  nand2_1 U9002 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [7]), .op(n7374)
         );
  not_ab_or_c_or_d U9003 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [9]), .ip2(n9363), 
        .ip3(n7379), .ip4(n7378), .op(n7383) );
  nand2_1 U9004 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [9]), .op(n7382)
         );
  nand2_1 U9005 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [9]), .op(n7381)
         );
  nand2_1 U9006 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [7]), .op(n7380)
         );
  not_ab_or_c_or_d U9007 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [9]), .ip2(n9347), 
        .ip3(n7385), .ip4(n7384), .op(n12166) );
  nor2_1 U9008 ( .ip1(n9371), .ip2(n12166), .op(n8024) );
  and2_1 U9009 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [8]), .op(n7397)
         );
  and2_1 U9010 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [8]), .op(n7391)
         );
  nand2_1 U9011 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [6]), .op(n7389)
         );
  nand2_1 U9012 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/M9dvx4 ), .op(
        n7388) );
  nand2_1 U9013 ( .ip1(\CORTEXM0DS_INST/u_logic/C8dvx4 ), .ip2(n7438), .op(
        n7387) );
  nand2_1 U9014 ( .ip1(n7437), .ip2(n9155), .op(n7386) );
  not_ab_or_c_or_d U9015 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [8]), .ip2(n9347), 
        .ip3(n7391), .ip4(n7390), .op(n7395) );
  nand2_1 U9016 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [8]), .op(n7394)
         );
  nand2_1 U9017 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [8]), .op(n7393)
         );
  nand2_1 U9018 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [6]), .op(n7392)
         );
  not_ab_or_c_or_d U9019 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [8]), .ip2(n9364), 
        .ip3(n7397), .ip4(n7396), .op(n9560) );
  nor2_1 U9020 ( .ip1(n9371), .ip2(n9560), .op(n8026) );
  inv_1 U9021 ( .ip(\CORTEXM0DS_INST/cm0_r14 [7]), .op(n7530) );
  nor2_1 U9022 ( .ip1(n7423), .ip2(n7530), .op(n7406) );
  inv_1 U9023 ( .ip(n8698), .op(n8791) );
  nor2_1 U9024 ( .ip1(n8791), .ip2(n9348), .op(n7400) );
  inv_1 U9025 ( .ip(\CORTEXM0DS_INST/u_logic/C8dvx4 ), .op(n12340) );
  nor2_1 U9026 ( .ip1(n7398), .ip2(n12340), .op(n7399) );
  not_ab_or_c_or_d U9027 ( .ip1(\CORTEXM0DS_INST/u_logic/S6dvx4 ), .ip2(n7438), 
        .ip3(n7400), .ip4(n7399), .op(n7404) );
  nand2_1 U9028 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [7]), .op(n7403)
         );
  nand2_1 U9029 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [7]), .op(n7402)
         );
  nand2_1 U9030 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [5]), .op(n7401)
         );
  not_ab_or_c_or_d U9031 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [7]), .ip2(n9364), 
        .ip3(n7406), .ip4(n7405), .op(n7410) );
  nand2_1 U9032 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [7]), .op(n7409)
         );
  nand2_1 U9033 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [7]), .op(n7408)
         );
  nand2_1 U9034 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [5]), .op(n7407)
         );
  and4_1 U9035 ( .ip1(n7410), .ip2(n7409), .ip3(n7408), .ip4(n7407), .op(
        n12331) );
  nor2_1 U9036 ( .ip1(n9371), .ip2(n12331), .op(n8028) );
  and2_1 U9037 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [6]), .op(n7422)
         );
  and2_1 U9038 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [6]), .op(n7416)
         );
  nand2_1 U9039 ( .ip1(n7437), .ip2(n8790), .op(n7414) );
  nand2_1 U9040 ( .ip1(\CORTEXM0DS_INST/u_logic/I5dvx4 ), .ip2(n7438), .op(
        n7413) );
  nand2_1 U9041 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/S6dvx4 ), .op(
        n7412) );
  nand2_1 U9042 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [4]), .op(n7411)
         );
  not_ab_or_c_or_d U9043 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [6]), .ip2(n9347), 
        .ip3(n7416), .ip4(n7415), .op(n7420) );
  nand2_1 U9044 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [6]), .op(n7419)
         );
  nand2_1 U9045 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [6]), .op(n7418)
         );
  nand2_1 U9046 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [4]), .op(n7417)
         );
  not_ab_or_c_or_d U9047 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [6]), .ip2(n9364), 
        .ip3(n7422), .ip4(n7421), .op(n9610) );
  nor2_1 U9048 ( .ip1(n9371), .ip2(n9610), .op(n8030) );
  inv_1 U9049 ( .ip(\CORTEXM0DS_INST/cm0_r14 [5]), .op(n7479) );
  nor2_1 U9050 ( .ip1(n7423), .ip2(n7479), .op(n7435) );
  and2_1 U9051 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [5]), .op(n7429)
         );
  nand2_1 U9052 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [3]), .op(n7427)
         );
  nand2_1 U9053 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/I5dvx4 ), .op(
        n7426) );
  nand2_1 U9054 ( .ip1(n7437), .ip2(n8643), .op(n7425) );
  nand2_1 U9055 ( .ip1(\CORTEXM0DS_INST/u_logic/Y3dvx4 ), .ip2(n7438), .op(
        n7424) );
  not_ab_or_c_or_d U9056 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [5]), .ip2(n9354), 
        .ip3(n7429), .ip4(n7428), .op(n7433) );
  nand2_1 U9057 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [5]), .op(n7432)
         );
  nand2_1 U9058 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [5]), .op(n7431)
         );
  nand2_1 U9059 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [3]), .op(n7430)
         );
  not_ab_or_c_or_d U9060 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [5]), 
        .ip3(n7435), .ip4(n7434), .op(n9458) );
  nor2_1 U9061 ( .ip1(n9371), .ip2(n9458), .op(n8032) );
  and2_1 U9062 ( .ip1(n9347), .ip2(\CORTEXM0DS_INST/cm0_r14 [4]), .op(n7450)
         );
  inv_1 U9063 ( .ip(\CORTEXM0DS_INST/cm0_r10 [4]), .op(n7453) );
  nor2_1 U9064 ( .ip1(n7436), .ip2(n7453), .op(n7444) );
  nand2_1 U9065 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [2]), .op(n7442)
         );
  nand2_1 U9066 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/Y3dvx4 ), .op(
        n7441) );
  nand2_1 U9067 ( .ip1(n7437), .ip2(n8462), .op(n7440) );
  nand2_1 U9068 ( .ip1(\CORTEXM0DS_INST/u_logic/O2dvx4 ), .ip2(n7438), .op(
        n7439) );
  not_ab_or_c_or_d U9069 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [4]), .ip2(n9354), 
        .ip3(n7444), .ip4(n7443), .op(n7448) );
  nand2_1 U9070 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [4]), .op(n7447)
         );
  nand2_1 U9071 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [4]), .op(n7446)
         );
  nand2_1 U9072 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [2]), .op(n7445)
         );
  not_ab_or_c_or_d U9073 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [4]), .ip2(n9364), 
        .ip3(n7450), .ip4(n7449), .op(n9571) );
  nor2_1 U9074 ( .ip1(n9371), .ip2(n9571), .op(n8034) );
  fulladder U9075 ( .a(n7452), .b(n7451), .ci(n9481), .co(n8033), .s(n8035) );
  nand2_1 U9076 ( .ip1(n7889), .ip2(\CORTEXM0DS_INST/u_logic/P39vx4 ), .op(
        n7476) );
  nand2_1 U9077 ( .ip1(\CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip2(n7478), .op(
        n7475) );
  nand2_1 U9078 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(n7551), .op(
        n7474) );
  and2_1 U9079 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [4]), .op(n7455)
         );
  nor2_1 U9080 ( .ip1(n7585), .ip2(n7453), .op(n7454) );
  not_ab_or_c_or_d U9081 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [2]), 
        .ip3(n7455), .ip4(n7454), .op(n7472) );
  nand2_1 U9082 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [4]), .ip2(n9344), .op(n7464)
         );
  and2_1 U9083 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [4]), .op(n7461)
         );
  nand2_1 U9084 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [4]), .op(n7459)
         );
  nand2_1 U9085 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [4]), .op(n7458)
         );
  nand2_1 U9086 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [4]), .op(n7457)
         );
  nand2_1 U9087 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [4]), .op(n7456)
         );
  not_ab_or_c_or_d U9088 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [4]), 
        .ip3(n7461), .ip4(n7460), .op(n7463) );
  nand2_1 U9089 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [4]), .op(n7462)
         );
  nand3_1 U9090 ( .ip1(n7464), .ip2(n7463), .ip3(n7462), .op(n8104) );
  nand2_1 U9091 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [4]), .ip2(n9326), .op(n7467)
         );
  nand2_1 U9092 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [4]), .op(n7466)
         );
  nand2_1 U9093 ( .ip1(n9325), .ip2(\CORTEXM0DS_INST/u_logic/Y3dvx4 ), .op(
        n7465) );
  nand3_1 U9094 ( .ip1(n7467), .ip2(n7466), .ip3(n7465), .op(n7468) );
  not_ab_or_c_or_d U9095 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [4]), .ip2(n9317), 
        .ip3(n8104), .ip4(n7468), .op(n7471) );
  nand2_1 U9096 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [2]), .op(n7470)
         );
  nand2_1 U9097 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [4]), .op(n7469)
         );
  nand2_1 U9098 ( .ip1(n7938), .ip2(n12675), .op(n7473) );
  mux2_1 U9099 ( .ip1(n7940), .ip2(n7941), .s(n7477), .op(n9566) );
  nand2_1 U9100 ( .ip1(n7889), .ip2(\CORTEXM0DS_INST/u_logic/W49vx4 ), .op(
        n7503) );
  nand2_1 U9101 ( .ip1(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .ip2(n7478), .op(
        n7502) );
  and2_1 U9102 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [5]), .op(n7481)
         );
  nor2_1 U9103 ( .ip1(n7857), .ip2(n7479), .op(n7480) );
  not_ab_or_c_or_d U9104 ( .ip1(\CORTEXM0DS_INST/vis_psp [3]), .ip2(n9323), 
        .ip3(n7481), .ip4(n7480), .op(n7499) );
  nand2_1 U9105 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [5]), .op(n7491)
         );
  nor2_1 U9106 ( .ip1(n7788), .ip2(n7482), .op(n7488) );
  nand2_1 U9107 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [5]), .op(n7486)
         );
  nand2_1 U9108 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [5]), .op(n7485)
         );
  nand2_1 U9109 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [5]), .op(n7484)
         );
  nand2_1 U9110 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [5]), .op(n7483)
         );
  not_ab_or_c_or_d U9111 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [5]), 
        .ip3(n7488), .ip4(n7487), .op(n7490) );
  nand2_1 U9112 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [5]), .op(n7489)
         );
  nand3_1 U9113 ( .ip1(n7491), .ip2(n7490), .ip3(n7489), .op(n8120) );
  nand2_1 U9114 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [5]), .op(n7494)
         );
  nand2_1 U9115 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [5]), .op(n7493)
         );
  nand2_1 U9116 ( .ip1(n9325), .ip2(\CORTEXM0DS_INST/u_logic/I5dvx4 ), .op(
        n7492) );
  nand3_1 U9117 ( .ip1(n7494), .ip2(n7493), .ip3(n7492), .op(n7495) );
  not_ab_or_c_or_d U9118 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [5]), .ip2(n9317), 
        .ip3(n8120), .ip4(n7495), .op(n7498) );
  nand2_1 U9119 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [3]), .op(n7497)
         );
  nand2_1 U9120 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [5]), .op(n7496)
         );
  nand2_1 U9121 ( .ip1(n7938), .ip2(n12679), .op(n7501) );
  nand2_1 U9122 ( .ip1(\CORTEXM0DS_INST/u_logic/Cq9vx4 ), .ip2(n7551), .op(
        n7500) );
  mux2_1 U9123 ( .ip1(n7940), .ip2(n7941), .s(n7504), .op(n9463) );
  and2_1 U9124 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [6]), .op(n7506)
         );
  and2_1 U9125 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [6]), .op(n7505)
         );
  not_ab_or_c_or_d U9126 ( .ip1(\CORTEXM0DS_INST/vis_psp [4]), .ip2(n9323), 
        .ip3(n7506), .ip4(n7505), .op(n7523) );
  nand2_1 U9127 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [6]), .op(n7515)
         );
  and2_1 U9128 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [6]), .op(n7512)
         );
  nand2_1 U9129 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [6]), .op(n7510)
         );
  nand2_1 U9130 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [6]), .op(n7509)
         );
  nand2_1 U9131 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [6]), .op(n7508)
         );
  nand2_1 U9132 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [6]), .op(n7507)
         );
  not_ab_or_c_or_d U9133 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [6]), .ip2(n9344), 
        .ip3(n7512), .ip4(n7511), .op(n7514) );
  nand2_1 U9134 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [6]), .op(n7513)
         );
  nand3_1 U9135 ( .ip1(n7515), .ip2(n7514), .ip3(n7513), .op(n8115) );
  nand2_1 U9136 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [6]), .op(n7518)
         );
  nand2_1 U9137 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [6]), .op(n7517)
         );
  nand2_1 U9138 ( .ip1(n9325), .ip2(\CORTEXM0DS_INST/u_logic/S6dvx4 ), .op(
        n7516) );
  nand3_1 U9139 ( .ip1(n7518), .ip2(n7517), .ip3(n7516), .op(n7519) );
  not_ab_or_c_or_d U9140 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [6]), .ip2(n9334), 
        .ip3(n8115), .ip4(n7519), .op(n7522) );
  nand2_1 U9141 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [4]), .op(n7521)
         );
  nand2_1 U9142 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [6]), .op(n7520)
         );
  nand2_1 U9143 ( .ip1(n7938), .ip2(n12681), .op(n7528) );
  nand2_1 U9144 ( .ip1(\CORTEXM0DS_INST/u_logic/Gr9vx4 ), .ip2(n7551), .op(
        n7527) );
  nor2_1 U9145 ( .ip1(n7524), .ip2(n9797), .op(n7583) );
  nand2_1 U9146 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(n7583), .op(
        n7526) );
  nand2_1 U9147 ( .ip1(n7889), .ip2(\CORTEXM0DS_INST/u_logic/D69vx4 ), .op(
        n7525) );
  mux2_1 U9148 ( .ip1(n7940), .ip2(n7941), .s(n7529), .op(n9611) );
  nor2_1 U9149 ( .ip1(n7857), .ip2(n7530), .op(n7532) );
  and2_1 U9150 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [7]), .op(n7531)
         );
  not_ab_or_c_or_d U9151 ( .ip1(\CORTEXM0DS_INST/vis_msp [5]), .ip2(n9333), 
        .ip3(n7532), .ip4(n7531), .op(n7550) );
  nand2_1 U9152 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [7]), .op(n7542)
         );
  nor2_1 U9153 ( .ip1(n7788), .ip2(n7533), .op(n7539) );
  nand2_1 U9154 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [7]), .op(n7537)
         );
  nand2_1 U9155 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [7]), .op(n7536)
         );
  nand2_1 U9156 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [7]), .op(n7535)
         );
  nand2_1 U9157 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [7]), .op(n7534)
         );
  not_ab_or_c_or_d U9158 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [7]), .ip2(n9314), 
        .ip3(n7539), .ip4(n7538), .op(n7541) );
  nand2_1 U9159 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [7]), .op(n7540)
         );
  nand3_1 U9160 ( .ip1(n7542), .ip2(n7541), .ip3(n7540), .op(n8116) );
  nand2_1 U9161 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [7]), .op(n7545)
         );
  nand2_1 U9162 ( .ip1(n9325), .ip2(\CORTEXM0DS_INST/u_logic/C8dvx4 ), .op(
        n7544) );
  nand2_1 U9163 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [7]), .op(n7543)
         );
  nand3_1 U9164 ( .ip1(n7545), .ip2(n7544), .ip3(n7543), .op(n7546) );
  not_ab_or_c_or_d U9165 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [7]), .ip2(n9317), 
        .ip3(n8116), .ip4(n7546), .op(n7549) );
  nand2_1 U9166 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [7]), .op(n7548)
         );
  nand2_1 U9167 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [5]), .op(n7547)
         );
  nand2_1 U9168 ( .ip1(n7938), .ip2(n12685), .op(n7555) );
  nand2_1 U9169 ( .ip1(\CORTEXM0DS_INST/u_logic/Ks9vx4 ), .ip2(n7551), .op(
        n7554) );
  nand2_1 U9170 ( .ip1(\CORTEXM0DS_INST/u_logic/Cq9vx4 ), .ip2(n7583), .op(
        n7553) );
  nand2_1 U9171 ( .ip1(n7889), .ip2(\CORTEXM0DS_INST/u_logic/K79vx4 ), .op(
        n7552) );
  mux2_1 U9172 ( .ip1(n7940), .ip2(n7941), .s(n7556), .op(n9447) );
  nand2_1 U9173 ( .ip1(n7889), .ip2(\CORTEXM0DS_INST/u_logic/R89vx4 ), .op(
        n7580) );
  inv_1 U9174 ( .ip(n7632), .op(n7582) );
  nand2_1 U9175 ( .ip1(\CORTEXM0DS_INST/u_logic/Ot9vx4 ), .ip2(n7582), .op(
        n7579) );
  nand2_1 U9176 ( .ip1(\CORTEXM0DS_INST/u_logic/Gr9vx4 ), .ip2(n7583), .op(
        n7578) );
  inv_1 U9177 ( .ip(\CORTEXM0DS_INST/u_logic/M9dvx4 ), .op(n12159) );
  nor2_1 U9178 ( .ip1(n9279), .ip2(n12159), .op(n7558) );
  and2_1 U9179 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [8]), .op(n7557)
         );
  not_ab_or_c_or_d U9180 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [8]), .ip2(n9338), 
        .ip3(n7558), .ip4(n7557), .op(n7576) );
  nand2_1 U9181 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [8]), .op(n7562)
         );
  nand2_1 U9182 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [8]), .op(n7561)
         );
  nand2_1 U9183 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [8]), .op(n7560)
         );
  nand2_1 U9184 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [8]), .op(n7559)
         );
  and4_1 U9185 ( .ip1(n7562), .ip2(n7561), .ip3(n7560), .ip4(n7559), .op(n7575) );
  nand2_1 U9186 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [8]), .op(n7566)
         );
  nand2_1 U9187 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [8]), .op(n7565)
         );
  nand2_1 U9188 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [8]), .op(n7564)
         );
  nand2_1 U9189 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [8]), .op(n7563)
         );
  nand2_1 U9190 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [6]), .op(n7570)
         );
  nand2_1 U9191 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [8]), .op(n7569)
         );
  nand2_1 U9192 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [8]), .op(n7568)
         );
  nand2_1 U9193 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [8]), .op(n7567)
         );
  not_ab_or_c_or_d U9194 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [6]), 
        .ip3(n7572), .ip4(n7571), .op(n7574) );
  nand2_1 U9195 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [8]), .op(n7573)
         );
  nand2_1 U9196 ( .ip1(n7938), .ip2(n12661), .op(n7577) );
  mux2_1 U9197 ( .ip1(n7940), .ip2(n7941), .s(n7581), .op(n11559) );
  nand2_1 U9198 ( .ip1(\CORTEXM0DS_INST/u_logic/Su9vx4 ), .ip2(n7582), .op(
        n7609) );
  nand2_1 U9199 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n7889), .op(
        n7608) );
  nand2_1 U9200 ( .ip1(\CORTEXM0DS_INST/u_logic/Ks9vx4 ), .ip2(n7583), .op(
        n7607) );
  nor2_1 U9201 ( .ip1(n7585), .ip2(n7584), .op(n7587) );
  nor2_1 U9202 ( .ip1(n9279), .ip2(n12170), .op(n7586) );
  not_ab_or_c_or_d U9203 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [9]), 
        .ip3(n7587), .ip4(n7586), .op(n7605) );
  nand2_1 U9204 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [9]), .op(n7591)
         );
  nand2_1 U9205 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [9]), .op(n7590)
         );
  nand2_1 U9206 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [9]), .op(n7589)
         );
  nand2_1 U9207 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [9]), .op(n7588)
         );
  and4_1 U9208 ( .ip1(n7591), .ip2(n7590), .ip3(n7589), .ip4(n7588), .op(n7604) );
  nand2_1 U9209 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [9]), .op(n7595)
         );
  nand2_1 U9210 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [9]), .op(n7594)
         );
  nand2_1 U9211 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [9]), .op(n7593)
         );
  nand2_1 U9212 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [9]), .op(n7592)
         );
  nand2_1 U9213 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [7]), .op(n7599)
         );
  nand2_1 U9214 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [7]), .op(n7598)
         );
  nand2_1 U9215 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [9]), .op(n7597)
         );
  nand2_1 U9216 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [9]), .op(n7596)
         );
  not_ab_or_c_or_d U9217 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [9]), 
        .ip3(n7601), .ip4(n7600), .op(n7603) );
  nand2_1 U9218 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [9]), .op(n7602)
         );
  nand2_1 U9219 ( .ip1(n7938), .ip2(n12662), .op(n7606) );
  mux2_1 U9220 ( .ip1(n7940), .ip2(n7941), .s(n7610), .op(n9466) );
  nand2_1 U9221 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [10]), .op(n7613)
         );
  nand2_1 U9222 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [10]), .op(n7612)
         );
  nand2_1 U9223 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [10]), .op(n7611)
         );
  nand3_1 U9224 ( .ip1(n7613), .ip2(n7612), .ip3(n7611), .op(n7631) );
  nand2_1 U9225 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [10]), .ip2(n9315), .op(n7629)
         );
  nand2_1 U9226 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [10]), .op(n7617)
         );
  nand2_1 U9227 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [10]), .op(n7616)
         );
  nand2_1 U9228 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [10]), .op(n7615)
         );
  nand2_1 U9229 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [10]), .op(n7614)
         );
  nand2_1 U9230 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [8]), .op(n7621)
         );
  nand2_1 U9231 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [8]), .op(n7620)
         );
  nand2_1 U9232 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [10]), .op(n7619)
         );
  nand2_1 U9233 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [10]), .op(n7618)
         );
  not_ab_or_c_or_d U9234 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [10]), 
        .ip3(n7623), .ip4(n7622), .op(n7628) );
  and2_1 U9235 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [10]), .op(n7626)
         );
  nor2_1 U9236 ( .ip1(n9279), .ip2(n7624), .op(n7625) );
  not_ab_or_c_or_d U9237 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [10]), .ip2(n9335), 
        .ip3(n7626), .ip4(n7625), .op(n7627) );
  nand3_1 U9238 ( .ip1(n7629), .ip2(n7628), .ip3(n7627), .op(n7630) );
  not_ab_or_c_or_d U9239 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [10]), 
        .ip3(n7631), .ip4(n7630), .op(n10063) );
  nor2_1 U9240 ( .ip1(n10063), .ip2(n7887), .op(n7634) );
  nor2_1 U9241 ( .ip1(n12362), .ip2(n7632), .op(n7633) );
  not_ab_or_c_or_d U9242 ( .ip1(n7889), .ip2(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), 
        .ip3(n7634), .ip4(n7633), .op(n7635) );
  mux2_1 U9243 ( .ip1(n7941), .ip2(n7940), .s(n7635), .op(n9497) );
  nand2_1 U9244 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [11]), .op(n7638)
         );
  nand2_1 U9245 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [11]), .op(n7637)
         );
  nand2_1 U9246 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [11]), .op(n7636)
         );
  nand3_1 U9247 ( .ip1(n7638), .ip2(n7637), .ip3(n7636), .op(n7655) );
  nand2_1 U9248 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [11]), .ip2(n9318), .op(n7653)
         );
  nand2_1 U9249 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [11]), .op(n7642)
         );
  nand2_1 U9250 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [11]), .op(n7641)
         );
  nand2_1 U9251 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [11]), .op(n7640)
         );
  nand2_1 U9252 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [11]), .op(n7639)
         );
  nand2_1 U9253 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [9]), .op(n7646)
         );
  nand2_1 U9254 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [9]), .op(n7645)
         );
  nand2_1 U9255 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [11]), .op(n7644)
         );
  nand2_1 U9256 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [11]), .op(n7643)
         );
  not_ab_or_c_or_d U9257 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [11]), 
        .ip3(n7648), .ip4(n7647), .op(n7652) );
  and2_1 U9258 ( .ip1(n9325), .ip2(\CORTEXM0DS_INST/u_logic/Rddvx4 ), .op(
        n7650) );
  and2_1 U9259 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [11]), .op(n7649)
         );
  not_ab_or_c_or_d U9260 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [11]), .ip2(n9317), 
        .ip3(n7650), .ip4(n7649), .op(n7651) );
  nand3_1 U9261 ( .ip1(n7653), .ip2(n7652), .ip3(n7651), .op(n7654) );
  not_ab_or_c_or_d U9262 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [11]), 
        .ip3(n7655), .ip4(n7654), .op(n12665) );
  nor2_1 U9263 ( .ip1(n12665), .ip2(n7887), .op(n7656) );
  not_ab_or_c_or_d U9264 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n7889), 
        .ip3(n7937), .ip4(n7656), .op(n7657) );
  mux2_1 U9265 ( .ip1(n7941), .ip2(n7940), .s(n7657), .op(n9618) );
  nand2_1 U9266 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [12]), .op(n7660)
         );
  nand2_1 U9267 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [12]), .op(n7659)
         );
  nand2_1 U9268 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [12]), .op(n7658)
         );
  nand3_1 U9269 ( .ip1(n7660), .ip2(n7659), .ip3(n7658), .op(n7679) );
  inv_1 U9270 ( .ip(\CORTEXM0DS_INST/u_logic/Cfdvx4 ), .op(n12202) );
  nor2_1 U9271 ( .ip1(n9279), .ip2(n12202), .op(n7661) );
  or2_1 U9272 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [12]), .ip2(n7661), .op(n7663)
         );
  or2_1 U9273 ( .ip1(n9308), .ip2(n7661), .op(n7662) );
  nand2_1 U9274 ( .ip1(n7663), .ip2(n7662), .op(n7677) );
  nand2_1 U9275 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [12]), .op(n7667)
         );
  nand2_1 U9276 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [12]), .op(n7666)
         );
  nand2_1 U9277 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [12]), .op(n7665)
         );
  nand2_1 U9278 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [12]), .op(n7664)
         );
  nand2_1 U9279 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [10]), .op(n7671)
         );
  nand2_1 U9280 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [10]), .op(n7670)
         );
  nand2_1 U9281 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [12]), .op(n7669)
         );
  nand2_1 U9282 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [12]), .op(n7668)
         );
  not_ab_or_c_or_d U9283 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [12]), 
        .ip3(n7673), .ip4(n7672), .op(n7676) );
  nand2_1 U9284 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [12]), .op(n7675)
         );
  nand2_1 U9285 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [12]), .op(n7674)
         );
  not_ab_or_c_or_d U9286 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [12]), 
        .ip3(n7679), .ip4(n7678), .op(n11315) );
  nor2_1 U9287 ( .ip1(n11315), .ip2(n7887), .op(n7680) );
  not_ab_or_c_or_d U9288 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n7889), 
        .ip3(n7937), .ip4(n7680), .op(n7681) );
  mux2_1 U9289 ( .ip1(n7941), .ip2(n7940), .s(n7681), .op(n9592) );
  nand2_1 U9290 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [13]), .op(n7684)
         );
  nand2_1 U9291 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [13]), .op(n7683)
         );
  nand2_1 U9292 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [13]), .op(n7682)
         );
  nand3_1 U9293 ( .ip1(n7684), .ip2(n7683), .ip3(n7682), .op(n7703) );
  nand2_1 U9294 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [13]), .ip2(n9314), .op(n7701)
         );
  nand2_1 U9295 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [13]), .op(n7688)
         );
  nand2_1 U9296 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [13]), .op(n7687)
         );
  nand2_1 U9297 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [13]), .op(n7686)
         );
  nand2_1 U9298 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [13]), .op(n7685)
         );
  nand2_1 U9299 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [11]), .op(n7692)
         );
  nand2_1 U9300 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [11]), .op(n7691)
         );
  nand2_1 U9301 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [13]), .op(n7690)
         );
  nand2_1 U9302 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [13]), .op(n7689)
         );
  not_ab_or_c_or_d U9303 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [13]), 
        .ip3(n7694), .ip4(n7693), .op(n7700) );
  nor2_1 U9304 ( .ip1(n7956), .ip2(n7695), .op(n7698) );
  nor2_1 U9305 ( .ip1(n9279), .ip2(n7696), .op(n7697) );
  not_ab_or_c_or_d U9306 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [13]), .ip2(n9308), 
        .ip3(n7698), .ip4(n7697), .op(n7699) );
  nand3_1 U9307 ( .ip1(n7701), .ip2(n7700), .ip3(n7699), .op(n7702) );
  not_ab_or_c_or_d U9308 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [13]), 
        .ip3(n7703), .ip4(n7702), .op(n11330) );
  nor2_1 U9309 ( .ip1(n11330), .ip2(n7887), .op(n7704) );
  not_ab_or_c_or_d U9310 ( .ip1(\CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip2(n7889), 
        .ip3(n7937), .ip4(n7704), .op(n7705) );
  mux2_1 U9311 ( .ip1(n7941), .ip2(n7940), .s(n7705), .op(n9616) );
  nand2_1 U9312 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [14]), .op(n7708)
         );
  nand2_1 U9313 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [14]), .op(n7707)
         );
  nand2_1 U9314 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [14]), .op(n7706)
         );
  nand3_1 U9315 ( .ip1(n7708), .ip2(n7707), .ip3(n7706), .op(n7725) );
  nand2_1 U9316 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [14]), .ip2(n9344), .op(n7723)
         );
  nand2_1 U9317 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [14]), .op(n7712)
         );
  nand2_1 U9318 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [14]), .op(n7711)
         );
  nand2_1 U9319 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [14]), .op(n7710)
         );
  nand2_1 U9320 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [14]), .op(n7709)
         );
  nand2_1 U9321 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [12]), .op(n7716)
         );
  nand2_1 U9322 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [14]), .op(n7715)
         );
  nand2_1 U9323 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [14]), .op(n7714)
         );
  nand2_1 U9324 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [14]), .op(n7713)
         );
  not_ab_or_c_or_d U9325 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [12]), 
        .ip3(n7718), .ip4(n7717), .op(n7722) );
  and2_1 U9326 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [14]), .op(n7720)
         );
  and2_1 U9327 ( .ip1(n9325), .ip2(\CORTEXM0DS_INST/u_logic/Yhdvx4 ), .op(
        n7719) );
  not_ab_or_c_or_d U9328 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [14]), .ip2(n9316), 
        .ip3(n7720), .ip4(n7719), .op(n7721) );
  nand3_1 U9329 ( .ip1(n7723), .ip2(n7722), .ip3(n7721), .op(n7724) );
  not_ab_or_c_or_d U9330 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [14]), 
        .ip3(n7725), .ip4(n7724), .op(n11340) );
  nor2_1 U9331 ( .ip1(n11340), .ip2(n7887), .op(n7726) );
  not_ab_or_c_or_d U9332 ( .ip1(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .ip2(n7889), 
        .ip3(n7937), .ip4(n7726), .op(n7727) );
  mux2_1 U9333 ( .ip1(n7941), .ip2(n7940), .s(n7727), .op(n9620) );
  nand2_1 U9334 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [15]), .op(n7730)
         );
  nand2_1 U9335 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [15]), .op(n7729)
         );
  nand2_1 U9336 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [15]), .op(n7728)
         );
  nand3_1 U9337 ( .ip1(n7730), .ip2(n7729), .ip3(n7728), .op(n7747) );
  nand2_1 U9338 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [15]), .ip2(n9308), .op(n7745)
         );
  nand2_1 U9339 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [15]), .op(n7734)
         );
  nand2_1 U9340 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [15]), .op(n7733)
         );
  nand2_1 U9341 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [15]), .op(n7732)
         );
  nand2_1 U9342 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [15]), .op(n7731)
         );
  nand2_1 U9343 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [13]), .op(n7738)
         );
  nand2_1 U9344 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [13]), .op(n7737)
         );
  nand2_1 U9345 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [15]), .op(n7736)
         );
  nand2_1 U9346 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [15]), .op(n7735)
         );
  not_ab_or_c_or_d U9347 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [15]), 
        .ip3(n7740), .ip4(n7739), .op(n7744) );
  and2_1 U9348 ( .ip1(n9325), .ip2(\CORTEXM0DS_INST/u_logic/Jjdvx4 ), .op(
        n7742) );
  and2_1 U9349 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [15]), .op(n7741)
         );
  not_ab_or_c_or_d U9350 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [15]), .ip2(n9317), 
        .ip3(n7742), .ip4(n7741), .op(n7743) );
  nand3_1 U9351 ( .ip1(n7745), .ip2(n7744), .ip3(n7743), .op(n7746) );
  not_ab_or_c_or_d U9352 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [15]), 
        .ip3(n7747), .ip4(n7746), .op(n10071) );
  nor2_1 U9353 ( .ip1(n10071), .ip2(n7887), .op(n7748) );
  not_ab_or_c_or_d U9354 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(n7889), 
        .ip3(n7937), .ip4(n7748), .op(n7749) );
  mux2_1 U9355 ( .ip1(n7941), .ip2(n7940), .s(n7749), .op(n9593) );
  nand2_1 U9356 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [16]), .op(n7752)
         );
  nand2_1 U9357 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [16]), .op(n7751)
         );
  nand2_1 U9358 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [16]), .op(n7750)
         );
  nand3_1 U9359 ( .ip1(n7752), .ip2(n7751), .ip3(n7750), .op(n7771) );
  inv_1 U9360 ( .ip(\CORTEXM0DS_INST/u_logic/Ukdvx4 ), .op(n12217) );
  nor2_1 U9361 ( .ip1(n9279), .ip2(n12217), .op(n7753) );
  or2_1 U9362 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [16]), .ip2(n7753), .op(n7755)
         );
  or2_1 U9363 ( .ip1(n9316), .ip2(n7753), .op(n7754) );
  nand2_1 U9364 ( .ip1(n7755), .ip2(n7754), .op(n7769) );
  nand2_1 U9365 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [16]), .op(n7759)
         );
  nand2_1 U9366 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [16]), .op(n7758)
         );
  nand2_1 U9367 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [16]), .op(n7757)
         );
  nand2_1 U9368 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [16]), .op(n7756)
         );
  nand2_1 U9369 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [14]), .op(n7763)
         );
  nand2_1 U9370 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [14]), .op(n7762)
         );
  nand2_1 U9371 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [16]), .op(n7761)
         );
  nand2_1 U9372 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [16]), .op(n7760)
         );
  not_ab_or_c_or_d U9373 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [16]), 
        .ip3(n7765), .ip4(n7764), .op(n7768) );
  nand2_1 U9374 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [16]), .op(n7767)
         );
  nand2_1 U9375 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [16]), .op(n7766)
         );
  not_ab_or_c_or_d U9376 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [16]), 
        .ip3(n7771), .ip4(n7770), .op(n9612) );
  nor2_1 U9377 ( .ip1(n9612), .ip2(n7887), .op(n7772) );
  not_ab_or_c_or_d U9378 ( .ip1(\CORTEXM0DS_INST/u_logic/Cq9vx4 ), .ip2(n7889), 
        .ip3(n7937), .ip4(n7772), .op(n7773) );
  mux2_1 U9379 ( .ip1(n7941), .ip2(n7940), .s(n7773), .op(n9596) );
  nand2_1 U9380 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [17]), .op(n7776)
         );
  nand2_1 U9381 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [17]), .op(n7775)
         );
  nand2_1 U9382 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [17]), .op(n7774)
         );
  nand3_1 U9383 ( .ip1(n7776), .ip2(n7775), .ip3(n7774), .op(n7795) );
  nand2_1 U9384 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [17]), .ip2(n9344), .op(n7793)
         );
  nand2_1 U9385 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [17]), .op(n7780)
         );
  nand2_1 U9386 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [17]), .op(n7779)
         );
  nand2_1 U9387 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [17]), .op(n7778)
         );
  nand2_1 U9388 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [17]), .op(n7777)
         );
  nand2_1 U9389 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [15]), .op(n7784)
         );
  nand2_1 U9390 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [15]), .op(n7783)
         );
  nand2_1 U9391 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [17]), .op(n7782)
         );
  nand2_1 U9392 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [17]), .op(n7781)
         );
  not_ab_or_c_or_d U9393 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [17]), 
        .ip3(n7786), .ip4(n7785), .op(n7792) );
  nor2_1 U9394 ( .ip1(n7788), .ip2(n7787), .op(n7790) );
  nor2_1 U9395 ( .ip1(n9279), .ip2(n12226), .op(n7789) );
  not_ab_or_c_or_d U9396 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [17]), .ip2(n9317), 
        .ip3(n7790), .ip4(n7789), .op(n7791) );
  nand3_1 U9397 ( .ip1(n7793), .ip2(n7792), .ip3(n7791), .op(n7794) );
  not_ab_or_c_or_d U9398 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [17]), 
        .ip3(n7795), .ip4(n7794), .op(n12672) );
  nor2_1 U9399 ( .ip1(n12672), .ip2(n7887), .op(n7796) );
  not_ab_or_c_or_d U9400 ( .ip1(\CORTEXM0DS_INST/u_logic/Gr9vx4 ), .ip2(n7889), 
        .ip3(n7937), .ip4(n7796), .op(n7797) );
  mux2_1 U9401 ( .ip1(n7941), .ip2(n7940), .s(n7797), .op(n11362) );
  nand2_1 U9402 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [18]), .op(n7800)
         );
  nand2_1 U9403 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [18]), .op(n7799)
         );
  nand2_1 U9404 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [18]), .op(n7798)
         );
  nand3_1 U9405 ( .ip1(n7800), .ip2(n7799), .ip3(n7798), .op(n7817) );
  and2_1 U9406 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [18]), .op(n7802)
         );
  inv_1 U9407 ( .ip(\CORTEXM0DS_INST/u_logic/Qndvx4 ), .op(n12236) );
  nor2_1 U9408 ( .ip1(n9279), .ip2(n12236), .op(n7801) );
  not_ab_or_c_or_d U9409 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [18]), .ip2(n9308), 
        .ip3(n7802), .ip4(n7801), .op(n7815) );
  nand2_1 U9410 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [18]), .op(n7806)
         );
  nand2_1 U9411 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [18]), .op(n7805)
         );
  nand2_1 U9412 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [18]), .op(n7804)
         );
  nand2_1 U9413 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [18]), .op(n7803)
         );
  nand2_1 U9414 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [18]), .op(n7809)
         );
  nand2_1 U9415 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [18]), .op(n7808)
         );
  nand2_1 U9416 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [18]), .op(n7807)
         );
  nand3_1 U9417 ( .ip1(n7809), .ip2(n7808), .ip3(n7807), .op(n7810) );
  not_ab_or_c_or_d U9418 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [18]), 
        .ip3(n7811), .ip4(n7810), .op(n7814) );
  nand2_1 U9419 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [16]), .op(n7813)
         );
  nand2_1 U9420 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [16]), .op(n7812)
         );
  not_ab_or_c_or_d U9421 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [18]), 
        .ip3(n7817), .ip4(n7816), .op(n12670) );
  nor2_1 U9422 ( .ip1(n12670), .ip2(n7887), .op(n7818) );
  not_ab_or_c_or_d U9423 ( .ip1(\CORTEXM0DS_INST/u_logic/Ks9vx4 ), .ip2(n7889), 
        .ip3(n7937), .ip4(n7818), .op(n7819) );
  mux2_1 U9424 ( .ip1(n7941), .ip2(n7940), .s(n7819), .op(n9594) );
  nand2_1 U9425 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [19]), .op(n7822)
         );
  nand2_1 U9426 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [19]), .op(n7821)
         );
  nand2_1 U9427 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [19]), .op(n7820)
         );
  nand3_1 U9428 ( .ip1(n7822), .ip2(n7821), .ip3(n7820), .op(n7840) );
  nand2_1 U9429 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [19]), .ip2(n9308), .op(n7838)
         );
  nand2_1 U9430 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [19]), .op(n7826)
         );
  nand2_1 U9431 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [19]), .op(n7825)
         );
  nand2_1 U9432 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [19]), .op(n7824)
         );
  nand2_1 U9433 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [19]), .op(n7823)
         );
  nand2_1 U9434 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [17]), .op(n7830)
         );
  nand2_1 U9435 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [17]), .op(n7829)
         );
  nand2_1 U9436 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [19]), .op(n7828)
         );
  nand2_1 U9437 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [19]), .op(n7827)
         );
  not_ab_or_c_or_d U9438 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [19]), 
        .ip3(n7832), .ip4(n7831), .op(n7837) );
  nor2_1 U9439 ( .ip1(n7857), .ip2(n7833), .op(n7835) );
  inv_1 U9440 ( .ip(\CORTEXM0DS_INST/u_logic/Bpdvx4 ), .op(n12247) );
  nor2_1 U9441 ( .ip1(n9279), .ip2(n12247), .op(n7834) );
  not_ab_or_c_or_d U9442 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [19]), .ip2(n9309), 
        .ip3(n7835), .ip4(n7834), .op(n7836) );
  nand3_1 U9443 ( .ip1(n7838), .ip2(n7837), .ip3(n7836), .op(n7839) );
  not_ab_or_c_or_d U9444 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [19]), 
        .ip3(n7840), .ip4(n7839), .op(n11382) );
  nor2_1 U9445 ( .ip1(n11382), .ip2(n7887), .op(n7841) );
  not_ab_or_c_or_d U9446 ( .ip1(\CORTEXM0DS_INST/u_logic/Ot9vx4 ), .ip2(n7889), 
        .ip3(n7937), .ip4(n7841), .op(n7842) );
  mux2_1 U9447 ( .ip1(n7941), .ip2(n7940), .s(n7842), .op(n11385) );
  nand2_1 U9448 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [20]), .op(n7845)
         );
  nand2_1 U9449 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [20]), .op(n7844)
         );
  nand2_1 U9450 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [20]), .op(n7843)
         );
  nand3_1 U9451 ( .ip1(n7845), .ip2(n7844), .ip3(n7843), .op(n7864) );
  nand2_1 U9452 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [20]), .ip2(n9308), .op(n7862)
         );
  nand2_1 U9453 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [20]), .op(n7849)
         );
  nand2_1 U9454 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [20]), .op(n7848)
         );
  nand2_1 U9455 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [20]), .op(n7847)
         );
  nand2_1 U9456 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [20]), .op(n7846)
         );
  nand2_1 U9457 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [18]), .op(n7853)
         );
  nand2_1 U9458 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [18]), .op(n7852)
         );
  nand2_1 U9459 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [20]), .op(n7851)
         );
  nand2_1 U9460 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [20]), .op(n7850)
         );
  not_ab_or_c_or_d U9461 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [20]), 
        .ip3(n7855), .ip4(n7854), .op(n7861) );
  nor2_1 U9462 ( .ip1(n7857), .ip2(n7856), .op(n7859) );
  inv_1 U9463 ( .ip(\CORTEXM0DS_INST/u_logic/Mqdvx4 ), .op(n12256) );
  nor2_1 U9464 ( .ip1(n9279), .ip2(n12256), .op(n7858) );
  not_ab_or_c_or_d U9465 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [20]), .ip2(n9326), 
        .ip3(n7859), .ip4(n7858), .op(n7860) );
  nand3_1 U9466 ( .ip1(n7862), .ip2(n7861), .ip3(n7860), .op(n7863) );
  not_ab_or_c_or_d U9467 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [20]), 
        .ip3(n7864), .ip4(n7863), .op(n12674) );
  nor2_1 U9468 ( .ip1(n12674), .ip2(n7887), .op(n7865) );
  not_ab_or_c_or_d U9469 ( .ip1(\CORTEXM0DS_INST/u_logic/Su9vx4 ), .ip2(n7889), 
        .ip3(n7937), .ip4(n7865), .op(n7866) );
  mux2_1 U9470 ( .ip1(n7941), .ip2(n7940), .s(n7866), .op(n9591) );
  nand2_1 U9471 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [21]), .op(n7869)
         );
  nand2_1 U9472 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [21]), .op(n7868)
         );
  nand2_1 U9473 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [21]), .op(n7867)
         );
  nand3_1 U9474 ( .ip1(n7869), .ip2(n7868), .ip3(n7867), .op(n7886) );
  nand2_1 U9475 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [21]), .ip2(n9315), .op(n7884)
         );
  nand2_1 U9476 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [21]), .op(n7873)
         );
  nand2_1 U9477 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [21]), .op(n7872)
         );
  nand2_1 U9478 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [21]), .op(n7871)
         );
  nand2_1 U9479 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [21]), .op(n7870)
         );
  nand2_1 U9480 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [19]), .op(n7877)
         );
  nand2_1 U9481 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [19]), .op(n7876)
         );
  nand2_1 U9482 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [21]), .op(n7875)
         );
  nand2_1 U9483 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [21]), .op(n7874)
         );
  not_ab_or_c_or_d U9484 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [21]), 
        .ip3(n7879), .ip4(n7878), .op(n7883) );
  nor2_1 U9485 ( .ip1(n9279), .ip2(n12267), .op(n7881) );
  and2_1 U9486 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [21]), .op(n7880)
         );
  not_ab_or_c_or_d U9487 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [21]), .ip2(n9314), 
        .ip3(n7881), .ip4(n7880), .op(n7882) );
  nand3_1 U9488 ( .ip1(n7884), .ip2(n7883), .ip3(n7882), .op(n7885) );
  not_ab_or_c_or_d U9489 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [21]), 
        .ip3(n7886), .ip4(n7885), .op(n9580) );
  nor2_1 U9490 ( .ip1(n9580), .ip2(n7887), .op(n7888) );
  not_ab_or_c_or_d U9491 ( .ip1(\CORTEXM0DS_INST/u_logic/Wv9vx4 ), .ip2(n7889), 
        .ip3(n7937), .ip4(n7888), .op(n7890) );
  mux2_1 U9492 ( .ip1(n7941), .ip2(n7940), .s(n7890), .op(n11405) );
  nand2_1 U9493 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [22]), .op(n7894)
         );
  nand2_1 U9494 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [22]), .op(n7893)
         );
  nand2_1 U9495 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [22]), .op(n7892)
         );
  nand2_1 U9496 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [22]), .op(n7891)
         );
  and4_1 U9497 ( .ip1(n7894), .ip2(n7893), .ip3(n7892), .ip4(n7891), .op(n7910) );
  inv_1 U9498 ( .ip(\CORTEXM0DS_INST/u_logic/Itdvx4 ), .op(n12277) );
  nor2_1 U9499 ( .ip1(n9279), .ip2(n12277), .op(n7896) );
  and2_1 U9500 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [22]), .op(n7895)
         );
  not_ab_or_c_or_d U9501 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [22]), .ip2(n9338), 
        .ip3(n7896), .ip4(n7895), .op(n7909) );
  nand2_1 U9502 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [22]), .op(n7900)
         );
  nand2_1 U9503 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [22]), .op(n7899)
         );
  nand2_1 U9504 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [22]), .op(n7898)
         );
  nand2_1 U9505 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [22]), .op(n7897)
         );
  nand2_1 U9506 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [20]), .op(n7904)
         );
  nand2_1 U9507 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [20]), .op(n7903)
         );
  nand2_1 U9508 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [22]), .op(n7902)
         );
  nand2_1 U9509 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [22]), .op(n7901)
         );
  not_ab_or_c_or_d U9510 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [22]), 
        .ip3(n7906), .ip4(n7905), .op(n7908) );
  nand2_1 U9511 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [22]), .op(n7907)
         );
  nor2_1 U9512 ( .ip1(n12384), .ip2(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .op(
        n7911) );
  not_ab_or_c_or_d U9513 ( .ip1(n12384), .ip2(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip3(n7911), .ip4(n7935), .op(n7912) );
  not_ab_or_c_or_d U9514 ( .ip1(n7938), .ip2(n12680), .ip3(n7937), .ip4(n7912), 
        .op(n7913) );
  mux2_1 U9515 ( .ip1(n7941), .ip2(n7940), .s(n7913), .op(n9597) );
  nand2_1 U9516 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [23]), .op(n7917)
         );
  nand2_1 U9517 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [23]), .op(n7916)
         );
  nand2_1 U9518 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [23]), .op(n7915)
         );
  nand2_1 U9519 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [23]), .op(n7914)
         );
  and4_1 U9520 ( .ip1(n7917), .ip2(n7916), .ip3(n7915), .ip4(n7914), .op(n7933) );
  and2_1 U9521 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [23]), .op(n7919)
         );
  nor2_1 U9522 ( .ip1(n9279), .ip2(n12149), .op(n7918) );
  not_ab_or_c_or_d U9523 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [23]), .ip2(n9308), 
        .ip3(n7919), .ip4(n7918), .op(n7932) );
  nand2_1 U9524 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [23]), .op(n7923)
         );
  nand2_1 U9525 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [23]), .op(n7922)
         );
  nand2_1 U9526 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [23]), .op(n7921)
         );
  nand2_1 U9527 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [23]), .op(n7920)
         );
  nand2_1 U9528 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [21]), .op(n7927)
         );
  nand2_1 U9529 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [21]), .op(n7926)
         );
  nand2_1 U9530 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [23]), .op(n7925)
         );
  nand2_1 U9531 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [23]), .op(n7924)
         );
  not_ab_or_c_or_d U9532 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [23]), 
        .ip3(n7929), .ip4(n7928), .op(n7931) );
  nand2_1 U9533 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [23]), .op(n7930)
         );
  nor2_1 U9534 ( .ip1(\CORTEXM0DS_INST/u_logic/Bx9vx4 ), .ip2(n12538), .op(
        n7934) );
  not_ab_or_c_or_d U9535 ( .ip1(\CORTEXM0DS_INST/u_logic/Bx9vx4 ), .ip2(n12538), .ip3(n7935), .ip4(n7934), .op(n7936) );
  not_ab_or_c_or_d U9536 ( .ip1(n7938), .ip2(n12682), .ip3(n7937), .ip4(n7936), 
        .op(n7939) );
  mux2_1 U9537 ( .ip1(n7941), .ip2(n7940), .s(n7939), .op(n9536) );
  nand2_1 U9538 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [24]), .op(n7944)
         );
  nand2_1 U9539 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [24]), .op(n7943)
         );
  nand2_1 U9540 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [24]), .op(n7942)
         );
  nand3_1 U9541 ( .ip1(n7944), .ip2(n7943), .ip3(n7942), .op(n7963) );
  nand2_1 U9542 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [24]), .ip2(n9344), .op(n7961)
         );
  nand2_1 U9543 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [24]), .op(n7948)
         );
  nand2_1 U9544 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [24]), .op(n7947)
         );
  nand2_1 U9545 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [24]), .op(n7946)
         );
  nand2_1 U9546 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [24]), .op(n7945)
         );
  nand2_1 U9547 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [22]), .op(n7952)
         );
  nand2_1 U9548 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [22]), .op(n7951)
         );
  nand2_1 U9549 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [24]), .op(n7950)
         );
  nand2_1 U9550 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [24]), .op(n7949)
         );
  not_ab_or_c_or_d U9551 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [24]), 
        .ip3(n7954), .ip4(n7953), .op(n7960) );
  nor2_1 U9552 ( .ip1(n7956), .ip2(n7955), .op(n7958) );
  nor2_1 U9553 ( .ip1(n9279), .ip2(n12354), .op(n7957) );
  not_ab_or_c_or_d U9554 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [24]), 
        .ip3(n7958), .ip4(n7957), .op(n7959) );
  nand3_1 U9555 ( .ip1(n7961), .ip2(n7960), .ip3(n7959), .op(n7962) );
  not_ab_or_c_or_d U9556 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [24]), 
        .ip3(n7963), .ip4(n7962), .op(n11455) );
  mux2_1 U9557 ( .ip1(n9346), .ip2(n9345), .s(n11455), .op(n9623) );
  nor2_1 U9558 ( .ip1(n9371), .ip2(n7964), .op(n7965) );
  xor2_1 U9559 ( .ip1(n11471), .ip2(n7965), .op(n8049) );
  nand2_1 U9560 ( .ip1(n8050), .ip2(n8049), .op(n7966) );
  nand2_1 U9561 ( .ip1(n7967), .ip2(n7966), .op(n7994) );
  nand2_1 U9562 ( .ip1(n7993), .ip2(n7994), .op(n7968) );
  nand2_1 U9563 ( .ip1(n7969), .ip2(n7968), .op(n8539) );
  nand2_1 U9564 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [28]), .op(n7972)
         );
  nand2_1 U9565 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [28]), .op(n7971)
         );
  nand2_1 U9566 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [28]), .op(n7970)
         );
  nand3_1 U9567 ( .ip1(n7972), .ip2(n7971), .ip3(n7970), .op(n7989) );
  and2_1 U9568 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [26]), .op(n7974)
         );
  nor2_1 U9569 ( .ip1(n9279), .ip2(n8564), .op(n7973) );
  not_ab_or_c_or_d U9570 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [28]), .ip2(n9316), 
        .ip3(n7974), .ip4(n7973), .op(n7987) );
  nand2_1 U9571 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [28]), .op(n7978)
         );
  nand2_1 U9572 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [28]), .op(n7977)
         );
  nand2_1 U9573 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [28]), .op(n7976)
         );
  nand2_1 U9574 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [28]), .op(n7975)
         );
  nand2_1 U9575 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [28]), .op(n7981)
         );
  nand2_1 U9576 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [28]), .op(n7980)
         );
  nand2_1 U9577 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [28]), .op(n7979)
         );
  nand3_1 U9578 ( .ip1(n7981), .ip2(n7980), .ip3(n7979), .op(n7982) );
  not_ab_or_c_or_d U9579 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [28]), 
        .ip3(n7983), .ip4(n7982), .op(n7986) );
  nand2_1 U9580 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [26]), .op(n7985)
         );
  nand2_1 U9581 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [28]), .op(n7984)
         );
  not_ab_or_c_or_d U9582 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [28]), 
        .ip3(n7989), .ip4(n7988), .op(n11052) );
  mux2_1 U9583 ( .ip1(n8562), .ip2(n8563), .s(n11052), .op(n9514) );
  inv_1 U9584 ( .ip(n9513), .op(n9516) );
  nor2_1 U9585 ( .ip1(n9514), .ip2(n9516), .op(n9520) );
  and2_1 U9586 ( .ip1(n9261), .ip2(n9520), .op(n8538) );
  nand2_1 U9587 ( .ip1(n9261), .ip2(n9513), .op(n7990) );
  nand2_1 U9588 ( .ip1(n9514), .ip2(n7990), .op(n8541) );
  inv_1 U9589 ( .ip(n8541), .op(n7991) );
  nor2_1 U9590 ( .ip1(n8538), .ip2(n7991), .op(n7992) );
  xor2_1 U9591 ( .ip1(n8539), .ip2(n7992), .op(n8535) );
  xor2_1 U9592 ( .ip1(n7994), .ip2(n7993), .op(n9436) );
  fulladder U9593 ( .a(n7996), .b(n9542), .ci(n7995), .co(n8050), .s(n9439) );
  fulladder U9594 ( .a(n7998), .b(n7997), .ci(n9623), .co(n7995), .s(n9412) );
  fulladder U9595 ( .a(n8000), .b(n7999), .ci(n9536), .co(n7997), .s(n9648) );
  fulladder U9596 ( .a(n8002), .b(n8001), .ci(n9597), .co(n7999), .s(n8898) );
  fulladder U9597 ( .a(n8004), .b(n8003), .ci(n11405), .co(n8001), .s(n9441)
         );
  inv_1 U9598 ( .ip(n9441), .op(n8047) );
  fulladder U9599 ( .a(n8006), .b(n8005), .ci(n9591), .co(n8003), .s(n9428) );
  fulladder U9600 ( .a(n8008), .b(n8007), .ci(n11385), .co(n8005), .s(n9640)
         );
  fulladder U9601 ( .a(n8010), .b(n8009), .ci(n9594), .co(n8007), .s(n9430) );
  inv_1 U9602 ( .ip(n9430), .op(n8046) );
  fulladder U9603 ( .a(n8012), .b(n8011), .ci(n11362), .co(n8009), .s(n9432)
         );
  fulladder U9604 ( .a(n8014), .b(n8013), .ci(n9596), .co(n8011), .s(n8840) );
  fulladder U9605 ( .a(n8016), .b(n8015), .ci(n9593), .co(n8013), .s(n9421) );
  fulladder U9606 ( .a(n8018), .b(n8017), .ci(n9620), .co(n8015), .s(n9423) );
  fulladder U9607 ( .a(n8020), .b(n8019), .ci(n9616), .co(n8017), .s(n9419) );
  fulladder U9608 ( .a(n8022), .b(n8021), .ci(n9497), .co(n8041), .s(n9642) );
  fulladder U9609 ( .a(n8024), .b(n8023), .ci(n9466), .co(n8021), .s(n8406) );
  fulladder U9610 ( .a(n8026), .b(n8025), .ci(n11559), .co(n8023), .s(n9414)
         );
  inv_1 U9611 ( .ip(n9414), .op(n8040) );
  fulladder U9612 ( .a(n8028), .b(n8027), .ci(n9447), .co(n8025), .s(n8845) );
  fulladder U9613 ( .a(n8030), .b(n8029), .ci(n9611), .co(n8027), .s(n8633) );
  inv_1 U9614 ( .ip(n8633), .op(n8039) );
  fulladder U9615 ( .a(n8032), .b(n8031), .ci(n9463), .co(n8029), .s(n8883) );
  fulladder U9616 ( .a(n8034), .b(n8033), .ci(n9566), .co(n8031), .s(n8870) );
  inv_1 U9617 ( .ip(n8035), .op(n8037) );
  nor2_1 U9618 ( .ip1(n8037), .ip2(n8036), .op(n8869) );
  nand2_1 U9619 ( .ip1(n8870), .ip2(n8869), .op(n8882) );
  inv_1 U9620 ( .ip(n8882), .op(n8038) );
  nand2_1 U9621 ( .ip1(n8883), .ip2(n8038), .op(n8632) );
  nor2_1 U9622 ( .ip1(n8039), .ip2(n8632), .op(n8844) );
  nand2_1 U9623 ( .ip1(n8845), .ip2(n8844), .op(n9413) );
  nor2_1 U9624 ( .ip1(n8040), .ip2(n9413), .op(n8405) );
  and2_1 U9625 ( .ip1(n8406), .ip2(n8405), .op(n9641) );
  nand2_1 U9626 ( .ip1(n9642), .ip2(n9641), .op(n8400) );
  fulladder U9627 ( .a(n8042), .b(n8041), .ci(n9618), .co(n8044), .s(n8401) );
  inv_1 U9628 ( .ip(n8401), .op(n8043) );
  nor2_1 U9629 ( .ip1(n8400), .ip2(n8043), .op(n9416) );
  fulladder U9630 ( .a(n8045), .b(n8044), .ci(n9592), .co(n8019), .s(n9417) );
  and2_1 U9631 ( .ip1(n9416), .ip2(n9417), .op(n9418) );
  and2_1 U9632 ( .ip1(n9419), .ip2(n9418), .op(n9422) );
  and2_1 U9633 ( .ip1(n9423), .ip2(n9422), .op(n9420) );
  and2_1 U9634 ( .ip1(n9421), .ip2(n9420), .op(n8839) );
  and2_1 U9635 ( .ip1(n8840), .ip2(n8839), .op(n9431) );
  nand2_1 U9636 ( .ip1(n9432), .ip2(n9431), .op(n9429) );
  nor2_1 U9637 ( .ip1(n8046), .ip2(n9429), .op(n9639) );
  and2_1 U9638 ( .ip1(n9640), .ip2(n9639), .op(n9427) );
  nand2_1 U9639 ( .ip1(n9428), .ip2(n9427), .op(n9440) );
  nor2_1 U9640 ( .ip1(n8047), .ip2(n9440), .op(n8897) );
  and2_1 U9641 ( .ip1(n8898), .ip2(n8897), .op(n9647) );
  and2_1 U9642 ( .ip1(n9648), .ip2(n9647), .op(n9411) );
  nand2_1 U9643 ( .ip1(n9412), .ip2(n9411), .op(n9438) );
  inv_1 U9644 ( .ip(n9438), .op(n8048) );
  nand2_1 U9645 ( .ip1(n9439), .ip2(n8048), .op(n9409) );
  xor2_1 U9646 ( .ip1(n8050), .ip2(n8049), .op(n9410) );
  inv_1 U9647 ( .ip(n9410), .op(n8051) );
  nor2_1 U9648 ( .ip1(n9409), .ip2(n8051), .op(n9437) );
  nand2_1 U9649 ( .ip1(n9436), .ip2(n9437), .op(n8537) );
  xor2_1 U9650 ( .ip1(n8535), .ip2(n8537), .op(n10232) );
  nor2_1 U9651 ( .ip1(n10232), .ip2(n12311), .op(n8052) );
  not_ab_or_c_or_d U9652 ( .ip1(n12316), .ip2(n9513), .ip3(n8053), .ip4(n8052), 
        .op(\CORTEXM0DS_INST/u_logic/V2qvx4 ) );
  or2_1 U9653 ( .ip1(n12355), .ip2(\CORTEXM0DS_INST/u_logic/V2qvx4 ), .op(
        n8054) );
  nand4_1 U9654 ( .ip1(n8057), .ip2(n8056), .ip3(n8055), .ip4(n8054), .op(
        n6073) );
  nand2_1 U9655 ( .ip1(\CORTEXM0DS_INST/u_logic/Ho8vx4 ), .ip2(n12575), .op(
        n8061) );
  nand3_1 U9656 ( .ip1(\CORTEXM0DS_INST/u_logic/Xyfvx4 ), .ip2(n12600), .ip3(
        n12660), .op(n8060) );
  nand2_1 U9657 ( .ip1(\CORTEXM0DS_INST/u_logic/R9fvx4 ), .ip2(n12598), .op(
        n8059) );
  nand2_1 U9658 ( .ip1(n12603), .ip2(\CORTEXM0DS_INST/u_logic/Mxfvx4 ), .op(
        n8058) );
  nand4_1 U9659 ( .ip1(n8061), .ip2(n8060), .ip3(n8059), .ip4(n8058), .op(
        \CORTEXM0DS_INST/u_logic/Llnvx4 ) );
  inv_1 U9660 ( .ip(n5814), .op(n10414) );
  nand2_1 U9661 ( .ip1(n10414), .ip2(n11061), .op(n10912) );
  inv_1 U9662 ( .ip(n8062), .op(n11059) );
  nor2_1 U9663 ( .ip1(n5814), .ip2(n11059), .op(n10916) );
  inv_1 U9664 ( .ip(n10916), .op(n10383) );
  nand2_1 U9665 ( .ip1(n10912), .ip2(n10383), .op(n10901) );
  inv_1 U9666 ( .ip(n10901), .op(n12113) );
  nand3_1 U9667 ( .ip1(\CORTEXM0DS_INST/vis_pc [2]), .ip2(
        \CORTEXM0DS_INST/vis_pc [3]), .ip3(\CORTEXM0DS_INST/vis_pc [4]), .op(
        n8635) );
  nand2_1 U9668 ( .ip1(\CORTEXM0DS_INST/vis_pc [0]), .ip2(
        \CORTEXM0DS_INST/vis_pc [1]), .op(n8586) );
  nand2_1 U9669 ( .ip1(\CORTEXM0DS_INST/vis_pc [5]), .ip2(
        \CORTEXM0DS_INST/vis_pc [6]), .op(n8063) );
  nor4_1 U9670 ( .ip1(n12154), .ip2(n8635), .ip3(n8586), .ip4(n8063), .op(
        n8532) );
  nand3_1 U9671 ( .ip1(n12113), .ip2(n8532), .ip3(n10414), .op(n10344) );
  nor2_1 U9672 ( .ip1(n8064), .ip2(n10344), .op(n10338) );
  inv_1 U9673 ( .ip(n10338), .op(n10192) );
  nand2_1 U9674 ( .ip1(n12113), .ip2(n10192), .op(n10345) );
  mux2_1 U9675 ( .ip1(n10192), .ip2(n10345), .s(\CORTEXM0DS_INST/vis_pc [10]), 
        .op(n8404) );
  nor2_1 U9676 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [0]), .ip2(n8942), .op(n12410)
         );
  and3_1 U9677 ( .ip1(n12403), .ip2(n12402), .ip3(
        \CORTEXM0DS_INST/u_logic/Mk8vx4 ), .op(n8066) );
  inv_1 U9678 ( .ip(n8065), .op(LOCKUP_top_out) );
  not_ab_or_c_or_d U9679 ( .ip1(\CORTEXM0DS_INST/u_logic/Ul8vx4 ), .ip2(n12410), .ip3(n8066), .ip4(LOCKUP_top_out), .op(n8067) );
  nor2_1 U9680 ( .ip1(n5814), .ip2(n8067), .op(n10467) );
  inv_1 U9681 ( .ip(n10467), .op(n10917) );
  inv_1 U9682 ( .ip(n10912), .op(n10475) );
  nor2_1 U9683 ( .ip1(n10851), .ip2(n10740), .op(n10992) );
  inv_1 U9684 ( .ip(n12618), .op(n12124) );
  nor3_1 U9685 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n12124), .ip3(
        n11693), .op(n8960) );
  nor4_1 U9686 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip3(n12117), .ip4(n12609), .op(
        n8377) );
  nor4_1 U9687 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n10992), .ip3(
        n8960), .ip4(n8377), .op(n8747) );
  inv_1 U9688 ( .ip(\CORTEXM0DS_INST/u_logic/Dw8vx4 ), .op(n9712) );
  nor2_1 U9689 ( .ip1(n8747), .ip2(n9712), .op(n8714) );
  inv_1 U9690 ( .ip(n8714), .op(n11871) );
  inv_1 U9691 ( .ip(\CORTEXM0DS_INST/u_logic/L9hvx4 ), .op(n11901) );
  inv_1 U9692 ( .ip(\CORTEXM0DS_INST/u_logic/B5hvx4 ), .op(n12433) );
  nand4_1 U9693 ( .ip1(n9146), .ip2(n11901), .ip3(n12433), .ip4(
        \CORTEXM0DS_INST/u_logic/N6hvx4 ), .op(n11899) );
  nor2_1 U9694 ( .ip1(n11871), .ip2(n11899), .op(n11829) );
  inv_1 U9695 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [11]), .op(n11727) );
  nand2_1 U9696 ( .ip1(\CORTEXM0DS_INST/u_logic/N6hvx4 ), .ip2(n11903), .op(
        n11860) );
  nor2_1 U9697 ( .ip1(n11871), .ip2(n11860), .op(n10272) );
  inv_1 U9698 ( .ip(n10272), .op(n11830) );
  nor2_1 U9699 ( .ip1(n11727), .ip2(n11830), .op(n8096) );
  nor2_1 U9700 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .op(n10653) );
  nor2_1 U9701 ( .ip1(n10653), .ip2(n12609), .op(n8605) );
  inv_1 U9702 ( .ip(n9377), .op(n11679) );
  nor3_1 U9703 ( .ip1(n8605), .ip2(n12133), .ip3(n11679), .op(n8068) );
  nor2_1 U9704 ( .ip1(n8068), .ip2(n9712), .op(n11853) );
  inv_1 U9705 ( .ip(n11853), .op(n11660) );
  nor2_1 U9706 ( .ip1(n9712), .ip2(n9751), .op(n8121) );
  nand2_1 U9707 ( .ip1(\CORTEXM0DS_INST/u_logic/Dw8vx4 ), .ip2(n11275), .op(
        n8114) );
  nor2_1 U9708 ( .ip1(n8069), .ip2(n8114), .op(n8070) );
  or2_1 U9709 ( .ip1(n8121), .ip2(n8070), .op(n8073) );
  or2_1 U9710 ( .ip1(n8071), .ip2(n8070), .op(n8072) );
  nand2_1 U9711 ( .ip1(n8073), .ip2(n8072), .op(n8079) );
  nor2_1 U9712 ( .ip1(n11517), .ip2(n8114), .op(n8074) );
  or2_1 U9713 ( .ip1(n8121), .ip2(n8074), .op(n8077) );
  or2_1 U9714 ( .ip1(n8075), .ip2(n8074), .op(n8076) );
  nand2_1 U9715 ( .ip1(n8077), .ip2(n8076), .op(n8081) );
  nor2_1 U9716 ( .ip1(n8081), .ip2(n11796), .op(n8078) );
  xor2_1 U9717 ( .ip1(n8079), .ip2(n8078), .op(n9228) );
  inv_1 U9718 ( .ip(n8081), .op(n8080) );
  nand2_1 U9719 ( .ip1(n9228), .ip2(n8080), .op(n9158) );
  inv_1 U9720 ( .ip(n9158), .op(n9179) );
  and2_1 U9721 ( .ip1(n8822), .ip2(n9179), .op(n8085) );
  inv_1 U9722 ( .ip(n8718), .op(n9150) );
  nand2_1 U9723 ( .ip1(n8079), .ip2(n8081), .op(n9243) );
  nor2_1 U9724 ( .ip1(n9150), .ip2(n9243), .op(n8084) );
  nor2_1 U9725 ( .ip1(n8080), .ip2(n8079), .op(n9183) );
  inv_1 U9726 ( .ip(n9183), .op(n9156) );
  nor2_1 U9727 ( .ip1(n8408), .ip2(n9156), .op(n8083) );
  nor2_1 U9728 ( .ip1(n8081), .ip2(n9228), .op(n9185) );
  inv_1 U9729 ( .ip(n9185), .op(n9160) );
  nor2_1 U9730 ( .ip1(n8821), .ip2(n9160), .op(n8082) );
  nor4_1 U9731 ( .ip1(n8085), .ip2(n8084), .ip3(n8083), .ip4(n8082), .op(n9168) );
  nor2_1 U9732 ( .ip1(n9161), .ip2(n9243), .op(n8089) );
  nor2_1 U9733 ( .ip1(n9149), .ip2(n9156), .op(n8088) );
  inv_1 U9734 ( .ip(n8690), .op(n9148) );
  nor2_1 U9735 ( .ip1(n9148), .ip2(n9158), .op(n8087) );
  nor2_1 U9736 ( .ip1(n9147), .ip2(n9160), .op(n8086) );
  nor4_1 U9737 ( .ip1(n8089), .ip2(n8088), .ip3(n8087), .ip4(n8086), .op(n9225) );
  or2_1 U9738 ( .ip1(n8114), .ip2(n10942), .op(n8092) );
  nand2_1 U9739 ( .ip1(n8121), .ip2(n8090), .op(n8091) );
  nand2_1 U9740 ( .ip1(n8092), .ip2(n8091), .op(n8111) );
  inv_1 U9741 ( .ip(n9243), .op(n9181) );
  nor2_1 U9742 ( .ip1(n9181), .ip2(n11796), .op(n8093) );
  xor2_1 U9743 ( .ip1(n8111), .ip2(n8093), .op(n8781) );
  inv_1 U9744 ( .ip(n8781), .op(n10256) );
  mux2_1 U9745 ( .ip1(n9168), .ip2(n9225), .s(n10256), .op(n8094) );
  nor2_1 U9746 ( .ip1(n11660), .ip2(n8094), .op(n8095) );
  not_ab_or_c_or_d U9747 ( .ip1(n11829), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [11]), .ip3(n8096), .ip4(n8095), .op(
        n8099) );
  nor2_1 U9748 ( .ip1(\CORTEXM0DS_INST/u_logic/N6hvx4 ), .ip2(n11898), .op(
        n8651) );
  nand2_1 U9749 ( .ip1(n11903), .ip2(n8651), .op(n8906) );
  nor2_1 U9750 ( .ip1(n11871), .ip2(n8906), .op(n10270) );
  nand2_1 U9751 ( .ip1(n10270), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [11]), 
        .op(n8098) );
  nor2_1 U9752 ( .ip1(\CORTEXM0DS_INST/u_logic/N6hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Xahvx4 ), .op(n11902) );
  inv_1 U9753 ( .ip(n11902), .op(n12689) );
  nor4_1 U9754 ( .ip1(n12689), .ip2(n11901), .ip3(n9146), .ip4(n12433), .op(
        n8746) );
  nand2_1 U9755 ( .ip1(n8714), .ip2(n8746), .op(n11875) );
  inv_1 U9756 ( .ip(n11875), .op(n10271) );
  nand2_1 U9757 ( .ip1(n10271), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [11]), 
        .op(n8097) );
  nand4_1 U9758 ( .ip1(n4190), .ip2(n8099), .ip3(n8098), .ip4(n8097), .op(
        n10436) );
  inv_1 U9759 ( .ip(n9956), .op(n11219) );
  nand2_1 U9760 ( .ip1(n11219), .ip2(n11228), .op(n10562) );
  inv_1 U9761 ( .ip(\CORTEXM0DS_INST/u_logic/Zph2z4 [1]), .op(n8614) );
  nor2_1 U9762 ( .ip1(n10478), .ip2(n8614), .op(n8101) );
  nor2_1 U9763 ( .ip1(n12125), .ip2(n10851), .op(n8944) );
  nor2_1 U9764 ( .ip1(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip2(n11693), .op(
        n8100) );
  nor2_1 U9765 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n8100), .op(
        n10872) );
  nor2_1 U9766 ( .ip1(n8944), .ip2(n10872), .op(n8613) );
  inv_1 U9767 ( .ip(n8613), .op(n8592) );
  ab_or_c_or_d U9768 ( .ip1(n10533), .ip2(n10562), .ip3(n8101), .ip4(n8592), 
        .op(n8127) );
  nor3_1 U9769 ( .ip1(n8592), .ip2(n8424), .ip3(n8494), .op(n8126) );
  nand2_1 U9770 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n12609), .op(
        n11067) );
  nand3_1 U9771 ( .ip1(n11067), .ip2(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Vdgvx4 ), .op(n8102) );
  nand2_1 U9772 ( .ip1(n8613), .ip2(n8102), .op(n8485) );
  nor2_1 U9773 ( .ip1(n12104), .ip2(n8114), .op(n8103) );
  or2_1 U9774 ( .ip1(n8121), .ip2(n8103), .op(n8106) );
  or2_1 U9775 ( .ip1(n8104), .ip2(n8103), .op(n8105) );
  nand2_1 U9776 ( .ip1(n8106), .ip2(n8105), .op(n8140) );
  inv_1 U9777 ( .ip(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .op(n11084) );
  nor2_1 U9778 ( .ip1(n8114), .ip2(n11084), .op(n8107) );
  or2_1 U9779 ( .ip1(n8121), .ip2(n8107), .op(n8110) );
  or2_1 U9780 ( .ip1(n8108), .ip2(n8107), .op(n8109) );
  nand2_1 U9781 ( .ip1(n8110), .ip2(n8109), .op(n8124) );
  nor2_1 U9782 ( .ip1(n9243), .ip2(n8111), .op(n8122) );
  and2_1 U9783 ( .ip1(n8124), .ip2(n8122), .op(n8125) );
  nand2_1 U9784 ( .ip1(n8140), .ip2(n8125), .op(n9704) );
  nand2_1 U9785 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n9704), .op(
        n9211) );
  inv_1 U9786 ( .ip(n9211), .op(n9202) );
  nand3_1 U9787 ( .ip1(n8112), .ip2(n11796), .ip3(n11084), .op(n8113) );
  nor4_1 U9788 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip3(n8114), .ip4(n8113), .op(n8119) );
  inv_1 U9789 ( .ip(n8121), .op(n8118) );
  nor2_1 U9790 ( .ip1(n8116), .ip2(n8115), .op(n8117) );
  nor2_1 U9791 ( .ip1(n8118), .ip2(n8117), .op(n9705) );
  not_ab_or_c_or_d U9792 ( .ip1(n8121), .ip2(n8120), .ip3(n8119), .ip4(n9705), 
        .op(n9707) );
  nor2_1 U9793 ( .ip1(n9707), .ip2(n8424), .op(n9251) );
  nor2_1 U9794 ( .ip1(n8122), .ip2(n11796), .op(n8123) );
  xor2_1 U9795 ( .ip1(n8124), .ip2(n8123), .op(n9673) );
  inv_1 U9796 ( .ip(n9673), .op(n8138) );
  or2_1 U9797 ( .ip1(n8125), .ip2(n11796), .op(n8137) );
  xor2_1 U9798 ( .ip1(n8140), .ip2(n8137), .op(n9672) );
  nor2_1 U9799 ( .ip1(n8138), .ip2(n9672), .op(n9691) );
  inv_1 U9800 ( .ip(n9691), .op(n9213) );
  nor2_1 U9801 ( .ip1(n9251), .ip2(n9213), .op(n9701) );
  nand2_1 U9802 ( .ip1(n9701), .ip2(n8592), .op(n8484) );
  or2_1 U9803 ( .ip1(n9202), .ip2(n8484), .op(n8762) );
  nand2_1 U9804 ( .ip1(n8485), .ip2(n8762), .op(n10439) );
  nor2_1 U9805 ( .ip1(n8126), .ip2(n10439), .op(n8610) );
  nand2_1 U9806 ( .ip1(n8127), .ip2(n8610), .op(n10362) );
  nand2_1 U9807 ( .ip1(n10436), .ip2(n10362), .op(n8399) );
  nor2_1 U9808 ( .ip1(n11689), .ip2(n8592), .op(n8596) );
  inv_1 U9809 ( .ip(n8596), .op(n8809) );
  nor2_1 U9810 ( .ip1(n9251), .ip2(n8613), .op(n8601) );
  inv_1 U9811 ( .ip(n8601), .op(n8594) );
  nor3_1 U9812 ( .ip1(n9673), .ip2(n9672), .ip3(n8594), .op(n8782) );
  nand2_1 U9813 ( .ip1(n8782), .ip2(n9211), .op(n8128) );
  nand2_1 U9814 ( .ip1(n8809), .ip2(n8128), .op(n10370) );
  nand2_1 U9815 ( .ip1(n10271), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [19]), 
        .op(n8136) );
  nand2_1 U9816 ( .ip1(n10270), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [19]), 
        .op(n8135) );
  nor2_1 U9817 ( .ip1(n8781), .ip2(n11660), .op(n10285) );
  nand2_1 U9818 ( .ip1(n9179), .ip2(n8815), .op(n8133) );
  nand2_1 U9819 ( .ip1(n9183), .ip2(n8814), .op(n8132) );
  nand2_1 U9820 ( .ip1(n9181), .ip2(n8824), .op(n8131) );
  inv_1 U9821 ( .ip(n8129), .op(n8816) );
  nand2_1 U9822 ( .ip1(n9185), .ip2(n8816), .op(n8130) );
  nand4_1 U9823 ( .ip1(n8133), .ip2(n8132), .ip3(n8131), .ip4(n8130), .op(
        n9196) );
  nand2_1 U9824 ( .ip1(n10285), .ip2(n9196), .op(n8134) );
  nand4_1 U9825 ( .ip1(n4185), .ip2(n8136), .ip3(n8135), .ip4(n8134), .op(
        n10438) );
  nand2_1 U9826 ( .ip1(n9673), .ip2(n9672), .op(n9670) );
  nand2_1 U9827 ( .ip1(n8140), .ip2(n8137), .op(n8139) );
  nand2_1 U9828 ( .ip1(n9672), .ip2(n8138), .op(n8595) );
  nand2_1 U9829 ( .ip1(n8139), .ip2(n8595), .op(n8600) );
  nor2_1 U9830 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n11256), .op(
        n9214) );
  inv_1 U9831 ( .ip(n9214), .op(n8526) );
  or2_1 U9832 ( .ip1(n8526), .ip2(n8140), .op(n9176) );
  nand2_1 U9833 ( .ip1(n8600), .ip2(n9176), .op(n9201) );
  nand2_1 U9834 ( .ip1(n9670), .ip2(n9201), .op(n9207) );
  nand2_1 U9835 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n11132), .op(
        n8495) );
  inv_1 U9836 ( .ip(n8495), .op(n8142) );
  nor2_1 U9837 ( .ip1(n12609), .ip2(n10944), .op(n8141) );
  nand2_1 U9838 ( .ip1(n8714), .ip2(n12608), .op(n8145) );
  nand2_1 U9839 ( .ip1(n8613), .ip2(n8145), .op(n8604) );
  not_ab_or_c_or_d U9840 ( .ip1(n8142), .ip2(n8424), .ip3(n8141), .ip4(n8604), 
        .op(n8357) );
  or2_1 U9841 ( .ip1(n9377), .ip2(n9349), .op(n8144) );
  nand2_1 U9842 ( .ip1(n11250), .ip2(n11796), .op(n11691) );
  or2_1 U9843 ( .ip1(n11691), .ip2(n9349), .op(n8143) );
  nand2_1 U9844 ( .ip1(n8144), .ip2(n8143), .op(n9256) );
  nand2_1 U9845 ( .ip1(\CORTEXM0DS_INST/u_logic/Dw8vx4 ), .ip2(n9256), .op(
        n9698) );
  inv_1 U9846 ( .ip(n9698), .op(n9247) );
  inv_1 U9847 ( .ip(n8145), .op(n8356) );
  inv_1 U9848 ( .ip(n11755), .op(n10611) );
  or2_1 U9849 ( .ip1(n11786), .ip2(n10611), .op(n8146) );
  inv_1 U9850 ( .ip(\CORTEXM0DS_INST/u_logic/Zph2z4 [0]), .op(n8593) );
  nand2_1 U9851 ( .ip1(n8614), .ip2(n8593), .op(n8606) );
  nand2_1 U9852 ( .ip1(n11224), .ip2(n8606), .op(n8148) );
  nand2_1 U9853 ( .ip1(n8146), .ip2(n8148), .op(n8147) );
  nor2_1 U9854 ( .ip1(n4149), .ip2(n8147), .op(n8355) );
  inv_1 U9855 ( .ip(n8148), .op(n8149) );
  not_ab_or_c_or_d U9856 ( .ip1(\CORTEXM0DS_INST/u_logic/Zph2z4 [1]), .ip2(
        n4130), .ip3(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip4(n9956), .op(n8153) );
  or2_1 U9857 ( .ip1(n8149), .ip2(n8153), .op(n8156) );
  nand2_1 U9858 ( .ip1(n10271), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [23]), 
        .op(n8151) );
  nand2_1 U9859 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [23]), .ip2(n10270), 
        .op(n8150) );
  nand3_1 U9860 ( .ip1(n8151), .ip2(n3020), .ip3(n8150), .op(n10454) );
  nand2_1 U9861 ( .ip1(\CORTEXM0DS_INST/u_logic/Zph2z4 [1]), .ip2(n4130), .op(
        n8152) );
  mux2_1 U9862 ( .ip1(n10454), .ip2(n8152), .s(
        \CORTEXM0DS_INST/u_logic/Zph2z4 [0]), .op(n8154) );
  or2_1 U9863 ( .ip1(n8154), .ip2(n8153), .op(n8155) );
  nand2_1 U9864 ( .ip1(n8156), .ip2(n8155), .op(n8351) );
  nand2_1 U9865 ( .ip1(n8351), .ip2(n8157), .op(n8350) );
  nand2_1 U9866 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [15]), .ip2(n10270), 
        .op(n8349) );
  nand2_1 U9867 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [1]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [1]), .op(n8159) );
  nand2_1 U9868 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [0]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [0]), .op(n8158) );
  nand2_1 U9869 ( .ip1(n8159), .ip2(n8158), .op(n8269) );
  nand2_1 U9870 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [3]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [3]), .op(n8161) );
  nand2_1 U9871 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [2]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [2]), .op(n8160) );
  nand2_1 U9872 ( .ip1(n8161), .ip2(n8160), .op(n8267) );
  nor2_1 U9873 ( .ip1(n8269), .ip2(n8267), .op(n8281) );
  inv_1 U9874 ( .ip(n8281), .op(n8166) );
  nand2_1 U9875 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [5]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [5]), .op(n8163) );
  nand2_1 U9876 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [4]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [4]), .op(n8162) );
  nand2_1 U9877 ( .ip1(n8163), .ip2(n8162), .op(n8250) );
  nand2_1 U9878 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [7]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [7]), .op(n8165) );
  nand2_1 U9879 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [6]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [6]), .op(n8164) );
  nand2_1 U9880 ( .ip1(n8165), .ip2(n8164), .op(n8248) );
  or2_1 U9881 ( .ip1(n8250), .ip2(n8248), .op(n8282) );
  nor2_1 U9882 ( .ip1(n8166), .ip2(n8282), .op(n8302) );
  inv_1 U9883 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [29]), .op(n8168) );
  nor2_1 U9884 ( .ip1(n8168), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [31]), .op(
        n8170) );
  inv_1 U9885 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [28]), .op(n8167) );
  not_ab_or_c_or_d U9886 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [31]), .ip2(
        n8168), .ip3(\CORTEXM0DS_INST/u_logic/Zuh2z4 [30]), .ip4(n8167), .op(
        n8169) );
  or2_1 U9887 ( .ip1(n8170), .ip2(n8169), .op(n8171) );
  nand3_1 U9888 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [15]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [15]), .ip3(n8171), .op(n8172) );
  and3_1 U9889 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [14]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [14]), .ip3(n8172), .op(n10105) );
  mux2_1 U9890 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [31]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [29]), .s(n10105), .op(n8189) );
  inv_1 U9891 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [25]), .op(n11855) );
  nor2_1 U9892 ( .ip1(n11855), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [27]), 
        .op(n8174) );
  not_ab_or_c_or_d U9893 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [27]), .ip2(
        n11855), .ip3(\CORTEXM0DS_INST/u_logic/Zuh2z4 [26]), .ip4(n8181), .op(
        n8173) );
  or2_1 U9894 ( .ip1(n8174), .ip2(n8173), .op(n8175) );
  nand3_1 U9895 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [13]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [13]), .ip3(n8175), .op(n8176) );
  nand3_1 U9896 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [12]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [12]), .ip3(n8176), .op(n10107) );
  mux2_1 U9897 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [25]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [27]), .s(n10107), .op(n8188) );
  nand2_1 U9898 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [15]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [15]), .op(n8178) );
  nand2_1 U9899 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [14]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [14]), .op(n8177) );
  nand2_1 U9900 ( .ip1(n8178), .ip2(n8177), .op(n8215) );
  and2_1 U9901 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [13]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [13]), .op(n8180) );
  and2_1 U9902 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [12]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [12]), .op(n8179) );
  nor2_1 U9903 ( .ip1(n8180), .ip2(n8179), .op(n8221) );
  or2_1 U9904 ( .ip1(n8215), .ip2(n8221), .op(n8187) );
  inv_1 U9905 ( .ip(n8188), .op(n8182) );
  nor2_1 U9906 ( .ip1(n8189), .ip2(n8182), .op(n8184) );
  mux2_1 U9907 ( .ip1(n8181), .ip2(n8739), .s(n10107), .op(n8216) );
  mux2_1 U9908 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [30]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [28]), .s(n10105), .op(n8291) );
  not_ab_or_c_or_d U9909 ( .ip1(n8182), .ip2(n8189), .ip3(n8216), .ip4(n8291), 
        .op(n8183) );
  or2_1 U9910 ( .ip1(n8184), .ip2(n8183), .op(n8185) );
  or2_1 U9911 ( .ip1(n8185), .ip2(n8221), .op(n8186) );
  nand2_1 U9912 ( .ip1(n8187), .ip2(n8186), .op(n10108) );
  mux2_1 U9913 ( .ip1(n8189), .ip2(n8188), .s(n10108), .op(n8230) );
  inv_1 U9914 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [21]), .op(n8191) );
  nor2_1 U9915 ( .ip1(n8191), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [23]), .op(
        n8193) );
  inv_1 U9916 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [20]), .op(n8190) );
  not_ab_or_c_or_d U9917 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [23]), .ip2(
        n8191), .ip3(\CORTEXM0DS_INST/u_logic/Zuh2z4 [22]), .ip4(n8190), .op(
        n8192) );
  or2_1 U9918 ( .ip1(n8193), .ip2(n8192), .op(n8194) );
  nand3_1 U9919 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [11]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [11]), .ip3(n8194), .op(n8195) );
  and3_1 U9920 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [10]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [10]), .ip3(n8195), .op(n10112) );
  mux2_1 U9921 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [23]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [21]), .s(n10112), .op(n8212) );
  nor2_1 U9922 ( .ip1(n8197), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [19]), .op(
        n8199) );
  not_ab_or_c_or_d U9923 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [19]), .ip2(
        n8197), .ip3(\CORTEXM0DS_INST/u_logic/Zuh2z4 [18]), .ip4(n8196), .op(
        n8198) );
  or2_1 U9924 ( .ip1(n8199), .ip2(n8198), .op(n8200) );
  nand3_1 U9925 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [9]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [9]), .ip3(n8200), .op(n8201) );
  and3_1 U9926 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [8]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [8]), .ip3(n8201), .op(n10115) );
  mux2_1 U9927 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [19]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [17]), .s(n10115), .op(n8211) );
  nand2_1 U9928 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [9]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [9]), .op(n8203) );
  nand2_1 U9929 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [8]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [8]), .op(n8202) );
  nand2_1 U9930 ( .ip1(n8203), .ip2(n8202), .op(n8225) );
  nand2_1 U9931 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [11]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [11]), .op(n8205) );
  nand2_1 U9932 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [10]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [10]), .op(n8204) );
  nand2_1 U9933 ( .ip1(n8205), .ip2(n8204), .op(n8224) );
  inv_1 U9934 ( .ip(n8211), .op(n8207) );
  nor2_1 U9935 ( .ip1(n8212), .ip2(n8207), .op(n8209) );
  mux2_1 U9936 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [18]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [16]), .s(n10115), .op(n8213) );
  inv_1 U9937 ( .ip(n8213), .op(n8206) );
  mux2_1 U9938 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [22]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [20]), .s(n10112), .op(n8214) );
  not_ab_or_c_or_d U9939 ( .ip1(n8207), .ip2(n8212), .ip3(n8206), .ip4(n8214), 
        .op(n8208) );
  or2_1 U9940 ( .ip1(n8209), .ip2(n8208), .op(n8210) );
  nand2_1 U9941 ( .ip1(n8224), .ip2(n8210), .op(n10113) );
  and2_1 U9942 ( .ip1(n8225), .ip2(n10113), .op(n8514) );
  mux2_1 U9943 ( .ip1(n8212), .ip2(n8211), .s(n8514), .op(n8229) );
  inv_1 U9944 ( .ip(n8229), .op(n8223) );
  mux2_1 U9945 ( .ip1(n8214), .ip2(n8213), .s(n8514), .op(n8294) );
  inv_1 U9946 ( .ip(n8294), .op(n8219) );
  inv_1 U9947 ( .ip(n8215), .op(n8220) );
  or2_1 U9948 ( .ip1(n8220), .ip2(n8291), .op(n8217) );
  inv_1 U9949 ( .ip(n8216), .op(n8288) );
  mux2_1 U9950 ( .ip1(n8217), .ip2(n8288), .s(n10108), .op(n8218) );
  ab_or_c_or_d U9951 ( .ip1(n8223), .ip2(n8230), .ip3(n8219), .ip4(n8218), 
        .op(n8228) );
  nand2_1 U9952 ( .ip1(n8221), .ip2(n8220), .op(n8287) );
  inv_1 U9953 ( .ip(n8287), .op(n8222) );
  nor3_1 U9954 ( .ip1(n8223), .ip2(n8230), .ip3(n8222), .op(n8227) );
  nor2_1 U9955 ( .ip1(n8225), .ip2(n8224), .op(n8226) );
  nor2_1 U9956 ( .ip1(n8227), .ip2(n8226), .op(n8290) );
  nand2_1 U9957 ( .ip1(n8228), .ip2(n8290), .op(n8513) );
  inv_1 U9958 ( .ip(n8513), .op(n10114) );
  mux2_1 U9959 ( .ip1(n8230), .ip2(n8229), .s(n10114), .op(n8303) );
  nor2_1 U9960 ( .ip1(n8232), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [15]), .op(
        n8234) );
  inv_1 U9961 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [12]), .op(n8231) );
  not_ab_or_c_or_d U9962 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [15]), .ip2(
        n8232), .ip3(\CORTEXM0DS_INST/u_logic/Zuh2z4 [14]), .ip4(n8231), .op(
        n8233) );
  or2_1 U9963 ( .ip1(n8234), .ip2(n8233), .op(n8235) );
  nand3_1 U9964 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [7]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [7]), .ip3(n8235), .op(n8236) );
  and3_1 U9965 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [6]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [6]), .ip3(n8236), .op(n10130) );
  mux2_1 U9966 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [15]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [13]), .s(n10130), .op(n8252) );
  nor2_1 U9967 ( .ip1(n8242), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [11]), .op(
        n8239) );
  not_ab_or_c_or_d U9968 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [11]), .ip2(
        n8242), .ip3(\CORTEXM0DS_INST/u_logic/Zuh2z4 [10]), .ip4(n8237), .op(
        n8238) );
  or2_1 U9969 ( .ip1(n8239), .ip2(n8238), .op(n8240) );
  nand3_1 U9970 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [5]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [5]), .ip3(n8240), .op(n8241) );
  and3_1 U9971 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [4]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [4]), .ip3(n8241), .op(n10120) );
  mux2_1 U9972 ( .ip1(n8243), .ip2(n8242), .s(n10120), .op(n8245) );
  inv_1 U9973 ( .ip(n8245), .op(n8251) );
  nor2_1 U9974 ( .ip1(n8252), .ip2(n8245), .op(n8247) );
  mux2_1 U9975 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [10]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [8]), .s(n10120), .op(n8274) );
  inv_1 U9976 ( .ip(n8274), .op(n8244) );
  mux2_1 U9977 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [14]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [12]), .s(n10130), .op(n8275) );
  not_ab_or_c_or_d U9978 ( .ip1(n8245), .ip2(n8252), .ip3(n8244), .ip4(n8275), 
        .op(n8246) );
  or2_1 U9979 ( .ip1(n8247), .ip2(n8246), .op(n8249) );
  nand2_1 U9980 ( .ip1(n8249), .ip2(n8248), .op(n10119) );
  and2_1 U9981 ( .ip1(n8250), .ip2(n10119), .op(n8511) );
  mux2_1 U9982 ( .ip1(n8252), .ip2(n8251), .s(n8511), .op(n8286) );
  nor2_1 U9983 ( .ip1(n11858), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [3]), .op(
        n8255) );
  inv_1 U9984 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [0]), .op(n8253) );
  not_ab_or_c_or_d U9985 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [3]), .ip2(
        n11858), .ip3(\CORTEXM0DS_INST/u_logic/Zuh2z4 [2]), .ip4(n8253), .op(
        n8254) );
  or2_1 U9986 ( .ip1(n8255), .ip2(n8254), .op(n8256) );
  nand3_1 U9987 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [1]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [1]), .ip3(n8256), .op(n8257) );
  and3_1 U9988 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [0]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [0]), .ip3(n8257), .op(n10123) );
  mux2_1 U9989 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [3]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [1]), .s(n10123), .op(n8271) );
  inv_1 U9990 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [5]), .op(n11833) );
  nor2_1 U9991 ( .ip1(n11833), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [7]), .op(
        n8260) );
  inv_1 U9992 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [4]), .op(n8258) );
  not_ab_or_c_or_d U9993 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [7]), .ip2(
        n11833), .ip3(\CORTEXM0DS_INST/u_logic/Zuh2z4 [6]), .ip4(n8258), .op(
        n8259) );
  or2_1 U9994 ( .ip1(n8260), .ip2(n8259), .op(n8261) );
  nand3_1 U9995 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [3]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [3]), .ip3(n8261), .op(n8262) );
  and3_1 U9996 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [2]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [2]), .ip3(n8262), .op(n10117) );
  mux2_1 U9997 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [7]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [5]), .s(n10117), .op(n8270) );
  inv_1 U9998 ( .ip(n8271), .op(n8264) );
  nor2_1 U9999 ( .ip1(n8270), .ip2(n8264), .op(n8266) );
  mux2_1 U10000 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [2]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [0]), .s(n10123), .op(n8273) );
  inv_1 U10001 ( .ip(n8273), .op(n8263) );
  mux2_1 U10002 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [6]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [4]), .s(n10117), .op(n8272) );
  not_ab_or_c_or_d U10003 ( .ip1(n8264), .ip2(n8270), .ip3(n8263), .ip4(n8272), 
        .op(n8265) );
  or2_1 U10004 ( .ip1(n8266), .ip2(n8265), .op(n8268) );
  nand2_1 U10005 ( .ip1(n8268), .ip2(n8267), .op(n10121) );
  nand2_1 U10006 ( .ip1(n8269), .ip2(n10121), .op(n10116) );
  mux2_1 U10007 ( .ip1(n8271), .ip2(n8270), .s(n10116), .op(n8285) );
  inv_1 U10008 ( .ip(n8285), .op(n8277) );
  nor2_1 U10009 ( .ip1(n8286), .ip2(n8277), .op(n8279) );
  mux2_1 U10010 ( .ip1(n8273), .ip2(n8272), .s(n10116), .op(n8295) );
  inv_1 U10011 ( .ip(n8295), .op(n8276) );
  mux2_1 U10012 ( .ip1(n8275), .ip2(n8274), .s(n8511), .op(n8296) );
  not_ab_or_c_or_d U10013 ( .ip1(n8277), .ip2(n8286), .ip3(n8276), .ip4(n8296), 
        .op(n8278) );
  or2_1 U10014 ( .ip1(n8279), .ip2(n8278), .op(n8280) );
  or2_1 U10015 ( .ip1(n8280), .ip2(n8281), .op(n8284) );
  or2_1 U10016 ( .ip1(n8282), .ip2(n8281), .op(n8283) );
  nand2_1 U10017 ( .ip1(n8284), .ip2(n8283), .op(n10122) );
  mux2_1 U10018 ( .ip1(n8286), .ip2(n8285), .s(n10122), .op(n8304) );
  inv_1 U10019 ( .ip(n8304), .op(n8298) );
  nor2_1 U10020 ( .ip1(n10114), .ip2(n8287), .op(n8301) );
  nor3_1 U10021 ( .ip1(n8303), .ip2(n8298), .ip3(n8301), .op(n8300) );
  nand2_1 U10022 ( .ip1(n10108), .ip2(n8288), .op(n8289) );
  nor2_1 U10023 ( .ip1(n8290), .ip2(n8289), .op(n8293) );
  nor2_1 U10024 ( .ip1(n10108), .ip2(n10114), .op(n8515) );
  and2_1 U10025 ( .ip1(n8291), .ip2(n8515), .op(n8292) );
  not_ab_or_c_or_d U10026 ( .ip1(n10114), .ip2(n8294), .ip3(n8293), .ip4(n8292), .op(n8305) );
  mux2_1 U10027 ( .ip1(n8296), .ip2(n8295), .s(n10122), .op(n8306) );
  nand2_1 U10028 ( .ip1(n8305), .ip2(n8306), .op(n8297) );
  not_ab_or_c_or_d U10029 ( .ip1(n8298), .ip2(n8303), .ip3(n8301), .ip4(n8297), 
        .op(n8299) );
  or2_1 U10030 ( .ip1(n8300), .ip2(n8299), .op(n8731) );
  nor2_1 U10031 ( .ip1(n8302), .ip2(n8731), .op(n10109) );
  nor2_1 U10032 ( .ip1(\CORTEXM0DS_INST/u_logic/Eqgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Krgvx4 ), .op(n8920) );
  nor2_1 U10033 ( .ip1(\CORTEXM0DS_INST/u_logic/Qsgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Wtgvx4 ), .op(n8331) );
  nand2_1 U10034 ( .ip1(n8302), .ip2(n8301), .op(n8312) );
  nor2_1 U10035 ( .ip1(\CORTEXM0DS_INST/u_logic/R3hvx4 ), .ip2(n8312), .op(
        n8327) );
  nand2_1 U10036 ( .ip1(n8331), .ip2(n8327), .op(n10104) );
  nand2_1 U10037 ( .ip1(n8920), .ip2(n10104), .op(n8811) );
  or2_1 U10038 ( .ip1(n10109), .ip2(n8811), .op(n8334) );
  inv_1 U10039 ( .ip(\CORTEXM0DS_INST/u_logic/Txh2z4 [1]), .op(n8308) );
  inv_1 U10040 ( .ip(n10109), .op(n10128) );
  mux2_1 U10041 ( .ip1(n8304), .ip2(n8303), .s(n10128), .op(n8314) );
  nor2_1 U10042 ( .ip1(n8308), .ip2(n8314), .op(n8310) );
  inv_1 U10043 ( .ip(\CORTEXM0DS_INST/u_logic/Txh2z4 [0]), .op(n8324) );
  inv_1 U10044 ( .ip(n8305), .op(n8307) );
  mux2_1 U10045 ( .ip1(n8307), .ip2(n8306), .s(n10109), .op(n8323) );
  not_ab_or_c_or_d U10046 ( .ip1(n8314), .ip2(n8308), .ip3(n8324), .ip4(n8323), 
        .op(n8309) );
  or2_1 U10047 ( .ip1(n8310), .ip2(n8309), .op(n8311) );
  inv_1 U10048 ( .ip(\CORTEXM0DS_INST/u_logic/R3hvx4 ), .op(n11730) );
  or2_1 U10049 ( .ip1(n8311), .ip2(n11730), .op(n8313) );
  nand2_1 U10050 ( .ip1(n8313), .ip2(n8312), .op(n8332) );
  mux2_1 U10051 ( .ip1(n8314), .ip2(\CORTEXM0DS_INST/u_logic/Txh2z4 [1]), .s(
        n8332), .op(n8931) );
  inv_1 U10052 ( .ip(\CORTEXM0DS_INST/u_logic/Wtgvx4 ), .op(n11885) );
  or2_1 U10053 ( .ip1(\CORTEXM0DS_INST/u_logic/Qsgvx4 ), .ip2(n11885), .op(
        n8321) );
  inv_1 U10054 ( .ip(\CORTEXM0DS_INST/u_logic/Uth2z4 [1]), .op(n8316) );
  nor2_1 U10055 ( .ip1(n8316), .ip2(\CORTEXM0DS_INST/u_logic/Psh2z4 [1]), .op(
        n8318) );
  not_ab_or_c_or_d U10056 ( .ip1(\CORTEXM0DS_INST/u_logic/Psh2z4 [1]), .ip2(
        n8316), .ip3(\CORTEXM0DS_INST/u_logic/Psh2z4 [0]), .ip4(n8315), .op(
        n8317) );
  or2_1 U10057 ( .ip1(n8318), .ip2(n8317), .op(n8319) );
  or2_1 U10058 ( .ip1(n8319), .ip2(n11885), .op(n8320) );
  nand2_1 U10059 ( .ip1(n8321), .ip2(n8320), .op(n10103) );
  mux2_1 U10060 ( .ip1(\CORTEXM0DS_INST/u_logic/Psh2z4 [1]), .ip2(
        \CORTEXM0DS_INST/u_logic/Uth2z4 [1]), .s(n10103), .op(n8322) );
  inv_1 U10061 ( .ip(n8322), .op(n8932) );
  nor3_1 U10062 ( .ip1(n8931), .ip2(n8932), .ip3(n8327), .op(n8329) );
  inv_1 U10063 ( .ip(n8323), .op(n8325) );
  mux2_1 U10064 ( .ip1(n8325), .ip2(n8324), .s(n8332), .op(n8927) );
  mux2_1 U10065 ( .ip1(\CORTEXM0DS_INST/u_logic/Psh2z4 [0]), .ip2(
        \CORTEXM0DS_INST/u_logic/Uth2z4 [0]), .s(n10103), .op(n8930) );
  nand2_1 U10066 ( .ip1(n8927), .ip2(n8930), .op(n8326) );
  not_ab_or_c_or_d U10067 ( .ip1(n8932), .ip2(n8931), .ip3(n8327), .ip4(n8326), 
        .op(n8328) );
  nor2_1 U10068 ( .ip1(n8329), .ip2(n8328), .op(n8738) );
  inv_1 U10069 ( .ip(n8738), .op(n8330) );
  nor2_1 U10070 ( .ip1(n8331), .ip2(n8330), .op(n10138) );
  nor2_1 U10071 ( .ip1(n8332), .ip2(n10138), .op(n8735) );
  or2_1 U10072 ( .ip1(n8735), .ip2(n8811), .op(n8333) );
  nand2_1 U10073 ( .ip1(n8334), .ip2(n8333), .op(n12471) );
  nand2_1 U10074 ( .ip1(\CORTEXM0DS_INST/u_logic/N6hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Xahvx4 ), .op(n9921) );
  nor3_1 U10075 ( .ip1(\CORTEXM0DS_INST/u_logic/L9hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/B5hvx4 ), .ip3(n9146), .op(n9134) );
  nand2_1 U10076 ( .ip1(n8714), .ip2(n9134), .op(n8474) );
  nor2_1 U10077 ( .ip1(n9921), .ip2(n8474), .op(n10246) );
  inv_1 U10078 ( .ip(n9196), .op(n8335) );
  mux2_1 U10079 ( .ip1(n8335), .ip2(n9168), .s(n10256), .op(n9669) );
  nor2_1 U10080 ( .ip1(n9669), .ip2(n11660), .op(n8347) );
  inv_1 U10081 ( .ip(n11899), .op(n11870) );
  nor3_1 U10082 ( .ip1(n11901), .ip2(n8337), .ip3(n9921), .op(n11842) );
  inv_1 U10083 ( .ip(n11842), .op(n11856) );
  nor2_1 U10084 ( .ip1(n8336), .ip2(n11856), .op(n8344) );
  nand2_1 U10085 ( .ip1(n8746), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [15]), 
        .op(n8342) );
  nand4_1 U10086 ( .ip1(\CORTEXM0DS_INST/u_logic/N6hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Z7hvx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/B5hvx4 ), .ip4(n11901), .op(n8338) );
  nor2_1 U10087 ( .ip1(n11898), .ip2(n8338), .op(n11864) );
  nand2_1 U10088 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [11]), .ip2(n11864), 
        .op(n8341) );
  nor3_1 U10089 ( .ip1(n11901), .ip2(n8337), .ip3(n8659), .op(n11863) );
  nand2_1 U10090 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [19]), .ip2(n11863), 
        .op(n8340) );
  nor2_1 U10091 ( .ip1(\CORTEXM0DS_INST/u_logic/Xahvx4 ), .ip2(n8338), .op(
        n11841) );
  nand2_1 U10092 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [3]), .ip2(n11841), 
        .op(n8339) );
  nand4_1 U10093 ( .ip1(n8342), .ip2(n8341), .ip3(n8340), .ip4(n8339), .op(
        n8343) );
  not_ab_or_c_or_d U10094 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [15]), .ip2(
        n11870), .ip3(n8344), .ip4(n8343), .op(n8345) );
  nor2_1 U10095 ( .ip1(n8345), .ip2(n11871), .op(n8346) );
  not_ab_or_c_or_d U10096 ( .ip1(n12471), .ip2(n10246), .ip3(n8347), .ip4(
        n8346), .op(n8348) );
  nand3_1 U10097 ( .ip1(n8349), .ip2(n8348), .ip3(n3045), .op(n10451) );
  nand2_1 U10098 ( .ip1(n8350), .ip2(n10451), .op(n8353) );
  or2_1 U10099 ( .ip1(n8614), .ip2(n8351), .op(n8352) );
  nand2_1 U10100 ( .ip1(n8353), .ip2(n8352), .op(n8354) );
  nor4_1 U10101 ( .ip1(n9247), .ip2(n8356), .ip3(n8355), .ip4(n8354), .op(
        n8599) );
  not_ab_or_c_or_d U10102 ( .ip1(n8601), .ip2(n9207), .ip3(n8357), .ip4(n8599), 
        .op(n10369) );
  inv_1 U10103 ( .ip(n8595), .op(n9686) );
  nand3_1 U10104 ( .ip1(n9686), .ip2(n8601), .ip3(n8526), .op(n8810) );
  inv_1 U10105 ( .ip(n8810), .op(n8361) );
  nand3_1 U10106 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n11051), .ip3(
        n8613), .op(n8784) );
  nand2_1 U10107 ( .ip1(n11065), .ip2(n8358), .op(n8359) );
  or2_1 U10108 ( .ip1(n8359), .ip2(n8592), .op(n8360) );
  nand2_1 U10109 ( .ip1(n8784), .ip2(n8360), .op(n8615) );
  nor2_1 U10110 ( .ip1(n8361), .ip2(n8615), .op(n10350) );
  inv_1 U10111 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [3]), .op(n11708) );
  nor2_1 U10112 ( .ip1(n11708), .ip2(n11830), .op(n8375) );
  nand2_1 U10113 ( .ip1(n9183), .ip2(n8699), .op(n8365) );
  nand2_1 U10114 ( .ip1(n9181), .ip2(n8698), .op(n8364) );
  nand2_1 U10115 ( .ip1(n9179), .ip2(n9155), .op(n8363) );
  inv_1 U10116 ( .ip(n9157), .op(n8691) );
  nand2_1 U10117 ( .ip1(n9185), .ip2(n8691), .op(n8362) );
  nand4_1 U10118 ( .ip1(n8365), .ip2(n8364), .ip3(n8363), .ip4(n8362), .op(
        n9223) );
  nor2_1 U10119 ( .ip1(n10256), .ip2(n9223), .op(n9215) );
  nand2_1 U10120 ( .ip1(n9181), .ip2(n8461), .op(n8369) );
  nand2_1 U10121 ( .ip1(n9183), .ip2(n8643), .op(n8368) );
  nand2_1 U10122 ( .ip1(n9179), .ip2(n8462), .op(n8367) );
  nand2_1 U10123 ( .ip1(n9185), .ip2(n8790), .op(n8366) );
  nand4_1 U10124 ( .ip1(n8369), .ip2(n8368), .ip3(n8367), .ip4(n8366), .op(
        n9242) );
  nor2_1 U10125 ( .ip1(n8781), .ip2(n9242), .op(n9217) );
  nor3_1 U10126 ( .ip1(n9215), .ip2(n9217), .ip3(n11660), .op(n8371) );
  and2_1 U10127 ( .ip1(n10271), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [3]), 
        .op(n8370) );
  not_ab_or_c_or_d U10128 ( .ip1(n10270), .ip2(
        \CORTEXM0DS_INST/u_logic/Czh2z4 [3]), .ip3(n8371), .ip4(n8370), .op(
        n8373) );
  inv_1 U10129 ( .ip(n8474), .op(n8372) );
  nand2_1 U10130 ( .ip1(n8651), .ip2(n8372), .op(n8446) );
  nand3_1 U10131 ( .ip1(n4203), .ip2(n8373), .ip3(n8446), .op(n8374) );
  not_ab_or_c_or_d U10132 ( .ip1(n11829), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [3]), .ip3(n8375), .ip4(n8374), .op(
        n10435) );
  nor2_1 U10133 ( .ip1(n10350), .ip2(n10435), .op(n8376) );
  not_ab_or_c_or_d U10134 ( .ip1(n10370), .ip2(n10438), .ip3(n10369), .ip4(
        n8376), .op(n8398) );
  nor2_1 U10135 ( .ip1(n9670), .ip2(n8594), .op(n8527) );
  inv_1 U10136 ( .ip(n9659), .op(n8378) );
  inv_1 U10137 ( .ip(n8377), .op(n8590) );
  not_ab_or_c_or_d U10138 ( .ip1(n8378), .ip2(n8590), .ip3(n8614), .ip4(n8592), 
        .op(n8379) );
  or2_1 U10139 ( .ip1(n8527), .ip2(n8379), .op(n10364) );
  nor2_1 U10140 ( .ip1(\CORTEXM0DS_INST/u_logic/Z7hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/B5hvx4 ), .op(n8380) );
  nand4_1 U10141 ( .ip1(\CORTEXM0DS_INST/u_logic/N6hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Xahvx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/L9hvx4 ), .ip4(n8380), .op(n12055) );
  or2_1 U10142 ( .ip1(n11871), .ip2(n12055), .op(n10259) );
  and2_1 U10143 ( .ip1(n9256), .ip2(n11853), .op(n10248) );
  nand2_1 U10144 ( .ip1(n8526), .ip2(n9704), .op(n8486) );
  nor2_1 U10145 ( .ip1(n8424), .ip2(n8486), .op(n9229) );
  nor2_1 U10146 ( .ip1(n10256), .ip2(n8486), .op(n8383) );
  nand2_1 U10147 ( .ip1(n10256), .ip2(n8486), .op(n8381) );
  nand2_1 U10148 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n8381), .op(
        n8382) );
  nor2_1 U10149 ( .ip1(n8383), .ip2(n8382), .op(n9230) );
  mux2_1 U10150 ( .ip1(n9229), .ip2(n9230), .s(n9243), .op(n8394) );
  nand2_1 U10151 ( .ip1(n10248), .ip2(n8394), .op(n8396) );
  nor2_1 U10152 ( .ip1(n8797), .ip2(n9158), .op(n8388) );
  inv_1 U10153 ( .ip(n8638), .op(n8796) );
  nor2_1 U10154 ( .ip1(n8796), .ip2(n9156), .op(n8387) );
  nor2_1 U10155 ( .ip1(n9349), .ip2(n9243), .op(n8386) );
  inv_1 U10156 ( .ip(n8384), .op(n8798) );
  nor2_1 U10157 ( .ip1(n8798), .ip2(n9160), .op(n8385) );
  nor4_1 U10158 ( .ip1(n8388), .ip2(n8387), .ip3(n8386), .ip4(n8385), .op(
        n9240) );
  nand2_1 U10159 ( .ip1(n9179), .ip2(n8774), .op(n8392) );
  inv_1 U10160 ( .ip(n8673), .op(n8775) );
  nand2_1 U10161 ( .ip1(n9183), .ip2(n8775), .op(n8391) );
  nand2_1 U10162 ( .ip1(n9181), .ip2(n8768), .op(n8390) );
  inv_1 U10163 ( .ip(n9287), .op(n8773) );
  nand2_1 U10164 ( .ip1(n9185), .ip2(n8773), .op(n8389) );
  nand4_1 U10165 ( .ip1(n8392), .ip2(n8391), .ip3(n8390), .ip4(n8389), .op(
        n9190) );
  nor2_1 U10166 ( .ip1(n9190), .ip2(n8781), .op(n8393) );
  not_ab_or_c_or_d U10167 ( .ip1(n9240), .ip2(n8781), .ip3(n8394), .ip4(n8393), 
        .op(n9237) );
  nand2_1 U10168 ( .ip1(n9237), .ip2(n11853), .op(n8395) );
  nand4_1 U10169 ( .ip1(n4175), .ip2(n10259), .ip3(n8396), .ip4(n8395), .op(
        n10440) );
  nand2_1 U10170 ( .ip1(n10364), .ip2(n10440), .op(n8397) );
  nand3_1 U10171 ( .ip1(n8399), .ip2(n8398), .ip3(n8397), .op(n11310) );
  nand2_1 U10172 ( .ip1(n10475), .ip2(n11310), .op(n8403) );
  xor2_1 U10173 ( .ip1(n8401), .ip2(n8400), .op(n12188) );
  inv_1 U10174 ( .ip(n12188), .op(n11312) );
  nand2_1 U10175 ( .ip1(n11312), .ip2(n10916), .op(n8402) );
  nand4_1 U10176 ( .ip1(n8404), .ip2(n10917), .ip3(n8403), .ip4(n8402), .op(
        \CORTEXM0DS_INST/u_logic/Uehvx4 ) );
  xor2_1 U10177 ( .ip1(n8406), .ip2(n8405), .op(n12169) );
  nand2_1 U10178 ( .ip1(n12169), .ip2(n10916), .op(n8483) );
  nand2_1 U10179 ( .ip1(n10344), .ip2(n12113), .op(n8407) );
  mux2_1 U10180 ( .ip1(n10344), .ip2(n8407), .s(\CORTEXM0DS_INST/vis_pc [8]), 
        .op(n8482) );
  nor2_1 U10181 ( .ip1(n10256), .ip2(n11660), .op(n11645) );
  nor2_1 U10182 ( .ip1(n8821), .ip2(n9158), .op(n8412) );
  nor2_1 U10183 ( .ip1(n8408), .ip2(n9243), .op(n8411) );
  inv_1 U10184 ( .ip(n8824), .op(n8724) );
  nor2_1 U10185 ( .ip1(n8724), .ip2(n9156), .op(n8410) );
  inv_1 U10186 ( .ip(n8815), .op(n8725) );
  nor2_1 U10187 ( .ip1(n8725), .ip2(n9160), .op(n8409) );
  nor4_1 U10188 ( .ip1(n8412), .ip2(n8411), .ip3(n8410), .ip4(n8409), .op(
        n9166) );
  inv_1 U10189 ( .ip(n10285), .op(n8467) );
  nor2_1 U10190 ( .ip1(n9166), .ip2(n8467), .op(n8417) );
  or2_1 U10191 ( .ip1(n11645), .ip2(n8417), .op(n8419) );
  nand2_1 U10192 ( .ip1(n9183), .ip2(n9180), .op(n8416) );
  nand2_1 U10193 ( .ip1(n9181), .ip2(n8814), .op(n8415) );
  nand2_1 U10194 ( .ip1(n9179), .ip2(n8816), .op(n8414) );
  nand2_1 U10195 ( .ip1(n9185), .ip2(n9178), .op(n8413) );
  nand4_1 U10196 ( .ip1(n8416), .ip2(n8415), .ip3(n8414), .ip4(n8413), .op(
        n9191) );
  or2_1 U10197 ( .ip1(n9191), .ip2(n8417), .op(n8418) );
  nand2_1 U10198 ( .ip1(n8419), .ip2(n8418), .op(n8422) );
  nand2_1 U10199 ( .ip1(n10270), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [17]), 
        .op(n8421) );
  nand2_1 U10200 ( .ip1(n10271), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [17]), 
        .op(n8420) );
  nand4_1 U10201 ( .ip1(n3197), .ip2(n8422), .ip3(n8421), .ip4(n8420), .op(
        n10911) );
  nand2_1 U10202 ( .ip1(n10911), .ip2(n10370), .op(n8480) );
  nand2_1 U10203 ( .ip1(n8781), .ip2(n9185), .op(n8425) );
  nor2_1 U10204 ( .ip1(n8486), .ip2(n8425), .op(n8423) );
  not_ab_or_c_or_d U10205 ( .ip1(n8486), .ip2(n8425), .ip3(n8424), .ip4(n8423), 
        .op(n8436) );
  nand2_1 U10206 ( .ip1(n8436), .ip2(n10248), .op(n8438) );
  inv_1 U10207 ( .ip(n8768), .op(n8670) );
  nor2_1 U10208 ( .ip1(n8670), .ip2(n9156), .op(n8430) );
  nor2_1 U10209 ( .ip1(n8426), .ip2(n9243), .op(n8429) );
  nor2_1 U10210 ( .ip1(n8672), .ip2(n9158), .op(n8428) );
  nor2_1 U10211 ( .ip1(n8671), .ip2(n9160), .op(n8427) );
  nor4_1 U10212 ( .ip1(n8430), .ip2(n8429), .ip3(n8428), .ip4(n8427), .op(
        n9192) );
  nand2_1 U10213 ( .ip1(n9181), .ip2(n8775), .op(n8434) );
  nand2_1 U10214 ( .ip1(n9183), .ip2(n8776), .op(n8433) );
  nand2_1 U10215 ( .ip1(n9179), .ip2(n8773), .op(n8432) );
  nand2_1 U10216 ( .ip1(n9185), .ip2(n8637), .op(n8431) );
  nand4_1 U10217 ( .ip1(n8434), .ip2(n8433), .ip3(n8432), .ip4(n8431), .op(
        n8488) );
  nor2_1 U10218 ( .ip1(n8488), .ip2(n10256), .op(n8435) );
  not_ab_or_c_or_d U10219 ( .ip1(n10256), .ip2(n9192), .ip3(n8436), .ip4(n8435), .op(n9250) );
  nand2_1 U10220 ( .ip1(n9250), .ip2(n11853), .op(n8437) );
  nand4_1 U10221 ( .ip1(n3212), .ip2(n10259), .ip3(n8438), .ip4(n8437), .op(
        n10905) );
  inv_1 U10222 ( .ip(n10362), .op(n10351) );
  inv_1 U10223 ( .ip(n9147), .op(n8719) );
  nand2_1 U10224 ( .ip1(n9179), .ip2(n8719), .op(n8442) );
  nand2_1 U10225 ( .ip1(n9181), .ip2(n8693), .op(n8441) );
  nand2_1 U10226 ( .ip1(n9183), .ip2(n8718), .op(n8440) );
  nand2_1 U10227 ( .ip1(n9185), .ip2(n8822), .op(n8439) );
  nand4_1 U10228 ( .ip1(n8442), .ip2(n8441), .ip3(n8440), .ip4(n8439), .op(
        n9172) );
  nand2_1 U10229 ( .ip1(n10271), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [9]), 
        .op(n8445) );
  nand2_1 U10230 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [9]), .ip2(n10272), 
        .op(n8444) );
  nand2_1 U10231 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [9]), .ip2(n11829), 
        .op(n8443) );
  nand4_1 U10232 ( .ip1(n8446), .ip2(n8445), .ip3(n8444), .ip4(n8443), .op(
        n8455) );
  nor2_1 U10233 ( .ip1(n8659), .ip2(n8474), .op(n4241) );
  inv_1 U10234 ( .ip(n4241), .op(n8453) );
  nand2_1 U10235 ( .ip1(n9179), .ip2(n8691), .op(n8450) );
  nand2_1 U10236 ( .ip1(n9183), .ip2(n8692), .op(n8449) );
  nand2_1 U10237 ( .ip1(n9181), .ip2(n8699), .op(n8448) );
  nand2_1 U10238 ( .ip1(n9185), .ip2(n8690), .op(n8447) );
  nand4_1 U10239 ( .ip1(n8450), .ip2(n8449), .ip3(n8448), .ip4(n8447), .op(
        n9170) );
  nand2_1 U10240 ( .ip1(n10285), .ip2(n9170), .op(n8452) );
  nand2_1 U10241 ( .ip1(n10270), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [9]), 
        .op(n8451) );
  nand4_1 U10242 ( .ip1(n3166), .ip2(n8453), .ip3(n8452), .ip4(n8451), .op(
        n8454) );
  not_ab_or_c_or_d U10243 ( .ip1(n11645), .ip2(n9172), .ip3(n8455), .ip4(n8454), .op(n10903) );
  nor2_1 U10244 ( .ip1(n10351), .ip2(n10903), .op(n8456) );
  not_ab_or_c_or_d U10245 ( .ip1(n10364), .ip2(n10905), .ip3(n10369), .ip4(
        n8456), .op(n8479) );
  inv_1 U10246 ( .ip(n10350), .op(n10361) );
  nand2_1 U10247 ( .ip1(n9179), .ip2(n8790), .op(n8460) );
  nand2_1 U10248 ( .ip1(n9181), .ip2(n8643), .op(n8459) );
  nand2_1 U10249 ( .ip1(n9183), .ip2(n8698), .op(n8458) );
  nand2_1 U10250 ( .ip1(n9185), .ip2(n9155), .op(n8457) );
  nand4_1 U10251 ( .ip1(n8460), .ip2(n8459), .ip3(n8458), .ip4(n8457), .op(
        n9220) );
  nor2_1 U10252 ( .ip1(n8798), .ip2(n9158), .op(n8466) );
  inv_1 U10253 ( .ip(n8461), .op(n8799) );
  nor2_1 U10254 ( .ip1(n8799), .ip2(n9156), .op(n8465) );
  nor2_1 U10255 ( .ip1(n8796), .ip2(n9243), .op(n8464) );
  inv_1 U10256 ( .ip(n8462), .op(n8789) );
  nor2_1 U10257 ( .ip1(n8789), .ip2(n9160), .op(n8463) );
  nor4_1 U10258 ( .ip1(n8466), .ip2(n8465), .ip3(n8464), .ip4(n8463), .op(
        n9218) );
  nor2_1 U10259 ( .ip1(n9218), .ip2(n8467), .op(n8473) );
  nand2_1 U10260 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [1]), .ip2(n11829), 
        .op(n8471) );
  nand3_1 U10261 ( .ip1(n8714), .ip2(n11902), .ip3(n11903), .op(n10281) );
  inv_1 U10262 ( .ip(n10281), .op(n8829) );
  nand2_1 U10263 ( .ip1(n8829), .ip2(\CORTEXM0DS_INST/u_logic/S0hvx4 ), .op(
        n8470) );
  nand2_1 U10264 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [1]), .ip2(n10272), 
        .op(n8469) );
  nand2_1 U10265 ( .ip1(n10271), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [1]), 
        .op(n8468) );
  nand4_1 U10266 ( .ip1(n8471), .ip2(n8470), .ip3(n8469), .ip4(n8468), .op(
        n8472) );
  not_ab_or_c_or_d U10267 ( .ip1(n11645), .ip2(n9220), .ip3(n8473), .ip4(n8472), .op(n8477) );
  nand2_1 U10268 ( .ip1(n10270), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [1]), 
        .op(n8476) );
  nor2_1 U10269 ( .ip1(n12689), .ip2(n8474), .op(n10278) );
  nand2_1 U10270 ( .ip1(\CORTEXM0DS_INST/u_logic/Eg8vx4 ), .ip2(n10278), .op(
        n8475) );
  nand4_1 U10271 ( .ip1(n3187), .ip2(n8477), .ip3(n8476), .ip4(n8475), .op(
        n10904) );
  nand2_1 U10272 ( .ip1(n10361), .ip2(n10904), .op(n8478) );
  nand3_1 U10273 ( .ip1(n8480), .ip2(n8479), .ip3(n8478), .op(n11761) );
  nand2_1 U10274 ( .ip1(n10475), .ip2(n11761), .op(n8481) );
  nand4_1 U10275 ( .ip1(n10917), .ip2(n8483), .ip3(n8482), .ip4(n8481), .op(
        \CORTEXM0DS_INST/u_logic/Bfhvx4 ) );
  nand2_1 U10276 ( .ip1(n8485), .ip2(n8484), .op(n10597) );
  inv_1 U10277 ( .ip(n9230), .op(n9245) );
  nand2_1 U10278 ( .ip1(n8486), .ip2(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .op(
        n9244) );
  mux2_1 U10279 ( .ip1(n9245), .ip2(n9244), .s(n9185), .op(n8487) );
  inv_1 U10280 ( .ip(n8487), .op(n8490) );
  nand2_1 U10281 ( .ip1(n10248), .ip2(n8490), .op(n8492) );
  nor2_1 U10282 ( .ip1(n8488), .ip2(n8781), .op(n8489) );
  not_ab_or_c_or_d U10283 ( .ip1(n9218), .ip2(n8781), .ip3(n8490), .ip4(n8489), 
        .op(n9238) );
  nand2_1 U10284 ( .ip1(n9238), .ip2(n11853), .op(n8491) );
  nand4_1 U10285 ( .ip1(n3068), .ip2(n10259), .ip3(n8492), .ip4(n8491), .op(
        n10374) );
  inv_1 U10286 ( .ip(n9701), .op(n8493) );
  inv_1 U10287 ( .ip(n9251), .op(n9208) );
  nand2_1 U10288 ( .ip1(n9208), .ip2(n8526), .op(n9695) );
  nand2_1 U10289 ( .ip1(n8493), .ip2(n9695), .op(n9697) );
  or2_1 U10290 ( .ip1(n8494), .ip2(n12117), .op(n8497) );
  or2_1 U10291 ( .ip1(n8495), .ip2(n12117), .op(n8496) );
  nand2_1 U10292 ( .ip1(n8497), .ip2(n8496), .op(n8498) );
  nor2_1 U10293 ( .ip1(n8498), .ip2(n8604), .op(n8765) );
  not_ab_or_c_or_d U10294 ( .ip1(n9697), .ip2(n8592), .ip3(n8765), .ip4(n8599), 
        .op(n10595) );
  nand2_1 U10295 ( .ip1(n8810), .ip2(n8784), .op(n10593) );
  nand2_1 U10296 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [21]), .ip2(n10270), 
        .op(n8502) );
  inv_1 U10297 ( .ip(n11645), .op(n10087) );
  nor2_1 U10298 ( .ip1(n9192), .ip2(n10087), .op(n8500) );
  inv_1 U10299 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [21]), .op(n12031) );
  nor2_1 U10300 ( .ip1(n11875), .ip2(n12031), .op(n8499) );
  not_ab_or_c_or_d U10301 ( .ip1(n10285), .ip2(n9191), .ip3(n8500), .ip4(n8499), .op(n8501) );
  nand3_1 U10302 ( .ip1(n8502), .ip2(n8501), .ip3(n3102), .op(n10379) );
  or2_1 U10303 ( .ip1(n8782), .ip2(n8596), .op(n8504) );
  or2_1 U10304 ( .ip1(n8526), .ip2(n8596), .op(n8503) );
  nand2_1 U10305 ( .ip1(n8504), .ip2(n8503), .op(n10589) );
  inv_1 U10306 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [5]), .op(n11739) );
  nor2_1 U10307 ( .ip1(n11739), .ip2(n11830), .op(n8508) );
  nand2_1 U10308 ( .ip1(n10285), .ip2(n9220), .op(n8506) );
  nand2_1 U10309 ( .ip1(n10270), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [5]), 
        .op(n8505) );
  nand3_1 U10310 ( .ip1(n8506), .ip2(n3085), .ip3(n8505), .op(n8507) );
  not_ab_or_c_or_d U10311 ( .ip1(n11645), .ip2(n9170), .ip3(n8508), .ip4(n8507), .op(n10187) );
  nor2_1 U10312 ( .ip1(n10589), .ip2(n10187), .op(n8529) );
  nor2_1 U10313 ( .ip1(n9166), .ip2(n10087), .op(n8525) );
  inv_1 U10314 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [13]), .op(n11718) );
  nor2_1 U10315 ( .ip1(n11718), .ip2(n11830), .op(n8510) );
  inv_1 U10316 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [13]), .op(n11994) );
  nor2_1 U10317 ( .ip1(n11875), .ip2(n11994), .op(n8509) );
  not_ab_or_c_or_d U10318 ( .ip1(n10270), .ip2(
        \CORTEXM0DS_INST/u_logic/Czh2z4 [13]), .ip3(n8510), .ip4(n8509), .op(
        n8523) );
  and2_1 U10319 ( .ip1(n10116), .ip2(n10122), .op(n8512) );
  nor2_1 U10320 ( .ip1(n8511), .ip2(n10122), .op(n10129) );
  nor2_1 U10321 ( .ip1(n8512), .ip2(n10129), .op(n8517) );
  nor2_1 U10322 ( .ip1(n8514), .ip2(n8513), .op(n10111) );
  nor2_1 U10323 ( .ip1(n8515), .ip2(n10111), .op(n8516) );
  mux2_1 U10324 ( .ip1(n8517), .ip2(n8516), .s(n10128), .op(n8518) );
  nand2_1 U10325 ( .ip1(n8518), .ip2(n8735), .op(n8519) );
  nand2_1 U10326 ( .ip1(n10104), .ip2(n8519), .op(n8520) );
  nand2_1 U10327 ( .ip1(n8920), .ip2(n8520), .op(n12458) );
  nand2_1 U10328 ( .ip1(n10246), .ip2(n12458), .op(n8522) );
  nand2_1 U10329 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [13]), .ip2(n11829), 
        .op(n8521) );
  nand4_1 U10330 ( .ip1(n2974), .ip2(n8523), .ip3(n8522), .ip4(n8521), .op(
        n8524) );
  not_ab_or_c_or_d U10331 ( .ip1(n10285), .ip2(n9172), .ip3(n8525), .ip4(n8524), .op(n10375) );
  nand2_1 U10332 ( .ip1(n8527), .ip2(n8526), .op(n10586) );
  nor2_1 U10333 ( .ip1(n10375), .ip2(n10586), .op(n8528) );
  ab_or_c_or_d U10334 ( .ip1(n10593), .ip2(n10379), .ip3(n8529), .ip4(n8528), 
        .op(n8530) );
  not_ab_or_c_or_d U10335 ( .ip1(n10597), .ip2(n10374), .ip3(n10595), .ip4(
        n8530), .op(n11821) );
  or2_1 U10336 ( .ip1(n11821), .ip2(n10912), .op(n8580) );
  inv_1 U10337 ( .ip(\CORTEXM0DS_INST/vis_pc [22]), .op(n12144) );
  inv_1 U10338 ( .ip(\CORTEXM0DS_INST/vis_pc [15]), .op(n12211) );
  nor3_1 U10339 ( .ip1(n11005), .ip2(n12211), .ip3(n12220), .op(n10081) );
  nand4_1 U10340 ( .ip1(\CORTEXM0DS_INST/vis_pc [17]), .ip2(
        \CORTEXM0DS_INST/vis_pc [18]), .ip3(\CORTEXM0DS_INST/vis_pc [19]), 
        .ip4(n10081), .op(n8894) );
  nor3_1 U10341 ( .ip1(n8531), .ip2(n12144), .ip3(n8894), .op(n10168) );
  nand4_1 U10342 ( .ip1(\CORTEXM0DS_INST/vis_pc [23]), .ip2(
        \CORTEXM0DS_INST/vis_pc [24]), .ip3(\CORTEXM0DS_INST/vis_pc [25]), 
        .ip4(n10168), .op(n10456) );
  nand2_1 U10343 ( .ip1(n8533), .ip2(n8532), .op(n10455) );
  nor2_1 U10344 ( .ip1(n5814), .ip2(n10455), .op(n10327) );
  inv_1 U10345 ( .ip(n10327), .op(n10164) );
  nor2_1 U10346 ( .ip1(n10456), .ip2(n10164), .op(n10290) );
  nand2_1 U10347 ( .ip1(\CORTEXM0DS_INST/vis_pc [26]), .ip2(n10290), .op(
        n10240) );
  nor2_1 U10348 ( .ip1(n10231), .ip2(n10240), .op(n10230) );
  or2_1 U10349 ( .ip1(\CORTEXM0DS_INST/vis_pc [28]), .ip2(n10230), .op(n8534)
         );
  nand2_1 U10350 ( .ip1(\CORTEXM0DS_INST/vis_pc [28]), .ip2(n10230), .op(
        n10603) );
  nand3_1 U10351 ( .ip1(n12113), .ip2(n8534), .ip3(n10603), .op(n8579) );
  inv_1 U10352 ( .ip(n8535), .op(n8536) );
  nor2_1 U10353 ( .ip1(n8537), .ip2(n8536), .op(n9303) );
  or2_1 U10354 ( .ip1(n8539), .ip2(n8538), .op(n8540) );
  nand2_1 U10355 ( .ip1(n8541), .ip2(n8540), .op(n9263) );
  nand2_1 U10356 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [29]), .op(n8544) );
  nand2_1 U10357 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [29]), .op(n8543) );
  nand2_1 U10358 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [29]), .op(n8542) );
  nand3_1 U10359 ( .ip1(n8544), .ip2(n8543), .ip3(n8542), .op(n8561) );
  and2_1 U10360 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [27]), .op(n8546)
         );
  inv_1 U10361 ( .ip(\CORTEXM0DS_INST/u_logic/H3evx4 ), .op(n9288) );
  nor2_1 U10362 ( .ip1(n9279), .ip2(n9288), .op(n8545) );
  not_ab_or_c_or_d U10363 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [29]), 
        .ip3(n8546), .ip4(n8545), .op(n8559) );
  nand2_1 U10364 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [29]), .op(n8550) );
  nand2_1 U10365 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [29]), .op(n8549) );
  nand2_1 U10366 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [29]), .op(n8548) );
  nand2_1 U10367 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [29]), .op(n8547) );
  nand2_1 U10368 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [29]), .op(n8553) );
  nand2_1 U10369 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [29]), .op(n8552) );
  nand2_1 U10370 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [29]), .op(n8551) );
  nand3_1 U10371 ( .ip1(n8553), .ip2(n8552), .ip3(n8551), .op(n8554) );
  not_ab_or_c_or_d U10372 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [29]), 
        .ip3(n8555), .ip4(n8554), .op(n8558) );
  nand2_1 U10373 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [27]), .op(n8557) );
  nand2_1 U10374 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [29]), .op(n8556) );
  not_ab_or_c_or_d U10375 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [29]), 
        .ip3(n8561), .ip4(n8560), .op(n11819) );
  inv_1 U10376 ( .ip(n11819), .op(n11488) );
  mux2_1 U10377 ( .ip1(n8563), .ip2(n8562), .s(n11488), .op(n9525) );
  and2_1 U10378 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [29]), .ip2(n9354), .op(n8572)
         );
  nor2_1 U10379 ( .ip1(n12088), .ip2(n8564), .op(n8566) );
  nor2_1 U10380 ( .ip1(n8673), .ip2(n9348), .op(n8565) );
  not_ab_or_c_or_d U10381 ( .ip1(\CORTEXM0DS_INST/vis_msp [27]), .ip2(n9366), 
        .ip3(n8566), .ip4(n8565), .op(n8570) );
  nand2_1 U10382 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [29]), .ip2(n9355), .op(n8569) );
  nand2_1 U10383 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [29]), .ip2(n9364), .op(n8568) );
  nand2_1 U10384 ( .ip1(\CORTEXM0DS_INST/u_logic/H3evx4 ), .ip2(n9353), .op(
        n8567) );
  not_ab_or_c_or_d U10385 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [29]), .ip2(n9363), 
        .ip3(n8572), .ip4(n8571), .op(n8576) );
  nand2_1 U10386 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [29]), .ip2(n9347), .op(n8575) );
  nand2_1 U10387 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [29]), .ip2(n9365), .op(n8574) );
  nand2_1 U10388 ( .ip1(\CORTEXM0DS_INST/vis_psp [27]), .ip2(n9356), .op(n8573) );
  inv_1 U10389 ( .ip(n9524), .op(n10040) );
  nor2_1 U10390 ( .ip1(n9371), .ip2(n10040), .op(n8577) );
  xor2_1 U10391 ( .ip1(n9525), .ip2(n8577), .op(n9262) );
  xor2_1 U10392 ( .ip1(n9263), .ip2(n9262), .op(n9302) );
  xor2_1 U10393 ( .ip1(n9303), .ip2(n9302), .op(n10033) );
  nand2_1 U10394 ( .ip1(n10033), .ip2(n10916), .op(n8578) );
  nand4_1 U10395 ( .ip1(n10917), .ip2(n8580), .ip3(n8579), .ip4(n8578), .op(
        \CORTEXM0DS_INST/u_logic/Mhhvx4 ) );
  nand2_1 U10396 ( .ip1(\CORTEXM0DS_INST/vis_pc [0]), .ip2(n12359), .op(n8585)
         );
  nand2_1 U10397 ( .ip1(\CORTEXM0DS_INST/u_logic/Uzcvx4 ), .ip2(n2119), .op(
        n8584) );
  nand2_1 U10398 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [1]), .ip2(n12358), .op(
        n8583) );
  inv_1 U10399 ( .ip(n12355), .op(n2118) );
  nand3_1 U10400 ( .ip1(n2118), .ip2(n8581), .ip3(n11201), .op(n8582) );
  nand4_1 U10401 ( .ip1(n8585), .ip2(n8584), .ip3(n8583), .ip4(n8582), .op(
        n6077) );
  inv_1 U10402 ( .ip(n9415), .op(n11432) );
  nand2_1 U10403 ( .ip1(n11432), .ip2(n10916), .op(n8622) );
  nor2_1 U10404 ( .ip1(n5814), .ip2(n8586), .op(n10415) );
  inv_1 U10405 ( .ip(n10415), .op(n8634) );
  nand2_1 U10406 ( .ip1(n8634), .ip2(n8587), .op(n8588) );
  nand2_1 U10407 ( .ip1(\CORTEXM0DS_INST/vis_pc [2]), .ip2(n10415), .op(n10400) );
  nand3_1 U10408 ( .ip1(n8588), .ip2(n12113), .ip3(n10400), .op(n8621) );
  inv_1 U10409 ( .ip(n9670), .op(n9682) );
  nand3_1 U10410 ( .ip1(n9211), .ip2(n9682), .ip3(n8601), .op(n8603) );
  nand3_1 U10411 ( .ip1(n12609), .ip2(n12118), .ip3(n8593), .op(n8589) );
  ab_or_c_or_d U10412 ( .ip1(n8590), .ip2(n8589), .ip3(n8614), .ip4(n8592), 
        .op(n8591) );
  nand2_1 U10413 ( .ip1(n8603), .ip2(n8591), .op(n11037) );
  nand2_1 U10414 ( .ip1(n10438), .ip2(n11037), .op(n8619) );
  nor2_1 U10415 ( .ip1(n8614), .ip2(n8592), .op(n8598) );
  nor3_1 U10416 ( .ip1(n8593), .ip2(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Fjgvx4 ), .op(n8612) );
  nor2_1 U10417 ( .ip1(n8595), .ip2(n8594), .op(n8597) );
  not_ab_or_c_or_d U10418 ( .ip1(n8598), .ip2(n8612), .ip3(n8597), .ip4(n8596), 
        .op(n11039) );
  inv_1 U10419 ( .ip(n11039), .op(n10906) );
  inv_1 U10420 ( .ip(n8599), .op(n8763) );
  nand2_1 U10421 ( .ip1(n8601), .ip2(n8600), .op(n8602) );
  nand4_1 U10422 ( .ip1(n8763), .ip2(n8604), .ip3(n8603), .ip4(n8602), .op(
        n11045) );
  inv_1 U10423 ( .ip(n11045), .op(n10376) );
  or2_1 U10424 ( .ip1(n8606), .ip2(n8605), .op(n8607) );
  nand3_1 U10425 ( .ip1(n10944), .ip2(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip3(
        n8607), .op(n8608) );
  nand2_1 U10426 ( .ip1(n8613), .ip2(n8608), .op(n8609) );
  nand2_1 U10427 ( .ip1(n8610), .ip2(n8609), .op(n11043) );
  inv_1 U10428 ( .ip(n11043), .op(n10408) );
  nor2_1 U10429 ( .ip1(n10408), .ip2(n10435), .op(n8611) );
  not_ab_or_c_or_d U10430 ( .ip1(n10906), .ip2(n10440), .ip3(n10376), .ip4(
        n8611), .op(n8618) );
  and3_1 U10431 ( .ip1(n8614), .ip2(n8613), .ip3(n8612), .op(n8616) );
  not_ab_or_c_or_d U10432 ( .ip1(n8782), .ip2(n9211), .ip3(n8616), .ip4(n8615), 
        .op(n11038) );
  inv_1 U10433 ( .ip(n11038), .op(n10391) );
  nand2_1 U10434 ( .ip1(n10391), .ip2(n10436), .op(n8617) );
  nand3_1 U10435 ( .ip1(n8619), .ip2(n8618), .ip3(n8617), .op(n11430) );
  nand2_1 U10436 ( .ip1(n10475), .ip2(n11430), .op(n8620) );
  nand4_1 U10437 ( .ip1(n10917), .ip2(n8622), .ip3(n8621), .ip4(n8620), .op(
        \CORTEXM0DS_INST/u_logic/Bmhvx4 ) );
  nor2_1 U10438 ( .ip1(n1156), .ip2(n12577), .op(n8623) );
  or2_1 U10439 ( .ip1(n12598), .ip2(n8623), .op(n8625) );
  or2_1 U10440 ( .ip1(\CORTEXM0DS_INST/u_logic/V6fvx4 ), .ip2(n8623), .op(
        n8624) );
  nand2_1 U10441 ( .ip1(n8625), .ip2(n8624), .op(n8628) );
  nand2_1 U10442 ( .ip1(n12603), .ip2(\CORTEXM0DS_INST/u_logic/Qufvx4 ), .op(
        n8627) );
  nand2_1 U10443 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n12575), .op(
        n8626) );
  nand4_1 U10444 ( .ip1(n1075), .ip2(n8628), .ip3(n8627), .ip4(n8626), .op(
        n6010) );
  nor2_1 U10445 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n8629), .op(
        n8631) );
  inv_1 U10446 ( .ip(\CORTEXM0DS_INST/u_logic/Xyfvx4 ), .op(n8630) );
  nor4_1 U10447 ( .ip1(n8631), .ip2(n12535), .ip3(n8630), .ip4(n12575), .op(
        n1147) );
  xor2_1 U10448 ( .ip1(n8633), .ip2(n8632), .op(n12282) );
  inv_1 U10449 ( .ip(n12282), .op(n11451) );
  nand2_1 U10450 ( .ip1(n11451), .ip2(n10916), .op(n8761) );
  nor2_1 U10451 ( .ip1(n8635), .ip2(n8634), .op(n10385) );
  or2_1 U10452 ( .ip1(n10385), .ip2(\CORTEXM0DS_INST/vis_pc [5]), .op(n8636)
         );
  nand2_1 U10453 ( .ip1(\CORTEXM0DS_INST/vis_pc [5]), .ip2(n10385), .op(n8846)
         );
  nand3_1 U10454 ( .ip1(n8636), .ip2(n12113), .ip3(n8846), .op(n8760) );
  nand2_1 U10455 ( .ip1(n9179), .ip2(n8776), .op(n8642) );
  nand2_1 U10456 ( .ip1(n9183), .ip2(n8637), .op(n8641) );
  nand2_1 U10457 ( .ip1(n9181), .ip2(n8773), .op(n8640) );
  nand2_1 U10458 ( .ip1(n9185), .ip2(n8638), .op(n8639) );
  nand4_1 U10459 ( .ip1(n8642), .ip2(n8641), .ip3(n8640), .ip4(n8639), .op(
        n9227) );
  nor2_1 U10460 ( .ip1(n8789), .ip2(n9156), .op(n8647) );
  nor2_1 U10461 ( .ip1(n8798), .ip2(n9243), .op(n8646) );
  nor2_1 U10462 ( .ip1(n8799), .ip2(n9158), .op(n8645) );
  inv_1 U10463 ( .ip(n8643), .op(n8788) );
  nor2_1 U10464 ( .ip1(n8788), .ip2(n9160), .op(n8644) );
  nor4_1 U10465 ( .ip1(n8647), .ip2(n8646), .ip3(n8645), .ip4(n8644), .op(
        n9219) );
  inv_1 U10466 ( .ip(n9219), .op(n10284) );
  mux2_1 U10467 ( .ip1(n9227), .ip2(n10284), .s(n8781), .op(n8649) );
  mux2_1 U10468 ( .ip1(n9244), .ip2(n9245), .s(n9228), .op(n8648) );
  mux2_1 U10469 ( .ip1(n9247), .ip2(n8649), .s(n8648), .op(n9249) );
  nand2_1 U10470 ( .ip1(n11853), .ip2(n9249), .op(n8665) );
  nand2_1 U10471 ( .ip1(n11863), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [22]), 
        .op(n8662) );
  nand4_1 U10472 ( .ip1(\CORTEXM0DS_INST/u_logic/L9hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Z7hvx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/B5hvx4 ), .ip4(n8651), .op(n8650) );
  nand2_1 U10473 ( .ip1(n12055), .ip2(n8650), .op(n11848) );
  nand2_1 U10474 ( .ip1(\CORTEXM0DS_INST/u_logic/L9hvx4 ), .ip2(n8651), .op(
        n8652) );
  nor3_1 U10475 ( .ip1(\CORTEXM0DS_INST/u_logic/Z7hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/B5hvx4 ), .ip3(n8652), .op(n12642) );
  nand2_1 U10476 ( .ip1(\CORTEXM0DS_INST/u_logic/Uth2z4 [0]), .ip2(n12642), 
        .op(n8656) );
  nand2_1 U10477 ( .ip1(n11841), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [6]), 
        .op(n8655) );
  nand2_1 U10478 ( .ip1(n11842), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [30]), 
        .op(n8654) );
  nand2_1 U10479 ( .ip1(n11864), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [14]), 
        .op(n8653) );
  nand4_1 U10480 ( .ip1(n8656), .ip2(n8655), .ip3(n8654), .ip4(n8653), .op(
        n8657) );
  not_ab_or_c_or_d U10481 ( .ip1(n8658), .ip2(n9134), .ip3(n11848), .ip4(n8657), .op(n8661) );
  nor4_1 U10482 ( .ip1(\CORTEXM0DS_INST/u_logic/B5hvx4 ), .ip2(n9146), .ip3(
        n11901), .ip4(n8659), .op(n12643) );
  nand2_1 U10483 ( .ip1(\CORTEXM0DS_INST/u_logic/Txh2z4 [0]), .ip2(n12643), 
        .op(n8660) );
  nand3_1 U10484 ( .ip1(n8662), .ip2(n8661), .ip3(n8660), .op(n8663) );
  nand2_1 U10485 ( .ip1(n8714), .ip2(n8663), .op(n8664) );
  nand3_1 U10486 ( .ip1(n8665), .ip2(n3485), .ip3(n8664), .op(n10596) );
  nand2_1 U10487 ( .ip1(n10906), .ip2(n10596), .op(n8758) );
  nand2_1 U10488 ( .ip1(n9181), .ip2(n8816), .op(n8669) );
  nand2_1 U10489 ( .ip1(n9183), .ip2(n9178), .op(n8668) );
  nand2_1 U10490 ( .ip1(n9179), .ip2(n9180), .op(n8667) );
  nand2_1 U10491 ( .ip1(n9185), .ip2(n9182), .op(n8666) );
  nand4_1 U10492 ( .ip1(n8669), .ip2(n8668), .ip3(n8667), .ip4(n8666), .op(
        n10253) );
  nand2_1 U10493 ( .ip1(n10285), .ip2(n10253), .op(n8689) );
  nor2_1 U10494 ( .ip1(n8670), .ip2(n9158), .op(n8677) );
  nor2_1 U10495 ( .ip1(n8671), .ip2(n9156), .op(n8676) );
  nor2_1 U10496 ( .ip1(n8672), .ip2(n9243), .op(n8675) );
  nor2_1 U10497 ( .ip1(n8673), .ip2(n9160), .op(n8674) );
  nor4_1 U10498 ( .ip1(n8677), .ip2(n8676), .ip3(n8675), .ip4(n8674), .op(
        n9232) );
  inv_1 U10499 ( .ip(n9232), .op(n9193) );
  nand2_1 U10500 ( .ip1(n11645), .ip2(n9193), .op(n8688) );
  nand2_1 U10501 ( .ip1(n8746), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [22]), 
        .op(n8681) );
  inv_1 U10502 ( .ip(n8906), .op(n11857) );
  nand2_1 U10503 ( .ip1(n11857), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [22]), 
        .op(n8680) );
  nand2_1 U10504 ( .ip1(n11863), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [20]), 
        .op(n8679) );
  nand2_1 U10505 ( .ip1(n11841), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [4]), 
        .op(n8678) );
  and4_1 U10506 ( .ip1(n8681), .ip2(n8680), .ip3(n8679), .ip4(n8678), .op(
        n8685) );
  nand2_1 U10507 ( .ip1(\CORTEXM0DS_INST/u_logic/Psh2z4 [0]), .ip2(n12643), 
        .op(n8684) );
  nand2_1 U10508 ( .ip1(n11864), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [12]), 
        .op(n8683) );
  nand2_1 U10509 ( .ip1(n11842), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [28]), 
        .op(n8682) );
  nand4_1 U10510 ( .ip1(n8685), .ip2(n8684), .ip3(n8683), .ip4(n8682), .op(
        n8686) );
  nand2_1 U10511 ( .ip1(n8714), .ip2(n8686), .op(n8687) );
  nand4_1 U10512 ( .ip1(n3554), .ip2(n8689), .ip3(n8688), .ip4(n8687), .op(
        n10592) );
  nand2_1 U10513 ( .ip1(n9183), .ip2(n8690), .op(n8697) );
  nand2_1 U10514 ( .ip1(n9181), .ip2(n8691), .op(n8696) );
  nand2_1 U10515 ( .ip1(n9179), .ip2(n8692), .op(n8695) );
  nand2_1 U10516 ( .ip1(n9185), .ip2(n8693), .op(n8694) );
  nand4_1 U10517 ( .ip1(n8697), .ip2(n8696), .ip3(n8695), .ip4(n8694), .op(
        n10263) );
  nand2_1 U10518 ( .ip1(n11645), .ip2(n10263), .op(n8717) );
  nand2_1 U10519 ( .ip1(n9183), .ip2(n9155), .op(n8703) );
  nand2_1 U10520 ( .ip1(n9181), .ip2(n8790), .op(n8702) );
  nand2_1 U10521 ( .ip1(n9179), .ip2(n8698), .op(n8701) );
  nand2_1 U10522 ( .ip1(n9185), .ip2(n8699), .op(n8700) );
  nand4_1 U10523 ( .ip1(n8703), .ip2(n8702), .ip3(n8701), .ip4(n8700), .op(
        n10277) );
  nand2_1 U10524 ( .ip1(n10285), .ip2(n10277), .op(n8716) );
  nand2_1 U10525 ( .ip1(n11870), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [6]), 
        .op(n8712) );
  inv_1 U10526 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [6]), .op(n11709) );
  nor2_1 U10527 ( .ip1(n11709), .ip2(n11860), .op(n8709) );
  nand2_1 U10528 ( .ip1(n11841), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [0]), 
        .op(n8707) );
  nand2_1 U10529 ( .ip1(n11864), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [8]), 
        .op(n8706) );
  nand2_1 U10530 ( .ip1(n11857), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [6]), 
        .op(n8705) );
  nand2_1 U10531 ( .ip1(n11842), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [24]), 
        .op(n8704) );
  nand4_1 U10532 ( .ip1(n8707), .ip2(n8706), .ip3(n8705), .ip4(n8704), .op(
        n8708) );
  not_ab_or_c_or_d U10533 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [6]), .ip2(
        n8746), .ip3(n8709), .ip4(n8708), .op(n8711) );
  nand2_1 U10534 ( .ip1(n11863), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [16]), 
        .op(n8710) );
  nand3_1 U10535 ( .ip1(n8712), .ip2(n8711), .ip3(n8710), .op(n8713) );
  nand2_1 U10536 ( .ip1(n8714), .ip2(n8713), .op(n8715) );
  and4_1 U10537 ( .ip1(n3514), .ip2(n8717), .ip3(n8716), .ip4(n8715), .op(
        n10588) );
  nor2_1 U10538 ( .ip1(n10588), .ip2(n10408), .op(n8756) );
  nand2_1 U10539 ( .ip1(n9179), .ip2(n8718), .op(n8723) );
  nand2_1 U10540 ( .ip1(n9181), .ip2(n8719), .op(n8722) );
  nand2_1 U10541 ( .ip1(n9183), .ip2(n8822), .op(n8721) );
  nand2_1 U10542 ( .ip1(n9185), .ip2(n8823), .op(n8720) );
  nand4_1 U10543 ( .ip1(n8723), .ip2(n8722), .ip3(n8721), .ip4(n8720), .op(
        n10269) );
  nor2_1 U10544 ( .ip1(n8724), .ip2(n9158), .op(n8730) );
  nor2_1 U10545 ( .ip1(n8725), .ip2(n9156), .op(n8729) );
  nor2_1 U10546 ( .ip1(n8821), .ip2(n9243), .op(n8728) );
  nor2_1 U10547 ( .ip1(n8726), .ip2(n9160), .op(n8727) );
  nor4_1 U10548 ( .ip1(n8730), .ip2(n8729), .ip3(n8728), .ip4(n8727), .op(
        n10255) );
  nor2_1 U10549 ( .ip1(n10255), .ip2(n10087), .op(n8754) );
  inv_1 U10550 ( .ip(n10122), .op(n10118) );
  nor2_1 U10551 ( .ip1(n8731), .ip2(n10118), .op(n8732) );
  or2_1 U10552 ( .ip1(n10114), .ip2(n8732), .op(n8734) );
  or2_1 U10553 ( .ip1(n10128), .ip2(n8732), .op(n8733) );
  nand2_1 U10554 ( .ip1(n8734), .ip2(n8733), .op(n8736) );
  inv_1 U10555 ( .ip(n8735), .op(n10131) );
  nor2_1 U10556 ( .ip1(n8736), .ip2(n10131), .op(n8737) );
  not_ab_or_c_or_d U10557 ( .ip1(n10103), .ip2(n8738), .ip3(n8737), .ip4(n8811), .op(n12470) );
  nand2_1 U10558 ( .ip1(n12470), .ip2(n10246), .op(n8752) );
  nor2_1 U10559 ( .ip1(n11856), .ip2(n8739), .op(n8745) );
  inv_1 U10560 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [14]), .op(n11726) );
  or2_1 U10561 ( .ip1(n11726), .ip2(n11860), .op(n8743) );
  nand2_1 U10562 ( .ip1(n11857), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [14]), 
        .op(n8742) );
  nand2_1 U10563 ( .ip1(n11863), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [18]), 
        .op(n8741) );
  nand2_1 U10564 ( .ip1(n11864), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [10]), 
        .op(n8740) );
  nand4_1 U10565 ( .ip1(n8743), .ip2(n8742), .ip3(n8741), .ip4(n8740), .op(
        n8744) );
  not_ab_or_c_or_d U10566 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [2]), .ip2(
        n11841), .ip3(n8745), .ip4(n8744), .op(n8749) );
  nand2_1 U10567 ( .ip1(n8746), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [14]), 
        .op(n8748) );
  not_ab_or_c_or_d U10568 ( .ip1(n8749), .ip2(n8748), .ip3(n8747), .ip4(n9712), 
        .op(n8750) );
  not_ab_or_c_or_d U10569 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [14]), .ip2(
        n11829), .ip3(n4241), .ip4(n8750), .op(n8751) );
  nand3_1 U10570 ( .ip1(n8752), .ip2(n8751), .ip3(n3420), .op(n8753) );
  not_ab_or_c_or_d U10571 ( .ip1(n10285), .ip2(n10269), .ip3(n8754), .ip4(
        n8753), .op(n10587) );
  nor2_1 U10572 ( .ip1(n10587), .ip2(n11038), .op(n8755) );
  not_ab_or_c_or_d U10573 ( .ip1(n10592), .ip2(n11037), .ip3(n8756), .ip4(
        n8755), .op(n8757) );
  nand3_1 U10574 ( .ip1(n8758), .ip2(n8757), .ip3(n11045), .op(n11449) );
  nand2_1 U10575 ( .ip1(n10475), .ip2(n11449), .op(n8759) );
  nand4_1 U10576 ( .ip1(n10917), .ip2(n8761), .ip3(n8760), .ip4(n8759), .op(
        \CORTEXM0DS_INST/u_logic/Glhvx4 ) );
  or2_1 U10577 ( .ip1(n10475), .ip2(n10467), .op(n8767) );
  nand4_1 U10578 ( .ip1(n8763), .ip2(n10586), .ip3(n8810), .ip4(n8762), .op(
        n8764) );
  nor3_1 U10579 ( .ip1(n8765), .ip2(n8782), .ip3(n8764), .op(n11355) );
  or2_1 U10580 ( .ip1(n11355), .ip2(n10467), .op(n8766) );
  nand2_1 U10581 ( .ip1(n8767), .ip2(n8766), .op(n10322) );
  nand2_1 U10582 ( .ip1(n9183), .ip2(n9184), .op(n8772) );
  nand2_1 U10583 ( .ip1(n9181), .ip2(n9178), .op(n8771) );
  nand2_1 U10584 ( .ip1(n9179), .ip2(n9182), .op(n8770) );
  nand2_1 U10585 ( .ip1(n9185), .ip2(n8768), .op(n8769) );
  nand4_1 U10586 ( .ip1(n8772), .ip2(n8771), .ip3(n8770), .ip4(n8769), .op(
        n10098) );
  nand2_1 U10587 ( .ip1(n9183), .ip2(n8773), .op(n8780) );
  nand2_1 U10588 ( .ip1(n9181), .ip2(n8774), .op(n8779) );
  nand2_1 U10589 ( .ip1(n9179), .ip2(n8775), .op(n8778) );
  nand2_1 U10590 ( .ip1(n9185), .ip2(n8776), .op(n8777) );
  nand4_1 U10591 ( .ip1(n8780), .ip2(n8779), .ip3(n8778), .ip4(n8777), .op(
        n9234) );
  mux2_1 U10592 ( .ip1(n10098), .ip2(n9234), .s(n8781), .op(n9685) );
  mux2_1 U10593 ( .ip1(n9685), .ip2(n9247), .s(n9229), .op(n9248) );
  not_ab_or_c_or_d U10594 ( .ip1(n11853), .ip2(n9248), .ip3(n3970), .ip4(n4241), .op(n11040) );
  inv_1 U10595 ( .ip(n11040), .op(n10468) );
  inv_1 U10596 ( .ip(n8782), .op(n8783) );
  nand2_1 U10597 ( .ip1(n8784), .ip2(n8783), .op(n10441) );
  nand2_1 U10598 ( .ip1(n10468), .ip2(n10441), .op(n8837) );
  inv_1 U10599 ( .ip(n10586), .op(n10452) );
  inv_1 U10600 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [0]), .op(n11716) );
  nor2_1 U10601 ( .ip1(n11716), .ip2(n11830), .op(n8785) );
  or2_1 U10602 ( .ip1(n10271), .ip2(n8785), .op(n8787) );
  or2_1 U10603 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [0]), .ip2(n8785), .op(
        n8786) );
  nand2_1 U10604 ( .ip1(n8787), .ip2(n8786), .op(n8808) );
  nor2_1 U10605 ( .ip1(n8788), .ip2(n9158), .op(n8795) );
  nor2_1 U10606 ( .ip1(n8789), .ip2(n9243), .op(n8794) );
  and2_1 U10607 ( .ip1(n8790), .ip2(n9183), .op(n8793) );
  nor2_1 U10608 ( .ip1(n8791), .ip2(n9160), .op(n8792) );
  nor4_1 U10609 ( .ip1(n8795), .ip2(n8794), .ip3(n8793), .ip4(n8792), .op(
        n10086) );
  nor2_1 U10610 ( .ip1(n8796), .ip2(n9158), .op(n8803) );
  nor2_1 U10611 ( .ip1(n8797), .ip2(n9243), .op(n8802) );
  nor2_1 U10612 ( .ip1(n8798), .ip2(n9156), .op(n8801) );
  nor2_1 U10613 ( .ip1(n8799), .ip2(n9160), .op(n8800) );
  nor4_1 U10614 ( .ip1(n8803), .ip2(n8802), .ip3(n8801), .ip4(n8800), .op(
        n9233) );
  mux2_1 U10615 ( .ip1(n10086), .ip2(n9233), .s(n10256), .op(n9680) );
  nor2_1 U10616 ( .ip1(n9680), .ip2(n11660), .op(n8805) );
  and2_1 U10617 ( .ip1(n8829), .ip2(\CORTEXM0DS_INST/u_logic/F2hvx4 ), .op(
        n8804) );
  not_ab_or_c_or_d U10618 ( .ip1(n10270), .ip2(
        \CORTEXM0DS_INST/u_logic/Czh2z4 [0]), .ip3(n8805), .ip4(n8804), .op(
        n8807) );
  nand2_1 U10619 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [0]), .ip2(n11829), 
        .op(n8806) );
  nand4_1 U10620 ( .ip1(n3973), .ip2(n8808), .ip3(n8807), .ip4(n8806), .op(
        n11044) );
  nand2_1 U10621 ( .ip1(n10452), .ip2(n11044), .op(n8836) );
  inv_1 U10622 ( .ip(n4286), .op(n10363) );
  nand2_1 U10623 ( .ip1(n8810), .ip2(n8809), .op(n10437) );
  nand2_1 U10624 ( .ip1(n10363), .ip2(n10437), .op(n8835) );
  nor2_1 U10625 ( .ip1(n8811), .ip2(n10131), .op(n12457) );
  nand2_1 U10626 ( .ip1(n10246), .ip2(n12457), .op(n8813) );
  nand2_1 U10627 ( .ip1(n10271), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [16]), 
        .op(n8812) );
  and4_1 U10628 ( .ip1(n3966), .ip2(n10259), .ip3(n8813), .ip4(n8812), .op(
        n8833) );
  nand2_1 U10629 ( .ip1(n9179), .ip2(n8814), .op(n8820) );
  nand2_1 U10630 ( .ip1(n9181), .ip2(n8815), .op(n8819) );
  nand2_1 U10631 ( .ip1(n9183), .ip2(n8816), .op(n8818) );
  nand2_1 U10632 ( .ip1(n9185), .ip2(n9180), .op(n8817) );
  nand4_1 U10633 ( .ip1(n8820), .ip2(n8819), .ip3(n8818), .ip4(n8817), .op(
        n10097) );
  or2_1 U10634 ( .ip1(n9156), .ip2(n8821), .op(n8828) );
  nand2_1 U10635 ( .ip1(n9181), .ip2(n8822), .op(n8827) );
  nand2_1 U10636 ( .ip1(n9179), .ip2(n8823), .op(n8826) );
  nand2_1 U10637 ( .ip1(n9185), .ip2(n8824), .op(n8825) );
  nand4_1 U10638 ( .ip1(n8828), .ip2(n8827), .ip3(n8826), .ip4(n8825), .op(
        n9167) );
  mux2_1 U10639 ( .ip1(n10097), .ip2(n9167), .s(n10256), .op(n9681) );
  nand2_1 U10640 ( .ip1(n9681), .ip2(n11853), .op(n8832) );
  nand2_1 U10641 ( .ip1(n10270), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [16]), 
        .op(n8831) );
  nand2_1 U10642 ( .ip1(\CORTEXM0DS_INST/u_logic/Izgvx4 ), .ip2(n8829), .op(
        n8830) );
  nand4_1 U10643 ( .ip1(n8833), .ip2(n8832), .ip3(n8831), .ip4(n8830), .op(
        n11036) );
  nand2_1 U10644 ( .ip1(n11036), .ip2(n10439), .op(n8834) );
  nand4_1 U10645 ( .ip1(n8837), .ip2(n8836), .ip3(n8835), .ip4(n8834), .op(
        n11356) );
  nand2_1 U10646 ( .ip1(n10475), .ip2(n11356), .op(n8843) );
  nor2_1 U10647 ( .ip1(n11005), .ip2(n10164), .op(n10163) );
  or2_1 U10648 ( .ip1(\CORTEXM0DS_INST/vis_pc [15]), .ip2(n10163), .op(n8838)
         );
  nand2_1 U10649 ( .ip1(\CORTEXM0DS_INST/vis_pc [15]), .ip2(n10163), .op(
        n10313) );
  nand3_1 U10650 ( .ip1(n12113), .ip2(n8838), .ip3(n10313), .op(n8842) );
  xor2_1 U10651 ( .ip1(n8840), .ip2(n8839), .op(n11357) );
  nand2_1 U10652 ( .ip1(n11357), .ip2(n10916), .op(n8841) );
  nand4_1 U10653 ( .ip1(n10322), .ip2(n8843), .ip3(n8842), .ip4(n8841), .op(
        \CORTEXM0DS_INST/u_logic/Qjhvx4 ) );
  xor2_1 U10654 ( .ip1(n8845), .ip2(n8844), .op(n12339) );
  nand2_1 U10655 ( .ip1(n12339), .ip2(n10916), .op(n8854) );
  inv_1 U10656 ( .ip(\CORTEXM0DS_INST/vis_pc [6]), .op(n12335) );
  nand2_1 U10657 ( .ip1(n8846), .ip2(n12335), .op(n8847) );
  nand3_1 U10658 ( .ip1(\CORTEXM0DS_INST/vis_pc [5]), .ip2(
        \CORTEXM0DS_INST/vis_pc [6]), .ip3(n10385), .op(n10360) );
  nand3_1 U10659 ( .ip1(n8847), .ip2(n12113), .ip3(n10360), .op(n8853) );
  nand2_1 U10660 ( .ip1(n10391), .ip2(n10451), .op(n8851) );
  nor2_1 U10661 ( .ip1(n4130), .ip2(n11039), .op(n8849) );
  nor2_1 U10662 ( .ip1(n4149), .ip2(n10408), .op(n8848) );
  not_ab_or_c_or_d U10663 ( .ip1(n10454), .ip2(n11037), .ip3(n8849), .ip4(
        n8848), .op(n8850) );
  nand3_1 U10664 ( .ip1(n8851), .ip2(n8850), .ip3(n11045), .op(n11513) );
  nand2_1 U10665 ( .ip1(n10475), .ip2(n11513), .op(n8852) );
  nand4_1 U10666 ( .ip1(n10917), .ip2(n8854), .ip3(n8853), .ip4(n8852), .op(
        \CORTEXM0DS_INST/u_logic/Zkhvx4 ) );
  nand2_1 U10667 ( .ip1(\CORTEXM0DS_INST/u_logic/E1dvx4 ), .ip2(n2119), .op(
        n8864) );
  nand2_1 U10668 ( .ip1(\CORTEXM0DS_INST/vis_pc [1]), .ip2(n12359), .op(n8863)
         );
  nand2_1 U10669 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [2]), .ip2(n12358), .op(
        n8862) );
  xor2_1 U10670 ( .ip1(n8856), .ip2(n8855), .op(n10418) );
  inv_1 U10671 ( .ip(n12316), .op(n12347) );
  nor2_1 U10672 ( .ip1(n11760), .ip2(n12347), .op(n8860) );
  not_ab_or_c_or_d U10673 ( .ip1(n8858), .ip2(n12401), .ip3(n8857), .ip4(
        n12343), .op(n8859) );
  not_ab_or_c_or_d U10674 ( .ip1(n12352), .ip2(n10418), .ip3(n8860), .ip4(
        n8859), .op(\CORTEXM0DS_INST/u_logic/Fvovx4 ) );
  inv_1 U10675 ( .ip(\CORTEXM0DS_INST/u_logic/Fvovx4 ), .op(n1850) );
  nand2_1 U10676 ( .ip1(n2118), .ip2(n1850), .op(n8861) );
  nand4_1 U10677 ( .ip1(n8864), .ip2(n8863), .ip3(n8862), .ip4(n8861), .op(
        n6075) );
  nand2_1 U10678 ( .ip1(\CORTEXM0DS_INST/vis_pc [2]), .ip2(n12359), .op(n8868)
         );
  nand2_1 U10679 ( .ip1(\CORTEXM0DS_INST/u_logic/O2dvx4 ), .ip2(n2119), .op(
        n8867) );
  nand2_1 U10680 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [3]), .ip2(n12358), .op(
        n8866) );
  or2_1 U10681 ( .ip1(n12355), .ip2(\CORTEXM0DS_INST/u_logic/Ekovx4 ), .op(
        n8865) );
  nand4_1 U10682 ( .ip1(n8868), .ip2(n8867), .ip3(n8866), .ip4(n8865), .op(
        n6085) );
  nand2_1 U10683 ( .ip1(\CORTEXM0DS_INST/vis_pc [3]), .ip2(n12359), .op(n8878)
         );
  nand2_1 U10684 ( .ip1(\CORTEXM0DS_INST/u_logic/Y3dvx4 ), .ip2(n2119), .op(
        n8877) );
  nand2_1 U10685 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [4]), .ip2(n12358), .op(
        n8876) );
  xor2_1 U10686 ( .ip1(n8870), .ip2(n8869), .op(n11437) );
  inv_1 U10687 ( .ip(\CORTEXM0DS_INST/vis_pc [3]), .op(n10401) );
  inv_1 U10688 ( .ip(n8871), .op(n8872) );
  nor2_1 U10689 ( .ip1(n10401), .ip2(n8872), .op(n8879) );
  not_ab_or_c_or_d U10690 ( .ip1(n10401), .ip2(n8872), .ip3(n8879), .ip4(
        n12343), .op(n8874) );
  nor2_1 U10691 ( .ip1(n9571), .ip2(n12347), .op(n8873) );
  not_ab_or_c_or_d U10692 ( .ip1(n12352), .ip2(n11437), .ip3(n8874), .ip4(
        n8873), .op(\CORTEXM0DS_INST/u_logic/Yuovx4 ) );
  inv_1 U10693 ( .ip(\CORTEXM0DS_INST/u_logic/Yuovx4 ), .op(n1943) );
  nand2_1 U10694 ( .ip1(n2118), .ip2(n1943), .op(n8875) );
  nand4_1 U10695 ( .ip1(n8878), .ip2(n8877), .ip3(n8876), .ip4(n8875), .op(
        n6084) );
  nand2_1 U10696 ( .ip1(\CORTEXM0DS_INST/u_logic/I5dvx4 ), .ip2(n2119), .op(
        n8889) );
  nand2_1 U10697 ( .ip1(\CORTEXM0DS_INST/vis_pc [4]), .ip2(n12359), .op(n8888)
         );
  nand2_1 U10698 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [5]), .ip2(n12358), .op(
        n8887) );
  inv_1 U10699 ( .ip(n9458), .op(n9462) );
  nor2_1 U10700 ( .ip1(\CORTEXM0DS_INST/vis_pc [4]), .ip2(n8879), .op(n8881)
         );
  inv_1 U10701 ( .ip(n12281), .op(n8880) );
  nor3_1 U10702 ( .ip1(n8881), .ip2(n8880), .ip3(n12343), .op(n8885) );
  xor2_1 U10703 ( .ip1(n8883), .ip2(n8882), .op(n10384) );
  nor2_1 U10704 ( .ip1(n10384), .ip2(n12311), .op(n8884) );
  not_ab_or_c_or_d U10705 ( .ip1(n12316), .ip2(n9462), .ip3(n8885), .ip4(n8884), .op(\CORTEXM0DS_INST/u_logic/Rxzvx4 ) );
  or2_1 U10706 ( .ip1(\CORTEXM0DS_INST/u_logic/Rxzvx4 ), .ip2(n12355), .op(
        n8886) );
  nand4_1 U10707 ( .ip1(n8889), .ip2(n8888), .ip3(n8887), .ip4(n8886), .op(
        n6083) );
  inv_1 U10708 ( .ip(n10437), .op(n10314) );
  nor2_1 U10709 ( .ip1(n10587), .ip2(n10314), .op(n8891) );
  nor2_1 U10710 ( .ip1(n10588), .ip2(n10586), .op(n8890) );
  not_ab_or_c_or_d U10711 ( .ip1(n10596), .ip2(n10441), .ip3(n8891), .ip4(
        n8890), .op(n8893) );
  nand2_1 U10712 ( .ip1(n10592), .ip2(n10439), .op(n8892) );
  nand2_1 U10713 ( .ip1(n8893), .ip2(n8892), .op(n11419) );
  nand2_1 U10714 ( .ip1(n10475), .ip2(n11419), .op(n8901) );
  nor2_1 U10715 ( .ip1(n8894), .ip2(n10164), .op(n10179) );
  nand2_1 U10716 ( .ip1(\CORTEXM0DS_INST/vis_pc [20]), .ip2(n10179), .op(n8895) );
  inv_1 U10717 ( .ip(\CORTEXM0DS_INST/vis_pc [21]), .op(n12272) );
  nand2_1 U10718 ( .ip1(n8895), .ip2(n12272), .op(n8896) );
  nand3_1 U10719 ( .ip1(\CORTEXM0DS_INST/vis_pc [20]), .ip2(
        \CORTEXM0DS_INST/vis_pc [21]), .ip3(n10179), .op(n10169) );
  nand3_1 U10720 ( .ip1(n8896), .ip2(n12113), .ip3(n10169), .op(n8900) );
  xor2_1 U10721 ( .ip1(n8898), .ip2(n8897), .op(n12276) );
  nand2_1 U10722 ( .ip1(n12276), .ip2(n10916), .op(n8899) );
  nand4_1 U10723 ( .ip1(n10322), .ip2(n8901), .ip3(n8900), .ip4(n8899), .op(
        \CORTEXM0DS_INST/u_logic/Vihvx4 ) );
  nand2_1 U10724 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [8]), .ip2(n11829), 
        .op(n8905) );
  nand2_1 U10725 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [8]), .ip2(n10272), 
        .op(n8904) );
  nand2_1 U10726 ( .ip1(n10270), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [8]), 
        .op(n8903) );
  nand2_1 U10727 ( .ip1(n10271), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [8]), 
        .op(n8902) );
  nand4_1 U10728 ( .ip1(n8905), .ip2(n8904), .ip3(n8903), .ip4(n8902), .op(
        n3958) );
  buf_1 U10729 ( .ip(n12697), .op(n12732) );
  buf_1 U10730 ( .ip(n12718), .op(n12734) );
  inv_1 U10731 ( .ip(\CORTEXM0DS_INST/u_logic/Mf8vx4 ), .op(n12687) );
  nor2_1 U10732 ( .ip1(n8906), .ip2(n12687), .op(n12691) );
  buf_1 U10733 ( .ip(n12691), .op(n12692) );
  buf_1 U10734 ( .ip(n12699), .op(n12694) );
  buf_1 U10735 ( .ip(n12703), .op(n12693) );
  nand4_1 U10736 ( .ip1(n3227), .ip2(n3226), .ip3(n3229), .ip4(n3228), .op(
        n3230) );
  nand2_1 U10737 ( .ip1(\CORTEXM0DS_INST/u_logic/D6evx4 ), .ip2(n2119), .op(
        n8909) );
  nand2_1 U10738 ( .ip1(\CORTEXM0DS_INST/vis_pc [30]), .ip2(n12359), .op(n8908) );
  nand2_1 U10739 ( .ip1(\CORTEXM0DS_INST/vis_apsr [3]), .ip2(n12358), .op(
        n8907) );
  nand4_1 U10740 ( .ip1(n2121), .ip2(n8909), .ip3(n8908), .ip4(n8907), .op(
        n6102) );
  nand2_1 U10741 ( .ip1(\CORTEXM0DS_INST/u_logic/S4evx4 ), .ip2(n2119), .op(
        n8912) );
  nand2_1 U10742 ( .ip1(\CORTEXM0DS_INST/vis_pc [29]), .ip2(n12359), .op(n8911) );
  nand2_1 U10743 ( .ip1(\CORTEXM0DS_INST/vis_apsr [2]), .ip2(n12358), .op(
        n8910) );
  nand4_1 U10744 ( .ip1(n1869), .ip2(n8912), .ip3(n8911), .ip4(n8910), .op(
        n6078) );
  nand2_1 U10745 ( .ip1(\CORTEXM0DS_INST/u_logic/H3evx4 ), .ip2(n2119), .op(
        n8915) );
  nand2_1 U10746 ( .ip1(\CORTEXM0DS_INST/vis_pc [28]), .ip2(n12359), .op(n8914) );
  nand2_1 U10747 ( .ip1(\CORTEXM0DS_INST/vis_apsr [1]), .ip2(n12358), .op(
        n8913) );
  nand4_1 U10748 ( .ip1(n1812), .ip2(n8915), .ip3(n8914), .ip4(n8913), .op(
        n6072) );
  inv_1 U10749 ( .ip(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .op(n12413) );
  nor2_1 U10750 ( .ip1(n10028), .ip2(n12413), .op(n12683) );
  inv_1 U10751 ( .ip(n11052), .op(n11508) );
  and2_1 U10752 ( .ip1(n10028), .ip2(n8917), .op(
        \CORTEXM0DS_INST/u_logic/Oq42z4 ) );
  nand2_1 U10753 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Oq42z4 ), .op(n10076) );
  nor2_1 U10754 ( .ip1(n11315), .ip2(n10076), .op(n8919) );
  nor3_1 U10755 ( .ip1(n8917), .ip2(n8916), .ip3(n12413), .op(n12664) );
  nand2_1 U10756 ( .ip1(n12664), .ip2(n12675), .op(n5990) );
  inv_1 U10757 ( .ip(n5990), .op(n8918) );
  not_ab_or_c_or_d U10758 ( .ip1(n12683), .ip2(n11508), .ip3(n8919), .ip4(
        n8918), .op(\CORTEXM0DS_INST/u_logic/Sx3wx4 ) );
  mux2_1 U10759 ( .ip1(n10058), .ip2(n9612), .s(n12683), .op(
        \CORTEXM0DS_INST/u_logic/O24wx4 ) );
  inv_1 U10760 ( .ip(n8942), .op(n12652) );
  nor2_1 U10761 ( .ip1(n8920), .ip2(n12652), .op(n8921) );
  or2_1 U10762 ( .ip1(\CORTEXM0DS_INST/u_logic/Eqgvx4 ), .ip2(n8921), .op(
        n8923) );
  or2_1 U10763 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [0]), .ip2(n8921), .op(n8922)
         );
  nand2_1 U10764 ( .ip1(n8923), .ip2(n8922), .op(n8973) );
  or2_1 U10765 ( .ip1(\CORTEXM0DS_INST/u_logic/Uth2z4 [0]), .ip2(n8924), .op(
        n8926) );
  or2_1 U10766 ( .ip1(n11884), .ip2(n8924), .op(n8925) );
  nand2_1 U10767 ( .ip1(n8926), .ip2(n8925), .op(n8929) );
  nor2_1 U10768 ( .ip1(n8927), .ip2(n10138), .op(n8928) );
  not_ab_or_c_or_d U10769 ( .ip1(n10138), .ip2(n8930), .ip3(n8929), .ip4(n8928), .op(n8940) );
  inv_1 U10770 ( .ip(n8931), .op(n8933) );
  mux2_1 U10771 ( .ip1(n8933), .ip2(n8932), .s(n10138), .op(n8939) );
  inv_1 U10772 ( .ip(n8934), .op(n8936) );
  nor2_1 U10773 ( .ip1(n8939), .ip2(n8940), .op(n8935) );
  nor2_1 U10774 ( .ip1(n8936), .ip2(n8935), .op(n8938) );
  ab_or_c_or_d U10775 ( .ip1(n8940), .ip2(n8939), .ip3(n8938), .ip4(n8937), 
        .op(n8941) );
  nand3_1 U10776 ( .ip1(n8942), .ip2(n8941), .ip3(n10104), .op(n8943) );
  nand2_1 U10777 ( .ip1(n8973), .ip2(n8943), .op(n5656) );
  nand4_1 U10778 ( .ip1(\CORTEXM0DS_INST/u_logic/I4gvx4 ), .ip2(n12112), .ip3(
        n9807), .ip4(n12536), .op(n11029) );
  or2_1 U10779 ( .ip1(n8944), .ip2(n12117), .op(n8953) );
  nand2_1 U10780 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .op(n9838) );
  nor2_1 U10781 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n12623), .op(
        n10701) );
  or2_1 U10782 ( .ip1(n9838), .ip2(n10701), .op(n8946) );
  or2_1 U10783 ( .ip1(n11681), .ip2(n10701), .op(n8945) );
  nand2_1 U10784 ( .ip1(n8946), .ip2(n8945), .op(n8952) );
  nor3_1 U10785 ( .ip1(n12609), .ip2(n11693), .ip3(n11793), .op(n8947) );
  nor3_1 U10786 ( .ip1(n8947), .ip2(n9385), .ip3(n11258), .op(n8950) );
  nand3_1 U10787 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n10632), .ip3(
        n11228), .op(n8949) );
  nand3_1 U10788 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(n9730), .ip3(
        n12118), .op(n8948) );
  nand4_1 U10789 ( .ip1(n8950), .ip2(n11754), .ip3(n8949), .ip4(n8948), .op(
        n8951) );
  not_ab_or_c_or_d U10790 ( .ip1(n12610), .ip2(n8953), .ip3(n8952), .ip4(n8951), .op(n11283) );
  nor2_1 U10791 ( .ip1(n11283), .ip2(n9091), .op(n8965) );
  nor2_1 U10792 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Whgvx4 ), .op(n12116) );
  nand2_1 U10793 ( .ip1(n12116), .ip2(n11679), .op(n9737) );
  inv_1 U10794 ( .ip(n9737), .op(n8958) );
  nor3_1 U10795 ( .ip1(n12117), .ip2(n12623), .ip3(n9956), .op(n8957) );
  nor2_1 U10796 ( .ip1(n11682), .ip2(n11681), .op(n11678) );
  inv_1 U10797 ( .ip(n12131), .op(n10962) );
  nor2_1 U10798 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n12627), .op(
        n12611) );
  nor2_1 U10799 ( .ip1(n11693), .ip2(n11232), .op(n8954) );
  not_ab_or_c_or_d U10800 ( .ip1(n10962), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip3(n12611), .ip4(n8954), .op(
        n8955) );
  nor2_1 U10801 ( .ip1(n8955), .ip2(n9807), .op(n8956) );
  nor4_1 U10802 ( .ip1(n8958), .ip2(n8957), .ip3(n11678), .ip4(n8956), .op(
        n11284) );
  nor2_1 U10803 ( .ip1(n11284), .ip2(n12373), .op(n8964) );
  nor2_1 U10804 ( .ip1(n12117), .ip2(n10988), .op(n12617) );
  nor3_1 U10805 ( .ip1(n9943), .ip2(n11683), .ip3(n10740), .op(n8959) );
  not_ab_or_c_or_d U10806 ( .ip1(n8960), .ip2(n9853), .ip3(n12617), .ip4(n8959), .op(n11285) );
  nor2_1 U10807 ( .ip1(n11285), .ip2(n9010), .op(n8963) );
  nand3_1 U10808 ( .ip1(n9807), .ip2(n9657), .ip3(
        \CORTEXM0DS_INST/u_logic/Efgvx4 ), .op(n8962) );
  nand2_1 U10809 ( .ip1(n8962), .ip2(n8961), .op(n11282) );
  nor4_1 U10810 ( .ip1(n8965), .ip2(n8964), .ip3(n8963), .ip4(n11282), .op(
        n11601) );
  nor4_1 U10811 ( .ip1(n11601), .ip2(n12131), .ip3(n12623), .ip4(n10673), .op(
        n8970) );
  inv_1 U10812 ( .ip(n9798), .op(n10610) );
  nor2_1 U10813 ( .ip1(n10610), .ip2(n10687), .op(n8966) );
  or2_1 U10814 ( .ip1(n10813), .ip2(n8966), .op(n8968) );
  or2_1 U10815 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n8966), .op(
        n8967) );
  nand2_1 U10816 ( .ip1(n8968), .ip2(n8967), .op(n11812) );
  nor2_1 U10817 ( .ip1(n11812), .ip2(n11516), .op(n8969) );
  nor2_1 U10818 ( .ip1(n8970), .ip2(n8969), .op(n12436) );
  nor2_1 U10819 ( .ip1(n12131), .ip2(n10673), .op(n8972) );
  nor2_1 U10820 ( .ip1(n10058), .ip2(n11812), .op(n8971) );
  not_ab_or_c_or_d U10821 ( .ip1(n8972), .ip2(\CORTEXM0DS_INST/u_logic/Fs8vx4 ), .ip3(n12436), .ip4(n8971), .op(n12439) );
  inv_1 U10822 ( .ip(n8973), .op(n8974) );
  ab_or_c_or_d U10823 ( .ip1(n12436), .ip2(n11515), .ip3(n12439), .ip4(n8974), 
        .op(n8975) );
  nand2_1 U10824 ( .ip1(n5656), .ip2(n8975), .op(n12064) );
  inv_1 U10825 ( .ip(\CORTEXM0DS_INST/u_logic/Xlevx4 ), .op(n12453) );
  nand2_1 U10826 ( .ip1(n12064), .ip2(n12453), .op(n9106) );
  or2_1 U10827 ( .ip1(n11029), .ip2(n9106), .op(n8978) );
  nand3_1 U10828 ( .ip1(n12112), .ip2(\CORTEXM0DS_INST/u_logic/V8evx4 ), .ip3(
        n12575), .op(n8976) );
  or2_1 U10829 ( .ip1(n8976), .ip2(n9106), .op(n8977) );
  nand2_1 U10830 ( .ip1(n8978), .ip2(n8977), .op(n6042) );
  nor2_1 U10831 ( .ip1(n12571), .ip2(n11089), .op(n9008) );
  inv_1 U10832 ( .ip(n10973), .op(n8979) );
  or2_1 U10833 ( .ip1(n8979), .ip2(n11779), .op(n8980) );
  nand2_1 U10834 ( .ip1(n10782), .ip2(n8980), .op(n12099) );
  inv_1 U10835 ( .ip(n12099), .op(n8981) );
  not_ab_or_c_or_d U10836 ( .ip1(n11108), .ip2(n9008), .ip3(n1769), .ip4(n8981), .op(n12392) );
  nand3_1 U10837 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n9807), .ip3(
        n12125), .op(n10885) );
  inv_1 U10838 ( .ip(n10885), .op(n10732) );
  or2_1 U10839 ( .ip1(n8982), .ip2(n10732), .op(n8983) );
  nand2_1 U10840 ( .ip1(n8983), .ip2(n12125), .op(n12386) );
  nand3_1 U10841 ( .ip1(n10206), .ip2(n10647), .ip3(n10818), .op(n8987) );
  nand2_1 U10842 ( .ip1(n10818), .ip2(n11090), .op(n10218) );
  inv_1 U10843 ( .ip(n10218), .op(n8985) );
  nor2_1 U10844 ( .ip1(n12592), .ip2(n10820), .op(n9882) );
  inv_1 U10845 ( .ip(n9882), .op(n10964) );
  nand2_1 U10846 ( .ip1(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip2(n10964), .op(
        n8984) );
  nand2_1 U10847 ( .ip1(n8985), .ip2(n8984), .op(n12385) );
  nand4_1 U10848 ( .ip1(n12386), .ip2(n8987), .ip3(n12385), .ip4(n8986), .op(
        n12374) );
  nand2_1 U10849 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n12374), .op(
        n8995) );
  nand2_1 U10850 ( .ip1(\CORTEXM0DS_INST/u_logic/R89vx4 ), .ip2(n12389), .op(
        n8994) );
  inv_1 U10851 ( .ip(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .op(n12583) );
  nor2_1 U10852 ( .ip1(n12592), .ip2(n12583), .op(n10724) );
  nand2_1 U10853 ( .ip1(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip2(n10481), .op(
        n9808) );
  nor3_1 U10854 ( .ip1(n10724), .ip2(n10218), .ip3(n9808), .op(n8988) );
  or2_1 U10855 ( .ip1(n11181), .ip2(n8988), .op(n8990) );
  or2_1 U10856 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(n8988), .op(
        n8989) );
  nand2_1 U10857 ( .ip1(n8990), .ip2(n8989), .op(n12390) );
  nand3_1 U10858 ( .ip1(n10647), .ip2(n10818), .ip3(n12599), .op(n11096) );
  inv_1 U10859 ( .ip(n9834), .op(n9869) );
  nand3_1 U10860 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n9870), .ip3(
        n9869), .op(n8992) );
  inv_1 U10861 ( .ip(n11090), .op(n10646) );
  nor2_1 U10862 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n10646), .op(
        n9899) );
  nand2_1 U10863 ( .ip1(n10818), .ip2(n9899), .op(n11105) );
  or2_1 U10864 ( .ip1(n12599), .ip2(n11105), .op(n8991) );
  nand4_1 U10865 ( .ip1(n12390), .ip2(n11096), .ip3(n8992), .ip4(n8991), .op(
        n12375) );
  nand2_1 U10866 ( .ip1(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), .ip2(n12375), .op(
        n8993) );
  and4_1 U10867 ( .ip1(n12392), .ip2(n8995), .ip3(n8994), .ip4(n8993), .op(
        n8996) );
  or2_1 U10868 ( .ip1(n1769), .ip2(n8996), .op(n8998) );
  or2_1 U10869 ( .ip1(n11206), .ip2(n8996), .op(n8997) );
  nand2_1 U10870 ( .ip1(n8998), .ip2(n8997), .op(n6067) );
  inv_1 U10871 ( .ip(n10041), .op(n1520) );
  nor2_1 U10872 ( .ip1(n11786), .ip2(n11789), .op(n10863) );
  nor3_1 U10873 ( .ip1(n10863), .ip2(n3348), .ip3(n10798), .op(n9006) );
  not_ab_or_c_or_d U10874 ( .ip1(n12384), .ip2(n12362), .ip3(
        \CORTEXM0DS_INST/u_logic/Ot9vx4 ), .ip4(
        \CORTEXM0DS_INST/u_logic/Su9vx4 ), .op(n8999) );
  nor2_1 U10875 ( .ip1(n9000), .ip2(n8999), .op(n9001) );
  nor2_1 U10876 ( .ip1(n10739), .ip2(n9001), .op(n9004) );
  nor2_1 U10877 ( .ip1(n12588), .ip2(n10646), .op(n9002) );
  nor2_1 U10878 ( .ip1(n10551), .ip2(n9002), .op(n9040) );
  nor2_1 U10879 ( .ip1(n9040), .ip2(n9881), .op(n9003) );
  not_ab_or_c_or_d U10880 ( .ip1(n9899), .ip2(\CORTEXM0DS_INST/u_logic/B19vx4 ), .ip3(n9004), .ip4(n9003), .op(n9005) );
  nand2_1 U10881 ( .ip1(n9006), .ip2(n9005), .op(n9007) );
  not_ab_or_c_or_d U10882 ( .ip1(n12653), .ip2(
        \CORTEXM0DS_INST/u_logic/Su9vx4 ), .ip3(n9008), .ip4(n9007), .op(n9009) );
  or2_1 U10883 ( .ip1(n3348), .ip2(n9009), .op(n9012) );
  or2_1 U10884 ( .ip1(n9010), .ip2(n9009), .op(n9011) );
  nand2_1 U10885 ( .ip1(n9012), .ip2(n9011), .op(
        \CORTEXM0DS_INST/u_logic/G2mvx4 ) );
  nor2_1 U10886 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n12623), .op(
        n9013) );
  nor4_1 U10887 ( .ip1(n9013), .ip2(n10863), .ip3(n3348), .ip4(n10798), .op(
        n9048) );
  inv_1 U10888 ( .ip(n9014), .op(n9021) );
  inv_1 U10889 ( .ip(\CORTEXM0DS_INST/u_logic/Ks9vx4 ), .op(n9015) );
  nor2_1 U10890 ( .ip1(n9043), .ip2(n9015), .op(n9020) );
  or2_1 U10891 ( .ip1(\CORTEXM0DS_INST/u_logic/Bx9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Su9vx4 ), .op(n9017) );
  or2_1 U10892 ( .ip1(n12362), .ip2(\CORTEXM0DS_INST/u_logic/Su9vx4 ), .op(
        n9016) );
  nand2_1 U10893 ( .ip1(n9017), .ip2(n9016), .op(n9018) );
  nor2_1 U10894 ( .ip1(\CORTEXM0DS_INST/u_logic/Ot9vx4 ), .ip2(n9018), .op(
        n9019) );
  not_ab_or_c_or_d U10895 ( .ip1(\CORTEXM0DS_INST/u_logic/Cq9vx4 ), .ip2(n9021), .ip3(n9020), .ip4(n9019), .op(n9022) );
  nor2_1 U10896 ( .ip1(n9022), .ip2(n10739), .op(n9024) );
  nor2_1 U10897 ( .ip1(n9040), .ip2(n12558), .op(n9023) );
  not_ab_or_c_or_d U10898 ( .ip1(n11146), .ip2(
        \CORTEXM0DS_INST/u_logic/K79vx4 ), .ip3(n9024), .ip4(n9023), .op(n9027) );
  nand2_1 U10899 ( .ip1(\CORTEXM0DS_INST/u_logic/Ot9vx4 ), .ip2(n12653), .op(
        n9026) );
  nand2_1 U10900 ( .ip1(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), .ip2(n9899), .op(
        n9025) );
  and4_1 U10901 ( .ip1(n9048), .ip2(n9027), .ip3(n9026), .ip4(n9025), .op(
        n9028) );
  or2_1 U10902 ( .ip1(n3348), .ip2(n9028), .op(n9030) );
  or2_1 U10903 ( .ip1(n11205), .ip2(n9028), .op(n9029) );
  nand2_1 U10904 ( .ip1(n9030), .ip2(n9029), .op(
        \CORTEXM0DS_INST/u_logic/Kuhvx4 ) );
  nor2_1 U10905 ( .ip1(n9040), .ip2(n12562), .op(n9035) );
  nand2_1 U10906 ( .ip1(\CORTEXM0DS_INST/u_logic/Wv9vx4 ), .ip2(n12653), .op(
        n9033) );
  nand2_1 U10907 ( .ip1(n9044), .ip2(n10203), .op(n9032) );
  nand2_1 U10908 ( .ip1(\CORTEXM0DS_INST/u_logic/I29vx4 ), .ip2(n9899), .op(
        n9031) );
  nand4_1 U10909 ( .ip1(n9048), .ip2(n9033), .ip3(n9032), .ip4(n9031), .op(
        n9034) );
  not_ab_or_c_or_d U10910 ( .ip1(n11146), .ip2(
        \CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip3(n9035), .ip4(n9034), .op(n9036) );
  or2_1 U10911 ( .ip1(n3348), .ip2(n9036), .op(n9039) );
  or2_1 U10912 ( .ip1(n9037), .ip2(n9036), .op(n9038) );
  nand2_1 U10913 ( .ip1(n9039), .ip2(n9038), .op(
        \CORTEXM0DS_INST/u_logic/Pfhvx4 ) );
  nor3_1 U10914 ( .ip1(n9040), .ip2(n12567), .ip3(n12588), .op(n9042) );
  nor2_1 U10915 ( .ip1(n12384), .ip2(n10865), .op(n9041) );
  not_ab_or_c_or_d U10916 ( .ip1(n9899), .ip2(\CORTEXM0DS_INST/u_logic/P39vx4 ), .ip3(n9042), .ip4(n9041), .op(n9047) );
  nor2_1 U10917 ( .ip1(\CORTEXM0DS_INST/u_logic/Ks9vx4 ), .ip2(n9043), .op(
        n10670) );
  nand2_1 U10918 ( .ip1(n10203), .ip2(n10670), .op(n9046) );
  nand4_1 U10919 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip3(n9044), .ip4(n10203), .op(
        n9045) );
  and4_1 U10920 ( .ip1(n9048), .ip2(n9047), .ip3(n9046), .ip4(n9045), .op(
        n9049) );
  or2_1 U10921 ( .ip1(n3348), .ip2(n9049), .op(n9052) );
  or2_1 U10922 ( .ip1(n9050), .ip2(n9049), .op(n9051) );
  nand2_1 U10923 ( .ip1(n9052), .ip2(n9051), .op(
        \CORTEXM0DS_INST/u_logic/Ifhvx4 ) );
  inv_1 U10924 ( .ip(n12072), .op(n10619) );
  or2_1 U10925 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n10619), .op(
        n9054) );
  nor4_1 U10926 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(n10492), .ip3(
        n9869), .ip4(n10782), .op(n9056) );
  or2_1 U10927 ( .ip1(n9056), .ip2(n10619), .op(n9053) );
  nand2_1 U10928 ( .ip1(n9054), .ip2(n9053), .op(n9055) );
  nor2_1 U10929 ( .ip1(n12571), .ip2(n9055), .op(n9063) );
  nor3_1 U10930 ( .ip1(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), .ip2(n12558), .ip3(
        n12072), .op(n11768) );
  inv_1 U10931 ( .ip(\CORTEXM0DS_INST/u_logic/B19vx4 ), .op(n12548) );
  inv_1 U10932 ( .ip(n10820), .op(n10636) );
  nor2_1 U10933 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n10636), .op(
        n9756) );
  nand2_1 U10934 ( .ip1(n12592), .ip2(n11190), .op(n10930) );
  inv_1 U10935 ( .ip(n10930), .op(n9057) );
  inv_1 U10936 ( .ip(n9056), .op(n9072) );
  nor3_1 U10937 ( .ip1(n9756), .ip2(n9057), .ip3(n9072), .op(n9058) );
  not_ab_or_c_or_d U10938 ( .ip1(n11768), .ip2(n12548), .ip3(n9058), .ip4(
        n3393), .op(n9086) );
  nand2_1 U10939 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Kg9vx4 ), .op(n9059) );
  nand2_1 U10940 ( .ip1(n10206), .ip2(n9059), .op(n9069) );
  nand2_1 U10941 ( .ip1(n12558), .ip2(n10619), .op(n9071) );
  nand2_1 U10942 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n10206), .op(
        n9081) );
  nand2_1 U10943 ( .ip1(n11782), .ip2(n9081), .op(n9060) );
  nand2_1 U10944 ( .ip1(n9071), .ip2(n9060), .op(n9062) );
  nand2_1 U10945 ( .ip1(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip2(n9082), .op(
        n9061) );
  nand4_1 U10946 ( .ip1(n9086), .ip2(n9069), .ip3(n9062), .ip4(n9061), .op(
        n9097) );
  nor2_1 U10947 ( .ip1(n9063), .ip2(n9097), .op(n9064) );
  or2_1 U10948 ( .ip1(n3393), .ip2(n9064), .op(n9067) );
  or2_1 U10949 ( .ip1(n9065), .ip2(n9064), .op(n9066) );
  nand2_1 U10950 ( .ip1(n9067), .ip2(n9066), .op(
        \CORTEXM0DS_INST/u_logic/Jxhvx4 ) );
  nand2_1 U10951 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n9834), .op(
        n9070) );
  or2_1 U10952 ( .ip1(n9948), .ip2(n10206), .op(n9068) );
  nand4_1 U10953 ( .ip1(n11782), .ip2(n9070), .ip3(n9069), .ip4(n9068), .op(
        n9094) );
  nor2_1 U10954 ( .ip1(n12558), .ip2(n9094), .op(n9077) );
  nand2_1 U10955 ( .ip1(n9072), .ip2(n9071), .op(n9089) );
  inv_1 U10956 ( .ip(n9089), .op(n9095) );
  nor2_1 U10957 ( .ip1(n9095), .ip2(n12542), .op(n9076) );
  nand2_1 U10958 ( .ip1(n9948), .ip2(n11100), .op(n9074) );
  nand2_1 U10959 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(n10492), .op(
        n9073) );
  nand3_1 U10960 ( .ip1(n9074), .ip2(n11782), .ip3(n9073), .op(n9096) );
  nor2_1 U10961 ( .ip1(n11190), .ip2(n9096), .op(n9075) );
  nor4_1 U10962 ( .ip1(n9077), .ip2(n9076), .ip3(n9075), .ip4(n9097), .op(
        n9078) );
  or2_1 U10963 ( .ip1(n3393), .ip2(n9078), .op(n9080) );
  or2_1 U10964 ( .ip1(n11207), .ip2(n9078), .op(n9079) );
  nand2_1 U10965 ( .ip1(n9080), .ip2(n9079), .op(
        \CORTEXM0DS_INST/u_logic/Awhvx4 ) );
  nor2_1 U10966 ( .ip1(n9881), .ip2(n9094), .op(n9088) );
  inv_1 U10967 ( .ip(n9081), .op(n10734) );
  nand2_1 U10968 ( .ip1(n10734), .ip2(n11782), .op(n9085) );
  or2_1 U10969 ( .ip1(n12583), .ip2(n9096), .op(n9084) );
  nand4_1 U10970 ( .ip1(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip2(n9082), .ip3(
        n11782), .ip4(n12592), .op(n9083) );
  nand4_1 U10971 ( .ip1(n9086), .ip2(n9085), .ip3(n9084), .ip4(n9083), .op(
        n9087) );
  not_ab_or_c_or_d U10972 ( .ip1(\CORTEXM0DS_INST/u_logic/B19vx4 ), .ip2(n9089), .ip3(n9088), .ip4(n9087), .op(n9090) );
  or2_1 U10973 ( .ip1(n3393), .ip2(n9090), .op(n9093) );
  or2_1 U10974 ( .ip1(n9091), .ip2(n9090), .op(n9092) );
  nand2_1 U10975 ( .ip1(n9093), .ip2(n9092), .op(
        \CORTEXM0DS_INST/u_logic/Pthvx4 ) );
  nor2_1 U10976 ( .ip1(n12562), .ip2(n9094), .op(n9100) );
  inv_1 U10977 ( .ip(\CORTEXM0DS_INST/u_logic/I29vx4 ), .op(n12552) );
  nor2_1 U10978 ( .ip1(n9095), .ip2(n12552), .op(n9099) );
  nor2_1 U10979 ( .ip1(n12588), .ip2(n9096), .op(n9098) );
  nor4_1 U10980 ( .ip1(n9100), .ip2(n9099), .ip3(n9098), .ip4(n9097), .op(
        n9101) );
  or2_1 U10981 ( .ip1(n3393), .ip2(n9101), .op(n9104) );
  or2_1 U10982 ( .ip1(n9102), .ip2(n9101), .op(n9103) );
  nand2_1 U10983 ( .ip1(n9104), .ip2(n9103), .op(
        \CORTEXM0DS_INST/u_logic/Rghvx4 ) );
  inv_1 U10984 ( .ip(n9106), .op(n12062) );
  nand2_1 U10985 ( .ip1(n12062), .ip2(n11029), .op(n4806) );
  nor2_1 U10986 ( .ip1(\CORTEXM0DS_INST/u_logic/R9fvx4 ), .ip2(n4806), .op(
        n9107) );
  or2_1 U10987 ( .ip1(n9105), .ip2(n9107), .op(n9109) );
  nor2_1 U10988 ( .ip1(n11029), .ip2(n9106), .op(n12519) );
  or2_1 U10989 ( .ip1(n12519), .ip2(n9107), .op(n9108) );
  nand2_1 U10990 ( .ip1(n9109), .ip2(n9108), .op(
        \CORTEXM0DS_INST/u_logic/Slnvx4 ) );
  inv_1 U10991 ( .ip(n11903), .op(n12688) );
  nor3_1 U10992 ( .ip1(n12688), .ip2(n9921), .ip3(n12687), .op(n2792) );
  nand2_1 U10993 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(n12685), .op(
        n6161) );
  inv_1 U10994 ( .ip(n2792), .op(n9111) );
  nor2_1 U10995 ( .ip1(n11705), .ip2(n6161), .op(n9110) );
  not_ab_or_c_or_d U10996 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [7]), .ip2(
        n9111), .ip3(n12748), .ip4(n9110), .op(n9112) );
  or2_1 U10997 ( .ip1(n3276), .ip2(n9112), .op(n9115) );
  or2_1 U10998 ( .ip1(n9113), .ip2(n9112), .op(n9114) );
  nand2_1 U10999 ( .ip1(n9115), .ip2(n9114), .op(
        \CORTEXM0DS_INST/u_logic/W0ivx4 ) );
  nand2_1 U11000 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(n12671), .op(
        n6166) );
  nor2_1 U11001 ( .ip1(n11705), .ip2(n6166), .op(n9116) );
  or2_1 U11002 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [2]), .ip2(n9116), .op(
        n9117) );
  nand2_1 U11003 ( .ip1(n2620), .ip2(n9117), .op(n9118) );
  or2_1 U11004 ( .ip1(n3276), .ip2(n9118), .op(n9121) );
  or2_1 U11005 ( .ip1(n9119), .ip2(n9118), .op(n9120) );
  nand2_1 U11006 ( .ip1(n9121), .ip2(n9120), .op(
        \CORTEXM0DS_INST/u_logic/F2ivx4 ) );
  inv_1 U11007 ( .ip(n12681), .op(n10077) );
  mux2_1 U11008 ( .ip1(n11340), .ip2(n10077), .s(n12664), .op(
        \CORTEXM0DS_INST/u_logic/Bq5wx4 ) );
  nor2_1 U11009 ( .ip1(\CORTEXM0DS_INST/u_logic/Bq5wx4 ), .ip2(n11705), .op(
        n9122) );
  or2_1 U11010 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [14]), .ip2(n9122), .op(
        n9123) );
  nand2_1 U11011 ( .ip1(n9123), .ip2(n2754), .op(n9124) );
  or2_1 U11012 ( .ip1(n3276), .ip2(n9124), .op(n9127) );
  or2_1 U11013 ( .ip1(n9125), .ip2(n9124), .op(n9126) );
  nand2_1 U11014 ( .ip1(n9127), .ip2(n9126), .op(
        \CORTEXM0DS_INST/u_logic/Zyhvx4 ) );
  inv_1 U11015 ( .ip(n11807), .op(n12673) );
  nand2_1 U11016 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(n12673), .op(
        n6184) );
  nor2_1 U11017 ( .ip1(n11705), .ip2(n6184), .op(n9128) );
  or2_1 U11018 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [1]), .ip2(n9128), .op(
        n9129) );
  nand2_1 U11019 ( .ip1(n9129), .ip2(n2776), .op(n9130) );
  or2_1 U11020 ( .ip1(n3276), .ip2(n9130), .op(n9133) );
  or2_1 U11021 ( .ip1(n9131), .ip2(n9130), .op(n9132) );
  nand2_1 U11022 ( .ip1(n9133), .ip2(n9132), .op(
        \CORTEXM0DS_INST/u_logic/M2ivx4 ) );
  inv_1 U11023 ( .ip(n9134), .op(n12686) );
  nor2_1 U11024 ( .ip1(n9921), .ip2(n12686), .op(n11851) );
  or2_1 U11025 ( .ip1(n11851), .ip2(\CORTEXM0DS_INST/u_logic/Eqgvx4 ), .op(
        n9136) );
  inv_1 U11026 ( .ip(n3227), .op(n12644) );
  or2_1 U11027 ( .ip1(n12644), .ip2(\CORTEXM0DS_INST/u_logic/Eqgvx4 ), .op(
        n9135) );
  nand2_1 U11028 ( .ip1(n9136), .ip2(n9135), .op(n9137) );
  or2_1 U11029 ( .ip1(n3276), .ip2(n9137), .op(n9139) );
  or2_1 U11030 ( .ip1(n12410), .ip2(n9137), .op(n9138) );
  nand2_1 U11031 ( .ip1(n9139), .ip2(n9138), .op(
        \CORTEXM0DS_INST/u_logic/Owgvx4 ) );
  or2_1 U11032 ( .ip1(n12343), .ip2(n10041), .op(n9141) );
  nand2_1 U11033 ( .ip1(n9141), .ip2(n9140), .op(
        \CORTEXM0DS_INST/u_logic/N4421 ) );
  inv_1 U11034 ( .ip(\interconnect_ip_inst/i_ahb_U_mux_hsel_prev [1]), .op(
        n5920) );
  or2_1 U11035 ( .ip1(n5920), .ip2(n5919), .op(n9145) );
  nor2_1 U11036 ( .ip1(\interconnect_ip_inst/i_ahb_U_dfltslv_current_state ), 
        .ip2(\interconnect_ip_inst/i_ahb_U_mux_hsel_prev [2]), .op(n9142) );
  not_ab_or_c_or_d U11037 ( .ip1(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [2]), .ip2(
        \interconnect_ip_inst/i_apb_hready_resp ), .ip3(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [3]), .ip4(n9142), .op(
        n9143) );
  or2_1 U11038 ( .ip1(\interconnect_ip_inst/i_ahb_U_mux_hsel_prev [4]), .ip2(
        n9143), .op(n9987) );
  or2_1 U11039 ( .ip1(n9987), .ip2(n5919), .op(n9144) );
  nand2_1 U11040 ( .ip1(n9145), .ip2(n9144), .op(\interconnect_ip_inst/n4861 )
         );
  nand4_1 U11041 ( .ip1(n11902), .ip2(n9146), .ip3(n11901), .ip4(n12433), .op(
        n11817) );
  nor3_1 U11042 ( .ip1(n11871), .ip2(n9986), .ip3(n11817), .op(n12690) );
  nor2_1 U11044 ( .ip1(n9147), .ip2(n9156), .op(n9154) );
  nor2_1 U11045 ( .ip1(n9148), .ip2(n9243), .op(n9153) );
  nor2_1 U11046 ( .ip1(n9149), .ip2(n9158), .op(n9152) );
  nor2_1 U11047 ( .ip1(n9150), .ip2(n9160), .op(n9151) );
  nor4_1 U11048 ( .ip1(n9154), .ip2(n9153), .ip3(n9152), .ip4(n9151), .op(
        n9171) );
  and2_1 U11049 ( .ip1(n9155), .ip2(n9181), .op(n9165) );
  nor2_1 U11050 ( .ip1(n9157), .ip2(n9156), .op(n9164) );
  nor2_1 U11051 ( .ip1(n9159), .ip2(n9158), .op(n9163) );
  nor2_1 U11052 ( .ip1(n9161), .ip2(n9160), .op(n9162) );
  nor4_1 U11053 ( .ip1(n9165), .ip2(n9164), .ip3(n9163), .ip4(n9162), .op(
        n10088) );
  mux2_1 U11054 ( .ip1(n9171), .ip2(n10088), .s(n10256), .op(n11661) );
  nand2_1 U11055 ( .ip1(n9166), .ip2(n10255), .op(n9195) );
  inv_1 U11056 ( .ip(n9195), .op(n9169) );
  nor2_1 U11057 ( .ip1(n10256), .ip2(n9167), .op(n10142) );
  nand3_1 U11058 ( .ip1(n9169), .ip2(n9168), .ip3(n10142), .op(n9174) );
  nor2_1 U11059 ( .ip1(n9170), .ip2(n10263), .op(n9216) );
  and2_1 U11060 ( .ip1(n10256), .ip2(n9171), .op(n10141) );
  nand3_1 U11061 ( .ip1(n9225), .ip2(n9216), .ip3(n10141), .op(n9173) );
  not_ab_or_c_or_d U11062 ( .ip1(n9174), .ip2(n9173), .ip3(n9172), .ip4(n10269), .op(n9175) );
  nand3_1 U11063 ( .ip1(n11661), .ip2(n9175), .ip3(n9669), .op(n9177) );
  nand2_1 U11064 ( .ip1(n9177), .ip2(n9176), .op(n9206) );
  nand2_1 U11065 ( .ip1(n9179), .ip2(n9178), .op(n9189) );
  nand2_1 U11066 ( .ip1(n9181), .ip2(n9180), .op(n9188) );
  nand2_1 U11067 ( .ip1(n9183), .ip2(n9182), .op(n9187) );
  nand2_1 U11068 ( .ip1(n9185), .ip2(n9184), .op(n9186) );
  nand4_1 U11069 ( .ip1(n9189), .ip2(n9188), .ip3(n9187), .ip4(n9186), .op(
        n11646) );
  mux2_1 U11070 ( .ip1(n9190), .ip2(n11646), .s(n10256), .op(n11832) );
  nor4_1 U11071 ( .ip1(n9681), .ip2(n11832), .ip3(n9191), .ip4(n10253), .op(
        n9200) );
  inv_1 U11072 ( .ip(n9192), .op(n9194) );
  nor4_1 U11073 ( .ip1(n11646), .ip2(n10098), .ip3(n9194), .ip4(n9193), .op(
        n9198) );
  nor3_1 U11074 ( .ip1(n10097), .ip2(n9196), .ip3(n9195), .op(n9197) );
  mux2_1 U11075 ( .ip1(n9198), .ip2(n9197), .s(n10256), .op(n9199) );
  nand2_1 U11076 ( .ip1(n9200), .ip2(n9199), .op(n9204) );
  nand2_1 U11077 ( .ip1(n9202), .ip2(n9201), .op(n9203) );
  nand2_1 U11078 ( .ip1(n9204), .ip2(n9203), .op(n9205) );
  nand2_1 U11079 ( .ip1(n9206), .ip2(n9205), .op(n9210) );
  and2_1 U11080 ( .ip1(n9208), .ip2(n9207), .op(n9209) );
  nand2_1 U11081 ( .ip1(n9210), .ip2(n9209), .op(n9260) );
  nor2_1 U11082 ( .ip1(n9211), .ip2(n9213), .op(n9212) );
  not_ab_or_c_or_d U11083 ( .ip1(n9214), .ip2(n9213), .ip3(n9251), .ip4(n9212), 
        .op(n9258) );
  nand3_1 U11084 ( .ip1(n10088), .ip2(n9216), .ip3(n9215), .op(n9222) );
  nand4_1 U11085 ( .ip1(n9219), .ip2(n9218), .ip3(n10086), .ip4(n9217), .op(
        n9221) );
  not_ab_or_c_or_d U11086 ( .ip1(n9222), .ip2(n9221), .ip3(n9220), .ip4(n10277), .op(n9226) );
  inv_1 U11087 ( .ip(n9223), .op(n9224) );
  mux2_1 U11088 ( .ip1(n9225), .ip2(n9224), .s(n10256), .op(n9671) );
  nand3_1 U11089 ( .ip1(n9226), .ip2(n9671), .ip3(n9680), .op(n9257) );
  nor2_1 U11090 ( .ip1(n9227), .ip2(n10256), .op(n9231) );
  mux2_1 U11091 ( .ip1(n9230), .ip2(n9229), .s(n9228), .op(n10247) );
  not_ab_or_c_or_d U11092 ( .ip1(n10256), .ip2(n9232), .ip3(n9231), .ip4(
        n10247), .op(n10249) );
  inv_1 U11093 ( .ip(n9233), .op(n9235) );
  mux2_1 U11094 ( .ip1(n9235), .ip2(n9234), .s(n10256), .op(n9236) );
  mux2_1 U11095 ( .ip1(n9247), .ip2(n9236), .s(n9245), .op(n10083) );
  nor4_1 U11096 ( .ip1(n9238), .ip2(n9237), .ip3(n10249), .ip4(n10083), .op(
        n9239) );
  or2_1 U11097 ( .ip1(n9239), .ip2(n9251), .op(n9254) );
  inv_1 U11098 ( .ip(n9240), .op(n9241) );
  mux2_1 U11099 ( .ip1(n9242), .ip2(n9241), .s(n10256), .op(n9677) );
  mux2_1 U11100 ( .ip1(n9245), .ip2(n9244), .s(n9243), .op(n9246) );
  mux2_1 U11101 ( .ip1(n9247), .ip2(n9677), .s(n9246), .op(n11840) );
  nor4_1 U11102 ( .ip1(n9250), .ip2(n11840), .ip3(n9249), .ip4(n9248), .op(
        n9252) );
  or2_1 U11103 ( .ip1(n9252), .ip2(n9251), .op(n9253) );
  nand2_1 U11104 ( .ip1(n9254), .ip2(n9253), .op(n9255) );
  not_ab_or_c_or_d U11105 ( .ip1(n9258), .ip2(n9257), .ip3(n9256), .ip4(n9255), 
        .op(n9259) );
  nand2_1 U11106 ( .ip1(n9260), .ip2(n9259), .op(n9654) );
  nor2_1 U11107 ( .ip1(n9525), .ip2(n10040), .op(n9530) );
  and2_1 U11108 ( .ip1(n9261), .ip2(n9530), .op(n9265) );
  nor2_1 U11109 ( .ip1(n9263), .ip2(n9262), .op(n9264) );
  nor2_1 U11110 ( .ip1(n9265), .ip2(n9264), .op(n9305) );
  nand2_1 U11111 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [30]), .op(n9268) );
  nand2_1 U11112 ( .ip1(n9338), .ip2(\CORTEXM0DS_INST/cm0_r00 [30]), .op(n9267) );
  nand2_1 U11113 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [30]), .op(n9266) );
  nand3_1 U11114 ( .ip1(n9268), .ip2(n9267), .ip3(n9266), .op(n9286) );
  nand2_1 U11115 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [30]), .ip2(n9310), .op(n9284) );
  nand2_1 U11116 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [30]), .op(n9272) );
  nand2_1 U11117 ( .ip1(n9314), .ip2(\CORTEXM0DS_INST/cm0_r06 [30]), .op(n9271) );
  nand2_1 U11118 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [30]), .op(n9270) );
  nand2_1 U11119 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [30]), .op(n9269) );
  nand2_1 U11120 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [28]), .op(n9276) );
  nand2_1 U11121 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [28]), .op(n9275) );
  nand2_1 U11122 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [30]), .op(n9274) );
  nand2_1 U11123 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [30]), .op(n9273) );
  not_ab_or_c_or_d U11124 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [30]), 
        .ip3(n9278), .ip4(n9277), .op(n9283) );
  inv_1 U11125 ( .ip(\CORTEXM0DS_INST/u_logic/S4evx4 ), .op(n9350) );
  nor2_1 U11126 ( .ip1(n9279), .ip2(n9350), .op(n9281) );
  and2_1 U11127 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [30]), .op(n9280)
         );
  not_ab_or_c_or_d U11128 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [30]), .ip2(n9309), 
        .ip3(n9281), .ip4(n9280), .op(n9282) );
  nand3_1 U11129 ( .ip1(n9284), .ip2(n9283), .ip3(n9282), .op(n9285) );
  not_ab_or_c_or_d U11130 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [30]), 
        .ip3(n9286), .ip4(n9285), .op(n11671) );
  mux2_1 U11131 ( .ip1(n9346), .ip2(n9345), .s(n11671), .op(n9622) );
  and2_1 U11132 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [30]), .op(n9296)
         );
  nor2_1 U11133 ( .ip1(n9287), .ip2(n9348), .op(n9290) );
  nor2_1 U11134 ( .ip1(n12088), .ip2(n9288), .op(n9289) );
  not_ab_or_c_or_d U11135 ( .ip1(\CORTEXM0DS_INST/vis_psp [28]), .ip2(n9356), 
        .ip3(n9290), .ip4(n9289), .op(n9294) );
  nand2_1 U11136 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [30]), .op(n9293) );
  nand2_1 U11137 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [30]), .op(n9292) );
  nand2_1 U11138 ( .ip1(n9353), .ip2(\CORTEXM0DS_INST/u_logic/S4evx4 ), .op(
        n9291) );
  not_ab_or_c_or_d U11139 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [30]), .ip2(n9364), 
        .ip3(n9296), .ip4(n9295), .op(n9300) );
  nand2_1 U11140 ( .ip1(n9363), .ip2(\CORTEXM0DS_INST/cm0_r11 [30]), .op(n9299) );
  nand2_1 U11141 ( .ip1(n9347), .ip2(\CORTEXM0DS_INST/cm0_r14 [30]), .op(n9298) );
  nand2_1 U11142 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [28]), .op(n9297) );
  nand2_1 U11143 ( .ip1(n9471), .ip2(n9261), .op(n9301) );
  xor2_1 U11144 ( .ip1(n9622), .ip2(n9301), .op(n9304) );
  xor2_1 U11145 ( .ip1(n9305), .ip2(n9304), .op(n9646) );
  and2_1 U11146 ( .ip1(n9303), .ip2(n9302), .op(n9645) );
  nand2_1 U11147 ( .ip1(n9646), .ip2(n9645), .op(n9718) );
  nand2_1 U11148 ( .ip1(n9622), .ip2(n9471), .op(n11500) );
  nor2_1 U11149 ( .ip1(n9371), .ip2(n11500), .op(n9307) );
  nor2_1 U11150 ( .ip1(n9305), .ip2(n9304), .op(n9306) );
  nor2_1 U11151 ( .ip1(n9307), .ip2(n9306), .op(n9716) );
  nand2_1 U11152 ( .ip1(n9308), .ip2(\CORTEXM0DS_INST/cm0_r01 [31]), .op(n9313) );
  nand2_1 U11153 ( .ip1(n9309), .ip2(\CORTEXM0DS_INST/cm0_r09 [31]), .op(n9312) );
  nand2_1 U11154 ( .ip1(n9310), .ip2(\CORTEXM0DS_INST/cm0_r05 [31]), .op(n9311) );
  nand3_1 U11155 ( .ip1(n9313), .ip2(n9312), .ip3(n9311), .op(n9343) );
  nand2_1 U11156 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [31]), .ip2(n9314), .op(n9341) );
  nand2_1 U11157 ( .ip1(n9315), .ip2(\CORTEXM0DS_INST/cm0_r07 [31]), .op(n9322) );
  nand2_1 U11158 ( .ip1(n9316), .ip2(\CORTEXM0DS_INST/cm0_r02 [31]), .op(n9321) );
  nand2_1 U11159 ( .ip1(n9317), .ip2(\CORTEXM0DS_INST/cm0_r12 [31]), .op(n9320) );
  nand2_1 U11160 ( .ip1(n9318), .ip2(\CORTEXM0DS_INST/cm0_r04 [31]), .op(n9319) );
  nand2_1 U11161 ( .ip1(n9323), .ip2(\CORTEXM0DS_INST/vis_psp [29]), .op(n9330) );
  nand2_1 U11162 ( .ip1(n9324), .ip2(\CORTEXM0DS_INST/cm0_r14 [31]), .op(n9329) );
  nand2_1 U11163 ( .ip1(n9325), .ip2(\CORTEXM0DS_INST/u_logic/D6evx4 ), .op(
        n9328) );
  nand2_1 U11164 ( .ip1(n9326), .ip2(\CORTEXM0DS_INST/cm0_r11 [31]), .op(n9327) );
  not_ab_or_c_or_d U11165 ( .ip1(n9333), .ip2(\CORTEXM0DS_INST/vis_msp [29]), 
        .ip3(n9332), .ip4(n9331), .op(n9340) );
  and2_1 U11166 ( .ip1(n9334), .ip2(\CORTEXM0DS_INST/cm0_r08 [31]), .op(n9337)
         );
  and2_1 U11167 ( .ip1(n9335), .ip2(\CORTEXM0DS_INST/cm0_r10 [31]), .op(n9336)
         );
  not_ab_or_c_or_d U11168 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [31]), .ip2(n9338), 
        .ip3(n9337), .ip4(n9336), .op(n9339) );
  nand3_1 U11169 ( .ip1(n9341), .ip2(n9340), .ip3(n9339), .op(n9342) );
  not_ab_or_c_or_d U11170 ( .ip1(n9344), .ip2(\CORTEXM0DS_INST/cm0_r03 [31]), 
        .ip3(n9343), .ip4(n9342), .op(n10072) );
  mux2_1 U11171 ( .ip1(n9346), .ip2(n9345), .s(n10072), .op(n9394) );
  and2_1 U11172 ( .ip1(n9347), .ip2(\CORTEXM0DS_INST/cm0_r14 [31]), .op(n9362)
         );
  nor2_1 U11173 ( .ip1(n9349), .ip2(n9348), .op(n9352) );
  nor2_1 U11174 ( .ip1(n12088), .ip2(n9350), .op(n9351) );
  not_ab_or_c_or_d U11175 ( .ip1(\CORTEXM0DS_INST/u_logic/D6evx4 ), .ip2(n9353), .ip3(n9352), .ip4(n9351), .op(n9360) );
  nand2_1 U11176 ( .ip1(n9354), .ip2(\CORTEXM0DS_INST/cm0_r08 [31]), .op(n9359) );
  nand2_1 U11177 ( .ip1(n9355), .ip2(\CORTEXM0DS_INST/cm0_r10 [31]), .op(n9358) );
  nand2_1 U11178 ( .ip1(n9356), .ip2(\CORTEXM0DS_INST/vis_psp [29]), .op(n9357) );
  not_ab_or_c_or_d U11179 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [31]), .ip2(n9363), 
        .ip3(n9362), .ip4(n9361), .op(n9370) );
  nand2_1 U11180 ( .ip1(n9364), .ip2(\CORTEXM0DS_INST/cm0_r09 [31]), .op(n9369) );
  nand2_1 U11181 ( .ip1(n9365), .ip2(\CORTEXM0DS_INST/cm0_r12 [31]), .op(n9368) );
  nand2_1 U11182 ( .ip1(n9366), .ip2(\CORTEXM0DS_INST/vis_msp [29]), .op(n9367) );
  nand2_1 U11183 ( .ip1(n9394), .ip2(n9990), .op(n9381) );
  nor2_1 U11184 ( .ip1(n9371), .ip2(n9381), .op(n9750) );
  or2_1 U11185 ( .ip1(n9261), .ip2(n9394), .op(n9373) );
  or2_1 U11186 ( .ip1(n9990), .ip2(n9394), .op(n9372) );
  nand2_1 U11187 ( .ip1(n9373), .ip2(n9372), .op(n9749) );
  nor2_1 U11188 ( .ip1(n9750), .ip2(n9749), .op(n9714) );
  xor2_1 U11189 ( .ip1(n9716), .ip2(n9714), .op(n9717) );
  xor2_1 U11190 ( .ip1(n9718), .ip2(n9717), .op(n10462) );
  not_ab_or_c_or_d U11191 ( .ip1(n12133), .ip2(n11796), .ip3(n10611), .ip4(
        n9374), .op(n9375) );
  mux2_1 U11192 ( .ip1(n9375), .ip2(n11016), .s(
        \CORTEXM0DS_INST/u_logic/Vdgvx4 ), .op(n9376) );
  nand2_1 U11193 ( .ip1(n9377), .ip2(n9376), .op(n9378) );
  nand2_1 U11194 ( .ip1(n9378), .ip2(\CORTEXM0DS_INST/u_logic/O8gvx4 ), .op(
        n9380) );
  nand2_1 U11195 ( .ip1(n9380), .ip2(n9379), .op(n11578) );
  inv_1 U11196 ( .ip(n9381), .op(n9397) );
  nor3_1 U11197 ( .ip1(n9797), .ip2(n9382), .ip3(n11239), .op(n11558) );
  nand2_1 U11198 ( .ip1(n9394), .ip2(n11558), .op(n9384) );
  inv_1 U11199 ( .ip(n9990), .op(n9383) );
  nand2_1 U11200 ( .ip1(n9384), .ip2(n9383), .op(n9396) );
  nand2_1 U11201 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(n9817) );
  nor2_1 U11202 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n9817), .op(
        n10805) );
  not_ab_or_c_or_d U11203 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(
        n11683), .ip3(n12125), .ip4(n10851), .op(n9386) );
  not_ab_or_c_or_d U11204 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        n10805), .ip3(n9386), .ip4(n9385), .op(n9387) );
  or2_1 U11205 ( .ip1(n9387), .ip2(n9797), .op(n9391) );
  nand3_1 U11206 ( .ip1(n9388), .ip2(n12623), .ip3(n11786), .op(n9389) );
  or2_1 U11207 ( .ip1(n9389), .ip2(n9797), .op(n9390) );
  nand2_1 U11208 ( .ip1(n9391), .ip2(n9390), .op(n9392) );
  or2_1 U11209 ( .ip1(n9393), .ip2(n9392), .op(n9445) );
  nor2_1 U11210 ( .ip1(n9445), .ip2(n11558), .op(n11564) );
  inv_1 U11211 ( .ip(n11564), .op(n11583) );
  or2_1 U11212 ( .ip1(n11583), .ip2(n9394), .op(n9395) );
  nand2_1 U11213 ( .ip1(n9396), .ip2(n9395), .op(n9399) );
  or2_1 U11214 ( .ip1(n9397), .ip2(n9399), .op(n9401) );
  nor2_1 U11215 ( .ip1(n11209), .ip2(n12369), .op(n9398) );
  not_ab_or_c_or_d U11216 ( .ip1(n11796), .ip2(n11786), .ip3(
        \CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip4(n9398), .op(n9446) );
  or2_1 U11217 ( .ip1(n9446), .ip2(n9445), .op(n11588) );
  inv_1 U11218 ( .ip(n11588), .op(n11501) );
  or2_1 U11219 ( .ip1(n11501), .ip2(n9399), .op(n9400) );
  nand2_1 U11220 ( .ip1(n9401), .ip2(n9400), .op(n9408) );
  inv_1 U11221 ( .ip(n10072), .op(n11667) );
  or2_1 U11222 ( .ip1(n9402), .ip2(n9797), .op(n9404) );
  or2_1 U11223 ( .ip1(n11277), .ip2(n9797), .op(n9403) );
  nand2_1 U11224 ( .ip1(n9404), .ip2(n9403), .op(n11594) );
  nand2_1 U11225 ( .ip1(n11667), .ip2(n11594), .op(n9406) );
  nor3_1 U11226 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n12117), .ip3(
        n11681), .op(n10650) );
  nand2_1 U11227 ( .ip1(\CORTEXM0DS_INST/u_logic/O8gvx4 ), .ip2(n10650), .op(
        n11522) );
  nor3_1 U11228 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip3(n11522), .op(n11496) );
  nand2_1 U11229 ( .ip1(n11496), .ip2(\CORTEXM0DS_INST/vis_apsr [3]), .op(
        n9405) );
  nand3_1 U11230 ( .ip1(\CORTEXM0DS_INST/u_logic/O8gvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip3(n11208), .op(n11438) );
  nand3_1 U11231 ( .ip1(n9406), .ip2(n9405), .ip3(n11438), .op(n9407) );
  not_ab_or_c_or_d U11232 ( .ip1(n10462), .ip2(n11578), .ip3(n9408), .ip4(
        n9407), .op(n11505) );
  nor2_1 U11233 ( .ip1(\CORTEXM0DS_INST/u_logic/Dw8vx4 ), .ip2(n11505), .op(
        n9743) );
  inv_1 U11234 ( .ip(n11578), .op(n9572) );
  nor2_1 U11235 ( .ip1(n9572), .ip2(n10232), .op(n11507) );
  xor2_1 U11236 ( .ip1(n9410), .ip2(n9409), .op(n12301) );
  nor2_1 U11237 ( .ip1(n9572), .ip2(n12301), .op(n11480) );
  xor2_1 U11238 ( .ip1(n9412), .ip2(n9411), .op(n12351) );
  xor2_1 U11239 ( .ip1(n9414), .ip2(n9413), .op(n12155) );
  nand4_1 U11240 ( .ip1(n12155), .ip2(n12282), .ip3(n11060), .ip4(n9415), .op(
        n9426) );
  xor2_1 U11241 ( .ip1(n9417), .ip2(n9416), .op(n11326) );
  inv_1 U11242 ( .ip(n11326), .op(n12198) );
  xor2_1 U11243 ( .ip1(n9419), .ip2(n9418), .op(n11337) );
  inv_1 U11244 ( .ip(n11337), .op(n10194) );
  nand3_1 U11245 ( .ip1(n12188), .ip2(n12198), .ip3(n10194), .op(n9425) );
  inv_1 U11246 ( .ip(n11357), .op(n12213) );
  xor2_1 U11247 ( .ip1(n9421), .ip2(n9420), .op(n11579) );
  inv_1 U11248 ( .ip(n11579), .op(n11007) );
  xor2_1 U11249 ( .ip1(n9423), .ip2(n9422), .op(n11347) );
  inv_1 U11250 ( .ip(n11347), .op(n10330) );
  nand3_1 U11251 ( .ip1(n12213), .ip2(n11007), .ip3(n10330), .op(n9424) );
  nor4_1 U11252 ( .ip1(n11437), .ip2(n9426), .ip3(n9425), .ip4(n9424), .op(
        n9433) );
  xor2_1 U11253 ( .ip1(n9428), .ip2(n9427), .op(n11401) );
  inv_1 U11254 ( .ip(n11401), .op(n12252) );
  xor2_1 U11255 ( .ip1(n9430), .ip2(n9429), .op(n12232) );
  xor2_1 U11256 ( .ip1(n9432), .ip2(n9431), .op(n11370) );
  inv_1 U11257 ( .ip(n11370), .op(n12222) );
  nand4_1 U11258 ( .ip1(n9433), .ip2(n12252), .ip3(n12232), .ip4(n12222), .op(
        n9434) );
  nor3_1 U11259 ( .ip1(n12351), .ip2(n9434), .ip3(n12276), .op(n9435) );
  nor2_1 U11260 ( .ip1(n9572), .ip2(n9435), .op(n9651) );
  xnor2_1 U11261 ( .ip1(n9437), .ip2(n9436), .op(n12312) );
  nor2_1 U11262 ( .ip1(n9572), .ip2(n12312), .op(n11483) );
  xor2_1 U11263 ( .ip1(n9439), .ip2(n9438), .op(n12291) );
  nor2_1 U11264 ( .ip1(n9572), .ip2(n12291), .op(n11466) );
  xor2_1 U11265 ( .ip1(n9441), .ip2(n9440), .op(n12263) );
  nor2_1 U11266 ( .ip1(n9572), .ip2(n12263), .op(n11415) );
  inv_1 U11267 ( .ip(n11438), .op(n11593) );
  or2_1 U11268 ( .ip1(n12169), .ip2(n11593), .op(n9443) );
  or2_1 U11269 ( .ip1(n11578), .ip2(n11593), .op(n9442) );
  nand2_1 U11270 ( .ip1(n9443), .ip2(n9442), .op(n11204) );
  inv_1 U11271 ( .ip(n11558), .op(n11581) );
  nor2_1 U11272 ( .ip1(n11581), .ip2(n9447), .op(n9444) );
  not_ab_or_c_or_d U11273 ( .ip1(n9446), .ip2(n9447), .ip3(n9445), .ip4(n9444), 
        .op(n9449) );
  nand2_1 U11274 ( .ip1(n11558), .ip2(n9447), .op(n9448) );
  mux2_1 U11275 ( .ip1(n9449), .ip2(n9448), .s(n12331), .op(n9452) );
  nand2_1 U11276 ( .ip1(n12339), .ip2(n11578), .op(n9451) );
  nand2_1 U11277 ( .ip1(n11594), .ip2(n12685), .op(n9450) );
  nand4_1 U11278 ( .ip1(n9452), .ip2(n11438), .ip3(n9451), .ip4(n9450), .op(
        n11514) );
  nand2_1 U11279 ( .ip1(n11558), .ip2(n9453), .op(n9457) );
  nor2_1 U11280 ( .ip1(n11583), .ip2(n9453), .op(n9456) );
  nand2_1 U11281 ( .ip1(n11501), .ip2(n9453), .op(n9454) );
  nor2_1 U11282 ( .ip1(n9454), .ip2(n11760), .op(n9455) );
  not_ab_or_c_or_d U11283 ( .ip1(n11760), .ip2(n9457), .ip3(n9456), .ip4(n9455), .op(n11301) );
  nand2_1 U11284 ( .ip1(n9463), .ip2(n11558), .op(n9459) );
  nand2_1 U11285 ( .ip1(n9459), .ip2(n9458), .op(n9461) );
  or2_1 U11286 ( .ip1(n11583), .ip2(n9463), .op(n9460) );
  nand2_1 U11287 ( .ip1(n9461), .ip2(n9460), .op(n9465) );
  and3_1 U11288 ( .ip1(n9463), .ip2(n11501), .ip3(n9462), .op(n9464) );
  nor2_1 U11289 ( .ip1(n9465), .ip2(n9464), .op(n11445) );
  nand2_1 U11290 ( .ip1(n11558), .ip2(n9466), .op(n9470) );
  nor2_1 U11291 ( .ip1(n11583), .ip2(n9466), .op(n9469) );
  nand2_1 U11292 ( .ip1(n11501), .ip2(n9466), .op(n9467) );
  nor2_1 U11293 ( .ip1(n9467), .ip2(n12166), .op(n9468) );
  not_ab_or_c_or_d U11294 ( .ip1(n12166), .ip2(n9470), .ip3(n9469), .ip4(n9468), .op(n11202) );
  nor3_1 U11295 ( .ip1(n11301), .ip2(n11445), .ip3(n11202), .op(n9512) );
  and2_1 U11296 ( .ip1(n9597), .ip2(n12273), .op(n11418) );
  and2_1 U11297 ( .ip1(n9620), .ip2(n9621), .op(n11343) );
  not_ab_or_c_or_d U11298 ( .ip1(n9557), .ip2(n11362), .ip3(n11418), .ip4(
        n11343), .op(n9480) );
  nand2_1 U11299 ( .ip1(n9617), .ip2(n9616), .op(n11331) );
  nand2_1 U11300 ( .ip1(n9590), .ip2(n9591), .op(n11396) );
  nand2_1 U11301 ( .ip1(n9595), .ip2(n9596), .op(n11350) );
  nand3_1 U11302 ( .ip1(n11331), .ip2(n11396), .ip3(n11350), .op(n9476) );
  and2_1 U11303 ( .ip1(n9618), .ip2(n9619), .op(n11308) );
  inv_1 U11304 ( .ip(n9594), .op(n9633) );
  nor2_1 U11305 ( .ip1(n9633), .ip2(n12235), .op(n11376) );
  not_ab_or_c_or_d U11306 ( .ip1(n11318), .ip2(n9592), .ip3(n11308), .ip4(
        n11376), .op(n9474) );
  inv_1 U11307 ( .ip(n9471), .op(n10029) );
  and2_1 U11308 ( .ip1(n9622), .ip2(n10029), .op(n11499) );
  nor2_1 U11309 ( .ip1(n11476), .ip2(n12304), .op(n9472) );
  not_ab_or_c_or_d U11310 ( .ip1(n9560), .ip2(n11559), .ip3(n11499), .ip4(
        n9472), .op(n9473) );
  nand2_1 U11311 ( .ip1(n9610), .ip2(n9611), .op(n11446) );
  nand2_1 U11312 ( .ip1(n12288), .ip2(n9542), .op(n11461) );
  nand4_1 U11313 ( .ip1(n9474), .ip2(n9473), .ip3(n11446), .ip4(n11461), .op(
        n9475) );
  not_ab_or_c_or_d U11314 ( .ip1(n11410), .ip2(n11405), .ip3(n9476), .ip4(
        n9475), .op(n9479) );
  nand2_1 U11315 ( .ip1(n11004), .ip2(n9593), .op(n9478) );
  nand2_1 U11316 ( .ip1(n12239), .ip2(n11385), .op(n9477) );
  nand4_1 U11317 ( .ip1(n9480), .ip2(n9479), .ip3(n9478), .ip4(n9477), .op(
        n9496) );
  nand2_1 U11318 ( .ip1(n11558), .ip2(n9481), .op(n9485) );
  nor2_1 U11319 ( .ip1(n11583), .ip2(n9481), .op(n9484) );
  nand2_1 U11320 ( .ip1(n11501), .ip2(n9481), .op(n9482) );
  nor2_1 U11321 ( .ip1(n9482), .ip2(n9486), .op(n9483) );
  not_ab_or_c_or_d U11322 ( .ip1(n9486), .ip2(n9485), .ip3(n9484), .ip4(n9483), 
        .op(n11431) );
  nand2_1 U11323 ( .ip1(n9489), .ip2(n11558), .op(n9488) );
  nand2_1 U11324 ( .ip1(n9488), .ip2(n9487), .op(n9491) );
  or2_1 U11325 ( .ip1(n11583), .ip2(n9489), .op(n9490) );
  nand2_1 U11326 ( .ip1(n9491), .ip2(n9490), .op(n9492) );
  or2_1 U11327 ( .ip1(n11501), .ip2(n9492), .op(n9495) );
  or2_1 U11328 ( .ip1(n9493), .ip2(n9492), .op(n9494) );
  nand2_1 U11329 ( .ip1(n9495), .ip2(n9494), .op(n11527) );
  not_ab_or_c_or_d U11330 ( .ip1(n11558), .ip2(n9496), .ip3(n11431), .ip4(
        n11527), .op(n9511) );
  nand3_1 U11331 ( .ip1(n9498), .ip2(n11501), .ip3(n9497), .op(n9503) );
  nand2_1 U11332 ( .ip1(n9497), .ip2(n9498), .op(n9501) );
  nand2_1 U11333 ( .ip1(n9497), .ip2(n11558), .op(n9500) );
  nand2_1 U11334 ( .ip1(n11583), .ip2(n9498), .op(n9499) );
  nand3_1 U11335 ( .ip1(n9501), .ip2(n9500), .ip3(n9499), .op(n9502) );
  nand2_1 U11336 ( .ip1(n9503), .ip2(n9502), .op(n11303) );
  nand3_1 U11337 ( .ip1(n9505), .ip2(n11501), .ip3(n9504), .op(n9510) );
  nand2_1 U11338 ( .ip1(n9504), .ip2(n9505), .op(n9508) );
  nand2_1 U11339 ( .ip1(n9504), .ip2(n11558), .op(n9507) );
  nand2_1 U11340 ( .ip1(n11583), .ip2(n9505), .op(n9506) );
  nand3_1 U11341 ( .ip1(n9508), .ip2(n9507), .ip3(n9506), .op(n9509) );
  nand2_1 U11342 ( .ip1(n9510), .ip2(n9509), .op(n11533) );
  nand4_1 U11343 ( .ip1(n9512), .ip2(n9511), .ip3(n11303), .ip4(n11533), .op(
        n9638) );
  nand2_1 U11344 ( .ip1(n9513), .ip2(n11583), .op(n9515) );
  nand2_1 U11345 ( .ip1(n9515), .ip2(n9514), .op(n9518) );
  nand2_1 U11346 ( .ip1(n11581), .ip2(n9516), .op(n9517) );
  nand2_1 U11347 ( .ip1(n9518), .ip2(n9517), .op(n9519) );
  or2_1 U11348 ( .ip1(n11501), .ip2(n9519), .op(n9522) );
  or2_1 U11349 ( .ip1(n9520), .ip2(n9519), .op(n9521) );
  nand2_1 U11350 ( .ip1(n9522), .ip2(n9521), .op(n9523) );
  not_ab_or_c_or_d U11351 ( .ip1(n11496), .ip2(\CORTEXM0DS_INST/vis_apsr [0]), 
        .ip3(n11593), .ip4(n9523), .op(n11512) );
  nand2_1 U11352 ( .ip1(n9524), .ip2(n11583), .op(n9526) );
  nand2_1 U11353 ( .ip1(n9526), .ip2(n9525), .op(n9528) );
  nand2_1 U11354 ( .ip1(n11581), .ip2(n10040), .op(n9527) );
  nand2_1 U11355 ( .ip1(n9528), .ip2(n9527), .op(n9529) );
  or2_1 U11356 ( .ip1(n11501), .ip2(n9529), .op(n9532) );
  or2_1 U11357 ( .ip1(n9530), .ip2(n9529), .op(n9531) );
  nand2_1 U11358 ( .ip1(n9532), .ip2(n9531), .op(n9533) );
  or2_1 U11359 ( .ip1(n11496), .ip2(n9533), .op(n9535) );
  or2_1 U11360 ( .ip1(\CORTEXM0DS_INST/vis_apsr [1]), .ip2(n9533), .op(n9534)
         );
  nand2_1 U11361 ( .ip1(n9535), .ip2(n9534), .op(n11493) );
  nand2_1 U11362 ( .ip1(n11558), .ip2(n9536), .op(n9540) );
  nor2_1 U11363 ( .ip1(n11583), .ip2(n9536), .op(n9539) );
  nand2_1 U11364 ( .ip1(n11501), .ip2(n9536), .op(n9537) );
  nor2_1 U11365 ( .ip1(n9537), .ip2(n12142), .op(n9538) );
  not_ab_or_c_or_d U11366 ( .ip1(n12142), .ip2(n9540), .ip3(n9539), .ip4(n9538), .op(n11574) );
  nor2_1 U11367 ( .ip1(n11583), .ip2(n9542), .op(n9541) );
  not_ab_or_c_or_d U11368 ( .ip1(n11501), .ip2(n9542), .ip3(n12288), .ip4(
        n9541), .op(n11465) );
  nor3_1 U11369 ( .ip1(n11564), .ip2(n9595), .ip3(n9596), .op(n11353) );
  nor3_1 U11370 ( .ip1(n11564), .ip2(n9590), .ip3(n9591), .op(n11400) );
  nor4_1 U11371 ( .ip1(n11574), .ip2(n11465), .ip3(n11353), .ip4(n11400), .op(
        n9549) );
  nor2_1 U11372 ( .ip1(n9546), .ip2(n11581), .op(n9545) );
  or2_1 U11373 ( .ip1(n9546), .ip2(n11588), .op(n9544) );
  inv_1 U11374 ( .ip(n9543), .op(n12315) );
  mux2_1 U11375 ( .ip1(n9545), .ip2(n9544), .s(n12315), .op(n9548) );
  nand2_1 U11376 ( .ip1(n9546), .ip2(n11564), .op(n9547) );
  nand2_1 U11377 ( .ip1(n9548), .ip2(n9547), .op(n11485) );
  nand4_1 U11378 ( .ip1(n11512), .ip2(n11493), .ip3(n9549), .ip4(n11485), .op(
        n9637) );
  nand3_1 U11379 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip3(
        \CORTEXM0DS_INST/cm0_control[1] ), .op(n9550) );
  or2_1 U11380 ( .ip1(n9550), .ip2(n11522), .op(n9553) );
  nand3_1 U11381 ( .ip1(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [1]), .ip3(n12104), .op(n9551) );
  or2_1 U11382 ( .ip1(n9551), .ip2(n11522), .op(n9552) );
  nand2_1 U11383 ( .ip1(n9553), .ip2(n9552), .op(n9554) );
  or2_1 U11384 ( .ip1(n10915), .ip2(n9554), .op(n9556) );
  or2_1 U11385 ( .ip1(n11578), .ip2(n9554), .op(n9555) );
  nand2_1 U11386 ( .ip1(n9556), .ip2(n9555), .op(n11535) );
  inv_1 U11387 ( .ip(n11362), .op(n11367) );
  inv_1 U11388 ( .ip(n9557), .op(n12225) );
  nor2_1 U11389 ( .ip1(n11318), .ip2(n9592), .op(n9559) );
  nor2_1 U11390 ( .ip1(n11004), .ip2(n9593), .op(n9558) );
  not_ab_or_c_or_d U11391 ( .ip1(n11367), .ip2(n12225), .ip3(n9559), .ip4(
        n9558), .op(n9564) );
  inv_1 U11392 ( .ip(n11559), .op(n11565) );
  inv_1 U11393 ( .ip(n9560), .op(n12158) );
  nand2_1 U11394 ( .ip1(n11565), .ip2(n12158), .op(n9563) );
  inv_1 U11395 ( .ip(n11385), .op(n11390) );
  inv_1 U11396 ( .ip(n12239), .op(n11384) );
  nand2_1 U11397 ( .ip1(n11390), .ip2(n11384), .op(n9562) );
  nand2_1 U11398 ( .ip1(n11476), .ip2(n12304), .op(n9561) );
  nand4_1 U11399 ( .ip1(n9564), .ip2(n9563), .ip3(n9562), .ip4(n9561), .op(
        n9565) );
  nor3_1 U11400 ( .ip1(n11564), .ip2(n12273), .ip3(n9597), .op(n11423) );
  nor3_1 U11401 ( .ip1(n11564), .ip2(n11410), .ip3(n11405), .op(n11406) );
  not_ab_or_c_or_d U11402 ( .ip1(n11583), .ip2(n9565), .ip3(n11423), .ip4(
        n11406), .op(n9635) );
  nand2_1 U11403 ( .ip1(n11558), .ip2(n9566), .op(n9570) );
  nor2_1 U11404 ( .ip1(n11583), .ip2(n9566), .op(n9569) );
  nand2_1 U11405 ( .ip1(n11501), .ip2(n9566), .op(n9567) );
  nor2_1 U11406 ( .ip1(n9567), .ip2(n9571), .op(n9568) );
  not_ab_or_c_or_d U11407 ( .ip1(n9571), .ip2(n9570), .ip3(n9569), .ip4(n9568), 
        .op(n11436) );
  nor2_1 U11408 ( .ip1(n9572), .ip2(n10384), .op(n11444) );
  nand4_1 U11409 ( .ip1(\CORTEXM0DS_INST/u_logic/O8gvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip3(n9573), .ip4(
        \CORTEXM0DS_INST/u_logic/Oy8vx4 ), .op(n9577) );
  nand2_1 U11410 ( .ip1(n11593), .ip2(\CORTEXM0DS_INST/cm0_control[1] ), .op(
        n9576) );
  nor3_1 U11411 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(n11517), .ip3(
        n11522), .op(n11427) );
  nand2_1 U11412 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [2]), .ip2(n11427), .op(
        n9575) );
  nand2_1 U11413 ( .ip1(n10418), .ip2(n11578), .op(n9574) );
  nand4_1 U11414 ( .ip1(n9577), .ip2(n9576), .ip3(n9575), .ip4(n9574), .op(
        n11299) );
  inv_1 U11415 ( .ip(n12662), .op(n9578) );
  nand4_1 U11416 ( .ip1(n10063), .ip2(n9578), .ip3(n11315), .ip4(n12665), .op(
        n9579) );
  nor3_1 U11417 ( .ip1(n11508), .ip2(n12661), .ip3(n9579), .op(n9588) );
  nand4_1 U11418 ( .ip1(n11819), .ip2(n11671), .ip3(n11462), .ip4(n11340), 
        .op(n9586) );
  inv_1 U11419 ( .ip(n9580), .op(n12678) );
  nor4_1 U11420 ( .ip1(n12682), .ip2(n12681), .ip3(n12678), .ip4(n12680), .op(
        n9581) );
  nand4_1 U11421 ( .ip1(n10058), .ip2(n11807), .ip3(n11455), .ip4(n9581), .op(
        n9585) );
  inv_1 U11422 ( .ip(n12671), .op(n11297) );
  nand4_1 U11423 ( .ip1(n11297), .ip2(n12670), .ip3(n11330), .ip4(n10071), 
        .op(n9584) );
  inv_1 U11424 ( .ip(n12677), .op(n9582) );
  nand4_1 U11425 ( .ip1(n12674), .ip2(n9582), .ip3(n12672), .ip4(n11382), .op(
        n9583) );
  nor4_1 U11426 ( .ip1(n9586), .ip2(n9585), .ip3(n9584), .ip4(n9583), .op(
        n9587) );
  nand4_1 U11427 ( .ip1(n10066), .ip2(n11477), .ip3(n9588), .ip4(n9587), .op(
        n9615) );
  nand2_1 U11428 ( .ip1(n11384), .ip2(n11385), .op(n11383) );
  nand2_1 U11429 ( .ip1(n12225), .ip2(n11362), .op(n11361) );
  nand4_1 U11430 ( .ip1(n11470), .ip2(n11500), .ip3(n11383), .ip4(n11361), 
        .op(n9602) );
  inv_1 U11431 ( .ip(n11410), .op(n12266) );
  nand2_1 U11432 ( .ip1(n12266), .ip2(n11405), .op(n9589) );
  nand2_1 U11433 ( .ip1(n10027), .ip2(n9620), .op(n11344) );
  nand2_1 U11434 ( .ip1(n12191), .ip2(n9618), .op(n11309) );
  nand2_1 U11435 ( .ip1(n12158), .ip2(n11559), .op(n11557) );
  nand4_1 U11436 ( .ip1(n9589), .ip2(n11344), .ip3(n11309), .ip4(n11557), .op(
        n9601) );
  inv_1 U11437 ( .ip(n9617), .op(n10022) );
  nand2_1 U11438 ( .ip1(n10022), .ip2(n9616), .op(n11334) );
  inv_1 U11439 ( .ip(n9590), .op(n12255) );
  nand2_1 U11440 ( .ip1(n12255), .ip2(n9591), .op(n11395) );
  inv_1 U11441 ( .ip(n9592), .op(n11316) );
  or2_1 U11442 ( .ip1(n11318), .ip2(n11316), .op(n11322) );
  inv_1 U11443 ( .ip(n9593), .op(n11580) );
  or2_1 U11444 ( .ip1(n11004), .ip2(n11580), .op(n11589) );
  nand4_1 U11445 ( .ip1(n11334), .ip2(n11395), .ip3(n11322), .ip4(n11589), 
        .op(n9600) );
  inv_1 U11446 ( .ip(n9610), .op(n12285) );
  nand2_1 U11447 ( .ip1(n12285), .ip2(n9611), .op(n11448) );
  nand2_1 U11448 ( .ip1(n12235), .ip2(n9594), .op(n11373) );
  inv_1 U11449 ( .ip(n9595), .op(n12216) );
  nand2_1 U11450 ( .ip1(n12216), .ip2(n9596), .op(n11351) );
  nand2_1 U11451 ( .ip1(n9598), .ip2(n9597), .op(n11421) );
  nand4_1 U11452 ( .ip1(n11448), .ip2(n11373), .ip3(n11351), .ip4(n11421), 
        .op(n9599) );
  nor4_1 U11453 ( .ip1(n9602), .ip2(n9601), .ip3(n9600), .ip4(n9599), .op(
        n9603) );
  nor2_1 U11454 ( .ip1(n11501), .ip2(n9603), .op(n9614) );
  inv_1 U11455 ( .ip(n11427), .op(n9606) );
  nor2_1 U11456 ( .ip1(n9606), .ip2(n9604), .op(n9605) );
  not_ab_or_c_or_d U11457 ( .ip1(n11594), .ip2(n12679), .ip3(n11593), .ip4(
        n9605), .op(n11441) );
  nor2_1 U11458 ( .ip1(n9606), .ip2(n11023), .op(n9607) );
  or2_1 U11459 ( .ip1(n11594), .ip2(n9607), .op(n9609) );
  or2_1 U11460 ( .ip1(n12675), .ip2(n9607), .op(n9608) );
  nand2_1 U11461 ( .ip1(n9609), .ip2(n9608), .op(n11440) );
  or3_1 U11462 ( .ip1(n9611), .ip2(n11564), .ip3(n9610), .op(n11452) );
  inv_1 U11463 ( .ip(n11594), .op(n11494) );
  or2_1 U11464 ( .ip1(n11494), .ip2(n9612), .op(n11358) );
  nand4_1 U11465 ( .ip1(n11441), .ip2(n11440), .ip3(n11452), .ip4(n11358), 
        .op(n9613) );
  not_ab_or_c_or_d U11466 ( .ip1(n11594), .ip2(n9615), .ip3(n9614), .ip4(n9613), .op(n9631) );
  nor3_1 U11467 ( .ip1(n11564), .ip2(n9617), .ip3(n9616), .op(n11333) );
  nor3_1 U11468 ( .ip1(n11564), .ip2(n9619), .ip3(n9618), .op(n11307) );
  nor3_1 U11469 ( .ip1(n11564), .ip2(n9621), .ip3(n9620), .op(n11342) );
  nor3_1 U11470 ( .ip1(n10029), .ip2(n11564), .ip3(n9622), .op(n11498) );
  nor4_1 U11471 ( .ip1(n11333), .ip2(n11307), .ip3(n11342), .ip4(n11498), .op(
        n9630) );
  nand3_1 U11472 ( .ip1(n9623), .ip2(n11501), .ip3(n9624), .op(n9629) );
  nand2_1 U11473 ( .ip1(n9623), .ip2(n9624), .op(n9627) );
  nand2_1 U11474 ( .ip1(n9623), .ip2(n11558), .op(n9626) );
  nand2_1 U11475 ( .ip1(n11583), .ip2(n9624), .op(n9625) );
  nand3_1 U11476 ( .ip1(n9627), .ip2(n9626), .ip3(n9625), .op(n9628) );
  nand2_1 U11477 ( .ip1(n9629), .ip2(n9628), .op(n11458) );
  nand3_1 U11478 ( .ip1(n9631), .ip2(n9630), .ip3(n11458), .op(n9632) );
  nor4_1 U11479 ( .ip1(n11436), .ip2(n11444), .ip3(n11299), .ip4(n9632), .op(
        n9634) );
  nand3_1 U11480 ( .ip1(n9633), .ip2(n11583), .ip3(n12235), .op(n11379) );
  nand4_1 U11481 ( .ip1(n11535), .ip2(n9635), .ip3(n9634), .ip4(n11379), .op(
        n9636) );
  nor4_1 U11482 ( .ip1(n11514), .ip2(n9638), .ip3(n9637), .ip4(n9636), .op(
        n9643) );
  xor2_1 U11483 ( .ip1(n9640), .ip2(n9639), .op(n12246) );
  nand2_1 U11484 ( .ip1(n12246), .ip2(n11578), .op(n11393) );
  xor2_1 U11485 ( .ip1(n9642), .ip2(n9641), .op(n12180) );
  nand2_1 U11486 ( .ip1(n12180), .ip2(n11578), .op(n11304) );
  nand4_1 U11487 ( .ip1(n11204), .ip2(n9643), .ip3(n11393), .ip4(n11304), .op(
        n9644) );
  nor4_1 U11488 ( .ip1(n11483), .ip2(n11466), .ip3(n11415), .ip4(n9644), .op(
        n9649) );
  xor2_1 U11489 ( .ip1(n9646), .ip2(n9645), .op(n10608) );
  nand2_1 U11490 ( .ip1(n10608), .ip2(n11578), .op(n11503) );
  nand2_1 U11491 ( .ip1(n10033), .ip2(n11578), .op(n11491) );
  xor2_1 U11492 ( .ip1(n9648), .ip2(n9647), .op(n12148) );
  nand2_1 U11493 ( .ip1(n12148), .ip2(n11578), .op(n11575) );
  nand4_1 U11494 ( .ip1(n9649), .ip2(n11503), .ip3(n11491), .ip4(n11575), .op(
        n9650) );
  nor4_1 U11495 ( .ip1(n11507), .ip2(n11480), .ip3(n9651), .ip4(n9650), .op(
        n9652) );
  nor2_1 U11496 ( .ip1(n9652), .ip2(\CORTEXM0DS_INST/u_logic/Dw8vx4 ), .op(
        n9653) );
  not_ab_or_c_or_d U11497 ( .ip1(\CORTEXM0DS_INST/u_logic/Dw8vx4 ), .ip2(n9654), .ip3(n9743), .ip4(n9653), .op(n11675) );
  and2_1 U11498 ( .ip1(n12633), .ip2(n9740), .op(n11263) );
  or2_1 U11499 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n11263), .op(
        n9665) );
  nor3_1 U11500 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip3(n11228), .op(n9655) );
  nor2_1 U11501 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(n10698), .op(
        n9725) );
  nor4_1 U11502 ( .ip1(n11209), .ip2(n12116), .ip3(n9655), .ip4(n9725), .op(
        n9662) );
  nand2_1 U11503 ( .ip1(n11250), .ip2(n11692), .op(n9656) );
  nand2_1 U11504 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n9656), .op(
        n9729) );
  nand2_1 U11505 ( .ip1(n9658), .ip2(n9657), .op(n9661) );
  nand3_1 U11506 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip3(n9659), .op(n9660) );
  nand4_1 U11507 ( .ip1(n9662), .ip2(n9729), .ip3(n9661), .ip4(n9660), .op(
        n9663) );
  or2_1 U11508 ( .ip1(n9663), .ip2(n11263), .op(n9664) );
  nand2_1 U11509 ( .ip1(n9665), .ip2(n9664), .op(n11669) );
  mux2_1 U11510 ( .ip1(n11675), .ip2(\CORTEXM0DS_INST/vis_apsr [2]), .s(n11669), .op(n9666) );
  mux2_1 U11511 ( .ip1(n9667), .ip2(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .s(
        n9666), .op(n9761) );
  inv_1 U11512 ( .ip(n9707), .op(n9668) );
  nor2_1 U11513 ( .ip1(n9668), .ip2(n9704), .op(n9713) );
  or2_1 U11514 ( .ip1(n9670), .ip2(n9669), .op(n9676) );
  nand2_1 U11515 ( .ip1(n9686), .ip2(n11832), .op(n9675) );
  inv_1 U11516 ( .ip(n9671), .op(n11854) );
  nor2_1 U11517 ( .ip1(n9673), .ip2(n9672), .op(n9683) );
  nand2_1 U11518 ( .ip1(n11854), .ip2(n9683), .op(n9674) );
  nand3_1 U11519 ( .ip1(n9676), .ip2(n9675), .ip3(n9674), .op(n9694) );
  or2_1 U11520 ( .ip1(n9677), .ip2(n9694), .op(n9679) );
  or2_1 U11521 ( .ip1(n9691), .ip2(n9694), .op(n9678) );
  nand2_1 U11522 ( .ip1(n9679), .ip2(n9678), .op(n9702) );
  inv_1 U11523 ( .ip(n9680), .op(n9692) );
  nand2_1 U11524 ( .ip1(n9682), .ip2(n9681), .op(n9689) );
  inv_1 U11525 ( .ip(n11661), .op(n9684) );
  nand2_1 U11526 ( .ip1(n9684), .ip2(n9683), .op(n9688) );
  nand2_1 U11527 ( .ip1(n9686), .ip2(n9685), .op(n9687) );
  nand3_1 U11528 ( .ip1(n9689), .ip2(n9688), .ip3(n9687), .op(n9690) );
  not_ab_or_c_or_d U11529 ( .ip1(n9692), .ip2(n9691), .ip3(n11796), .ip4(n9690), .op(n9693) );
  not_ab_or_c_or_d U11530 ( .ip1(n9702), .ip2(n11796), .ip3(n9693), .ip4(n9713), .op(n9710) );
  inv_1 U11531 ( .ip(n9694), .op(n9696) );
  nor2_1 U11532 ( .ip1(n9696), .ip2(n9695), .op(n9700) );
  nor2_1 U11533 ( .ip1(n9698), .ip2(n9697), .op(n9699) );
  not_ab_or_c_or_d U11534 ( .ip1(n9701), .ip2(n11840), .ip3(n9700), .ip4(n9699), .op(n9742) );
  or2_1 U11535 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n9702), .op(
        n9703) );
  nand2_1 U11536 ( .ip1(n9742), .ip2(n9703), .op(n9709) );
  nor2_1 U11537 ( .ip1(n9705), .ip2(n9704), .op(n9706) );
  nor2_1 U11538 ( .ip1(n9707), .ip2(n9706), .op(n9708) );
  mux2_1 U11539 ( .ip1(n9710), .ip2(n9709), .s(n9708), .op(n9711) );
  not_ab_or_c_or_d U11540 ( .ip1(n9713), .ip2(\CORTEXM0DS_INST/vis_apsr [1]), 
        .ip3(n9712), .ip4(n9711), .op(n9722) );
  inv_1 U11541 ( .ip(n9714), .op(n9715) );
  nor2_1 U11542 ( .ip1(n9716), .ip2(n9715), .op(n9720) );
  nor2_1 U11543 ( .ip1(n9718), .ip2(n9717), .op(n9719) );
  nor4_1 U11544 ( .ip1(\CORTEXM0DS_INST/u_logic/Dw8vx4 ), .ip2(n9750), .ip3(
        n9720), .ip4(n9719), .op(n9721) );
  nor2_1 U11545 ( .ip1(n9722), .ip2(n9721), .op(n11824) );
  inv_1 U11546 ( .ip(n9853), .op(n9723) );
  nand2_1 U11547 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n11275), .op(
        n10690) );
  nand4_1 U11548 ( .ip1(n11796), .ip2(n9724), .ip3(n9723), .ip4(n10690), .op(
        n9739) );
  inv_1 U11549 ( .ip(n9725), .op(n9726) );
  or2_1 U11550 ( .ip1(n9726), .ip2(n9807), .op(n9728) );
  nand2_1 U11551 ( .ip1(n9728), .ip2(n9727), .op(n9738) );
  inv_1 U11552 ( .ip(n9729), .op(n9731) );
  or2_1 U11553 ( .ip1(n9730), .ip2(n9731), .op(n9733) );
  or2_1 U11554 ( .ip1(n10962), .ip2(n9731), .op(n9732) );
  nand2_1 U11555 ( .ip1(n9733), .ip2(n9732), .op(n9734) );
  or2_1 U11556 ( .ip1(n9807), .ip2(n9734), .op(n9735) );
  nand3_1 U11557 ( .ip1(n9737), .ip2(n9736), .ip3(n9735), .op(n9752) );
  not_ab_or_c_or_d U11558 ( .ip1(n9740), .ip2(n9739), .ip3(n9738), .ip4(n9752), 
        .op(n11826) );
  mux2_1 U11559 ( .ip1(n11824), .ip2(\CORTEXM0DS_INST/vis_apsr [1]), .s(n11826), .op(n9741) );
  not_ab_or_c_or_d U11560 ( .ip1(n10481), .ip2(n9963), .ip3(n10724), .ip4(
        n9741), .op(n9760) );
  nor2_1 U11561 ( .ip1(n10724), .ip2(n10932), .op(n9748) );
  or2_1 U11562 ( .ip1(\CORTEXM0DS_INST/u_logic/Dw8vx4 ), .ip2(n9743), .op(
        n9746) );
  inv_1 U11563 ( .ip(n9742), .op(n9744) );
  or2_1 U11564 ( .ip1(n9744), .ip2(n9743), .op(n9745) );
  nand2_1 U11565 ( .ip1(n9746), .ip2(n9745), .op(n11664) );
  nor2_1 U11566 ( .ip1(n11664), .ip2(n11669), .op(n9747) );
  not_ab_or_c_or_d U11567 ( .ip1(n11669), .ip2(\CORTEXM0DS_INST/vis_apsr [3]), 
        .ip3(n9748), .ip4(n9747), .op(n9758) );
  mux2_1 U11568 ( .ip1(n9750), .ip2(n9749), .s(n10462), .op(n11055) );
  nor3_1 U11569 ( .ip1(n9751), .ip2(n10944), .ip3(n11241), .op(n9753) );
  not_ab_or_c_or_d U11570 ( .ip1(n9754), .ip2(n10421), .ip3(n9753), .ip4(n9752), .op(n11056) );
  mux2_1 U11571 ( .ip1(n11055), .ip2(\CORTEXM0DS_INST/vis_apsr [0]), .s(n11056), .op(n9755) );
  nor3_1 U11572 ( .ip1(n10500), .ip2(n9756), .ip3(n9755), .op(n9757) );
  xor2_1 U11573 ( .ip1(n9758), .ip2(n9757), .op(n9759) );
  not_ab_or_c_or_d U11574 ( .ip1(n9761), .ip2(n12583), .ip3(n9760), .ip4(n9759), .op(n9762) );
  mux2_1 U11575 ( .ip1(n11190), .ip2(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .s(
        n9762), .op(n10963) );
  nor4_1 U11576 ( .ip1(n9882), .ip2(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip3(
        n10963), .ip4(n11100), .op(n9770) );
  nand2_1 U11577 ( .ip1(n12588), .ip2(n10930), .op(n9764) );
  nor4_1 U11578 ( .ip1(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/I29vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/P39vx4 ), .ip4(n11112), .op(n10496) );
  inv_1 U11579 ( .ip(n10496), .op(n10826) );
  nor2_1 U11580 ( .ip1(\CORTEXM0DS_INST/u_logic/K79vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/W49vx4 ), .op(n9947) );
  nand3_1 U11581 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n9947), .ip3(
        n12571), .op(n10825) );
  nand2_1 U11582 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n12562), .op(
        n10494) );
  nor4_1 U11583 ( .ip1(n12588), .ip2(n10826), .ip3(n10825), .ip4(n10494), .op(
        n9763) );
  not_ab_or_c_or_d U11584 ( .ip1(n12583), .ip2(n9764), .ip3(n9763), .ip4(
        n12538), .op(n9765) );
  nor3_1 U11585 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n9765), .ip3(
        n11100), .op(n9769) );
  nor2_1 U11586 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n10835), .op(
        n10620) );
  nor3_1 U11587 ( .ip1(n9834), .ip2(n10620), .ip3(n10539), .op(n9768) );
  nand2_1 U11588 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n12567), .op(
        n10546) );
  nor4_1 U11589 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/K79vx4 ), .ip3(n11190), .ip4(n12571), .op(
        n9939) );
  inv_1 U11590 ( .ip(n10500), .op(n9766) );
  not_ab_or_c_or_d U11591 ( .ip1(n12571), .ip2(n10546), .ip3(n9939), .ip4(
        n9766), .op(n10976) );
  nor2_1 U11592 ( .ip1(n10976), .ip2(n10542), .op(n9767) );
  or4_1 U11593 ( .ip1(n9770), .ip2(n9769), .ip3(n9768), .ip4(n9767), .op(n9795) );
  nor4_1 U11594 ( .ip1(n11232), .ip2(n11080), .ip3(n9771), .ip4(n10697), .op(
        n9877) );
  nor3_1 U11595 ( .ip1(n11131), .ip2(n9772), .ip3(n12118), .op(n9775) );
  nand2_1 U11596 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(n5639), .op(
        n10706) );
  mux2_1 U11597 ( .ip1(n12567), .ip2(\CORTEXM0DS_INST/u_logic/K79vx4 ), .s(
        \CORTEXM0DS_INST/u_logic/D69vx4 ), .op(n11111) );
  nand4_1 U11598 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/R89vx4 ), .ip4(n11111), .op(n10621) );
  nor4_1 U11599 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n10848), .ip3(
        n10706), .ip4(n10621), .op(n9774) );
  nor2_1 U11600 ( .ip1(n5932), .ip2(n9773), .op(n10752) );
  inv_1 U11601 ( .ip(n9817), .op(n10677) );
  nand2_1 U11602 ( .ip1(n10677), .ip2(n9785), .op(n12637) );
  nand2_1 U11603 ( .ip1(n10752), .ip2(n12637), .op(n9863) );
  nor4_1 U11604 ( .ip1(n9877), .ip2(n9775), .ip3(n9774), .ip4(n9863), .op(
        n9793) );
  not_ab_or_c_or_d U11605 ( .ip1(n10734), .ip2(n9776), .ip3(n11686), .ip4(
        n11803), .op(n9792) );
  nor2_1 U11606 ( .ip1(n12592), .ip2(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .op(
        n11102) );
  and4_1 U11607 ( .ip1(n12122), .ip2(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip3(
        n11102), .ip4(n10551), .op(n9778) );
  not_ab_or_c_or_d U11608 ( .ip1(n12610), .ip2(n9962), .ip3(n9778), .ip4(n9777), .op(n9781) );
  nand3_1 U11609 ( .ip1(n9781), .ip2(n9780), .ip3(n9779), .op(n9784) );
  nor3_1 U11610 ( .ip1(n10512), .ip2(n10842), .ip3(n10706), .op(n9783) );
  nor2_1 U11611 ( .ip1(n11253), .ip2(n9927), .op(n9782) );
  not_ab_or_c_or_d U11612 ( .ip1(n5639), .ip2(n9784), .ip3(n9783), .ip4(n9782), 
        .op(n9791) );
  nand2_1 U11613 ( .ip1(n9785), .ip2(n12117), .op(n11136) );
  nor3_1 U11614 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n11786), .ip3(
        n11136), .op(n11751) );
  or2_1 U11615 ( .ip1(n12624), .ip2(n9785), .op(n9787) );
  or2_1 U11616 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n9785), .op(
        n9786) );
  nand2_1 U11617 ( .ip1(n9787), .ip2(n9786), .op(n11011) );
  nor2_1 U11618 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Ki8vx4 ), .op(n9929) );
  nor3_1 U11619 ( .ip1(n11011), .ip2(n9929), .ip3(n12126), .op(n9788) );
  nor4_1 U11620 ( .ip1(n11802), .ip2(n9789), .ip3(n11751), .ip4(n9788), .op(
        n9790) );
  nand4_1 U11621 ( .ip1(n9793), .ip2(n9792), .ip3(n9791), .ip4(n9790), .op(
        n9794) );
  not_ab_or_c_or_d U11622 ( .ip1(n12618), .ip2(n9795), .ip3(n10052), .ip4(
        n9794), .op(n9796) );
  not_ab_or_c_or_d U11623 ( .ip1(n5932), .ip2(n9797), .ip3(1'b0), .ip4(n9796), 
        .op(\CORTEXM0DS_INST/u_logic/Eyhvx4 ) );
  nand3_1 U11624 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n9798), .ip3(
        n10632), .op(n9801) );
  nand2_1 U11625 ( .ip1(n9799), .ip2(n9962), .op(n9800) );
  nand2_1 U11626 ( .ip1(n9801), .ip2(n9800), .op(n9851) );
  not_ab_or_c_or_d U11627 ( .ip1(n10944), .ip2(n10690), .ip3(n10892), .ip4(
        n12628), .op(n9803) );
  nor2_1 U11628 ( .ip1(n10670), .ip2(n10671), .op(n9802) );
  not_ab_or_c_or_d U11629 ( .ip1(n12116), .ip2(n10770), .ip3(n9803), .ip4(
        n9802), .op(n9804) );
  nor2_1 U11630 ( .ip1(n9804), .ip2(n10851), .op(n9850) );
  nand2_1 U11631 ( .ip1(n9955), .ip2(n12588), .op(n10540) );
  inv_1 U11632 ( .ip(n10540), .op(n9814) );
  nand2_1 U11633 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n12583), .op(
        n10718) );
  inv_1 U11634 ( .ip(n10718), .op(n10713) );
  nor2_1 U11635 ( .ip1(\CORTEXM0DS_INST/u_logic/K79vx4 ), .ip2(n10713), .op(
        n9805) );
  nor2_1 U11636 ( .ip1(n11190), .ip2(n12571), .op(n10625) );
  not_ab_or_c_or_d U11637 ( .ip1(n9828), .ip2(n12583), .ip3(n9805), .ip4(
        n10625), .op(n9806) );
  nor2_1 U11638 ( .ip1(n9806), .ip2(n10491), .op(n9810) );
  not_ab_or_c_or_d U11639 ( .ip1(n11102), .ip2(n9808), .ip3(
        \CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip4(n9807), .op(n9809) );
  not_ab_or_c_or_d U11640 ( .ip1(n12320), .ip2(
        \CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip3(n9810), .ip4(n9809), .op(n9811) );
  nor2_1 U11641 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(n9811), .op(
        n9813) );
  nor4_1 U11642 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n9929), .ip3(
        n11240), .ip4(n11223), .op(n9812) );
  not_ab_or_c_or_d U11643 ( .ip1(n9814), .ip2(n10512), .ip3(n9813), .ip4(n9812), .op(n9848) );
  nor2_1 U11644 ( .ip1(n9815), .ip2(n10770), .op(n9816) );
  nor4_1 U11645 ( .ip1(n11679), .ip2(n10611), .ip3(n9816), .ip4(n11277), .op(
        n9819) );
  nor2_1 U11646 ( .ip1(n9817), .ip2(n11136), .op(n9818) );
  not_ab_or_c_or_d U11647 ( .ip1(n9946), .ip2(n12369), .ip3(n9819), .ip4(n9818), .op(n9847) );
  nor2_1 U11648 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n9807), .op(
        n9825) );
  inv_1 U11649 ( .ip(n10690), .op(n9821) );
  nor3_1 U11650 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip3(n11786), .op(n9820) );
  not_ab_or_c_or_d U11651 ( .ip1(n12641), .ip2(n10611), .ip3(n9821), .ip4(
        n9820), .op(n9822) );
  nor2_1 U11652 ( .ip1(n9822), .ip2(n10865), .op(n9824) );
  and4_1 U11653 ( .ip1(n10932), .ip2(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip4(n10647), .op(n9823) );
  not_ab_or_c_or_d U11654 ( .ip1(n9825), .ip2(n10734), .ip3(n9824), .ip4(n9823), .op(n9846) );
  and2_1 U11655 ( .ip1(n12125), .ip2(n10556), .op(n9844) );
  or4_1 U11656 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n9947), .ip3(
        n12562), .ip4(n12571), .op(n9826) );
  nand2_1 U11657 ( .ip1(n9955), .ip2(n9826), .op(n9827) );
  not_ab_or_c_or_d U11658 ( .ip1(n10491), .ip2(n9827), .ip3(n10492), .ip4(
        n12538), .op(n9843) );
  not_ab_or_c_or_d U11659 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(
        n12567), .ip3(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip4(n9828), .op(
        n9829) );
  nor2_1 U11660 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n12599), .op(
        n10884) );
  inv_1 U11661 ( .ip(n10884), .op(n10624) );
  nor2_1 U11662 ( .ip1(n9829), .ip2(n10624), .op(n9830) );
  or2_1 U11663 ( .ip1(n10481), .ip2(n9830), .op(n9831) );
  nand2_1 U11664 ( .ip1(n10206), .ip2(n9831), .op(n9832) );
  nor2_1 U11665 ( .ip1(n9832), .ip2(n10646), .op(n9842) );
  inv_1 U11666 ( .ip(n9833), .op(n10422) );
  not_ab_or_c_or_d U11667 ( .ip1(n11786), .ip2(n10422), .ip3(
        \CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip4(n10631), .op(n9840) );
  nand3_1 U11668 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip3(n9834), .op(n10705) );
  or2_1 U11669 ( .ip1(n10705), .ip2(n11100), .op(n9837) );
  nor2_1 U11670 ( .ip1(n10835), .ip2(n12321), .op(n11093) );
  inv_1 U11671 ( .ip(n11093), .op(n9835) );
  or2_1 U11672 ( .ip1(n9835), .ip2(n11100), .op(n9836) );
  nand2_1 U11673 ( .ip1(n9837), .ip2(n9836), .op(n9839) );
  nor2_1 U11674 ( .ip1(n9838), .ip2(n10851), .op(n11787) );
  or4_1 U11675 ( .ip1(n9840), .ip2(n9839), .ip3(n11787), .ip4(n5420), .op(
        n9841) );
  nor4_1 U11676 ( .ip1(n9844), .ip2(n9843), .ip3(n9842), .ip4(n9841), .op(
        n9845) );
  nand4_1 U11677 ( .ip1(n9848), .ip2(n9847), .ip3(n9846), .ip4(n9845), .op(
        n9849) );
  not_ab_or_c_or_d U11678 ( .ip1(n10892), .ip2(n9851), .ip3(n9850), .ip4(n9849), .op(n9852) );
  not_ab_or_c_or_d U11679 ( .ip1(n5932), .ip2(n11228), .ip3(1'b0), .ip4(n9852), 
        .op(\CORTEXM0DS_INST/u_logic/Fvhvx4 ) );
  nand2_1 U11680 ( .ip1(n11051), .ip2(n10992), .op(n10956) );
  nor2_1 U11681 ( .ip1(n12117), .ip2(n10956), .op(n9857) );
  nand2_1 U11682 ( .ip1(n11208), .ip2(n10992), .op(n10987) );
  nor2_1 U11683 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n10987), .op(
        n9856) );
  nand2_1 U11684 ( .ip1(n9853), .ip2(n10670), .op(n10950) );
  nor3_1 U11685 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n10949), .ip3(
        n11788), .op(n10981) );
  inv_1 U11686 ( .ip(n10981), .op(n9854) );
  nor2_1 U11687 ( .ip1(n10950), .ip2(n9854), .op(n9855) );
  or4_1 U11688 ( .ip1(n9858), .ip2(n9857), .ip3(n9856), .ip4(n9855), .op(n9911) );
  nor2_1 U11689 ( .ip1(n10971), .ip2(n12070), .op(n11247) );
  inv_1 U11690 ( .ip(n11249), .op(n9859) );
  nand3_1 U11691 ( .ip1(n10805), .ip2(n10734), .ip3(n11782), .op(n10569) );
  nor2_1 U11692 ( .ip1(n9859), .ip2(n10569), .op(n9862) );
  nor3_1 U11693 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip3(n10722), .op(n11791) );
  inv_1 U11694 ( .ip(n11076), .op(n9860) );
  nor3_1 U11695 ( .ip1(\CORTEXM0DS_INST/u_logic/Q5gvx4 ), .ip2(n11786), .ip3(
        n9860), .op(n10045) );
  nor2_1 U11696 ( .ip1(n11791), .ip2(n10045), .op(n10996) );
  inv_1 U11697 ( .ip(n10996), .op(n9861) );
  not_ab_or_c_or_d U11698 ( .ip1(n11247), .ip2(
        \CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip3(n9862), .ip4(n9861), .op(n9880) );
  nand2_1 U11699 ( .ip1(n12656), .ip2(n10652), .op(n11184) );
  nor2_1 U11700 ( .ip1(n11796), .ip2(n11184), .op(n9864) );
  not_ab_or_c_or_d U11701 ( .ip1(n9865), .ip2(n10478), .ip3(n9864), .ip4(n9863), .op(n9879) );
  nor2_1 U11702 ( .ip1(n8424), .ip2(n10949), .op(n10741) );
  inv_1 U11703 ( .ip(n10741), .op(n9887) );
  or2_1 U11704 ( .ip1(n9887), .ip2(n12131), .op(n9867) );
  or2_1 U11705 ( .ip1(n10988), .ip2(n12131), .op(n9866) );
  nand2_1 U11706 ( .ip1(n9867), .ip2(n9866), .op(n9876) );
  nand3_1 U11707 ( .ip1(n9870), .ip2(n9869), .ip3(n9868), .op(n9871) );
  or2_1 U11708 ( .ip1(n9871), .ip2(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .op(
        n9874) );
  nand2_1 U11709 ( .ip1(n10636), .ip2(n11190), .op(n10824) );
  nand2_1 U11710 ( .ip1(n10965), .ip2(n10824), .op(n9872) );
  or2_1 U11711 ( .ip1(n9872), .ip2(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .op(
        n9873) );
  nand2_1 U11712 ( .ip1(n9874), .ip2(n9873), .op(n9875) );
  not_ab_or_c_or_d U11713 ( .ip1(n9877), .ip2(n12125), .ip3(n9876), .ip4(n9875), .op(n9878) );
  nor2_1 U11714 ( .ip1(n10706), .ip2(n10218), .op(n10928) );
  nand2_1 U11715 ( .ip1(n10928), .ip2(n12599), .op(n10936) );
  nand4_1 U11716 ( .ip1(n9880), .ip2(n9879), .ip3(n9878), .ip4(n10936), .op(
        n9910) );
  nor2_1 U11717 ( .ip1(n12567), .ip2(n9881), .op(n9883) );
  nand4_1 U11718 ( .ip1(n9882), .ip2(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip3(
        n10496), .ip4(n10928), .op(n10926) );
  nor4_1 U11719 ( .ip1(\CORTEXM0DS_INST/u_logic/D69vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/R89vx4 ), .ip3(n9883), .ip4(n10926), .op(
        n9891) );
  nand2_1 U11720 ( .ip1(n10500), .ip2(n11146), .op(n9965) );
  nor2_1 U11721 ( .ip1(n9884), .ip2(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .op(
        n10991) );
  nand2_1 U11722 ( .ip1(n10991), .ip2(n10492), .op(n9885) );
  not_ab_or_c_or_d U11723 ( .ip1(n9886), .ip2(n9965), .ip3(n12592), .ip4(n9885), .op(n9890) );
  nor3_1 U11724 ( .ip1(n11796), .ip2(n11793), .ip3(n9887), .op(n9889) );
  inv_1 U11725 ( .ip(n10992), .op(n10563) );
  nor3_1 U11726 ( .ip1(n12117), .ip2(n10971), .ip3(n10563), .op(n9888) );
  nor4_1 U11727 ( .ip1(n9891), .ip2(n9890), .ip3(n9889), .ip4(n9888), .op(
        n9908) );
  inv_1 U11728 ( .ip(n11243), .op(n9893) );
  inv_1 U11729 ( .ip(n9892), .op(n10984) );
  nand2_1 U11730 ( .ip1(n10928), .ip2(n9933), .op(n10978) );
  nor2_1 U11731 ( .ip1(n10979), .ip2(n10978), .op(n10939) );
  nor4_1 U11732 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip3(n12623), .ip4(n11789), .op(
        n10044) );
  not_ab_or_c_or_d U11733 ( .ip1(n9893), .ip2(n10984), .ip3(n10939), .ip4(
        n10044), .op(n9907) );
  nand2_1 U11734 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Cf9vx4 ), .op(n9895) );
  or2_1 U11735 ( .ip1(n12538), .ip2(n10715), .op(n9894) );
  not_ab_or_c_or_d U11736 ( .ip1(n9895), .ip2(n9894), .ip3(n11088), .ip4(
        n10740), .op(n9904) );
  nor2_1 U11737 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n12571), .op(
        n9897) );
  nand2_1 U11738 ( .ip1(n11190), .ip2(n12567), .op(n9950) );
  nand4_1 U11739 ( .ip1(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/B19vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/I29vx4 ), .ip4(
        \CORTEXM0DS_INST/u_logic/R89vx4 ), .op(n10841) );
  nor3_1 U11740 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip3(n10841), .op(n9896) );
  not_ab_or_c_or_d U11741 ( .ip1(n9897), .ip2(n9950), .ip3(n10500), .ip4(n9896), .op(n9898) );
  nand3_1 U11742 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n10636), .ip3(
        n12571), .op(n10493) );
  nand3_1 U11743 ( .ip1(n10635), .ip2(n10551), .ip3(n10991), .op(n10921) );
  not_ab_or_c_or_d U11744 ( .ip1(n9898), .ip2(n10493), .ip3(n10921), .ip4(
        n10492), .op(n9903) );
  nand2_1 U11745 ( .ip1(n9899), .ip2(n11190), .op(n9901) );
  nand3_1 U11746 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(n12592), .ip3(
        n12125), .op(n9900) );
  not_ab_or_c_or_d U11747 ( .ip1(n10806), .ip2(n9901), .ip3(
        \CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip4(n9900), .op(n9902) );
  nor3_1 U11748 ( .ip1(n9904), .ip2(n9903), .ip3(n9902), .op(n9906) );
  nand4_1 U11749 ( .ip1(n9908), .ip2(n9907), .ip3(n9906), .ip4(n9905), .op(
        n9909) );
  not_ab_or_c_or_d U11750 ( .ip1(n10892), .ip2(n9911), .ip3(n9910), .ip4(n9909), .op(n9912) );
  not_ab_or_c_or_d U11751 ( .ip1(n5932), .ip2(n12623), .ip3(1'b0), .ip4(n9912), 
        .op(\CORTEXM0DS_INST/u_logic/Ruhvx4 ) );
  nor2_1 U11752 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [10]), .ip2(n9919), 
        .op(n9913) );
  or2_1 U11753 ( .ip1(n12739), .ip2(n9913), .op(n2543) );
  nor2_1 U11754 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [15]), .ip2(n9919), 
        .op(n9914) );
  or2_1 U11755 ( .ip1(n12741), .ip2(n9914), .op(n2463) );
  nor2_1 U11756 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [8]), .ip2(n9919), .op(
        n9915) );
  or2_1 U11757 ( .ip1(n12742), .ip2(n9915), .op(n2511) );
  nor2_1 U11758 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [12]), .ip2(n9919), 
        .op(n9916) );
  or2_1 U11759 ( .ip1(n12743), .ip2(n9916), .op(n2647) );
  nor2_1 U11760 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [0]), .ip2(n9919), .op(
        n9917) );
  or2_1 U11761 ( .ip1(n12744), .ip2(n9917), .op(n2790) );
  nor2_1 U11762 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [3]), .ip2(n9919), .op(
        n9918) );
  or2_1 U11763 ( .ip1(n12745), .ip2(n9918), .op(n2626) );
  nor2_1 U11764 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [6]), .ip2(n9919), .op(
        n9920) );
  or2_1 U11765 ( .ip1(n12746), .ip2(n9920), .op(n2713) );
  nor3_1 U11766 ( .ip1(n9921), .ip2(n12686), .ip3(n12687), .op(n3224) );
  inv_1 U11767 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [6]), .op(n11941) );
  inv_1 U11768 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [5]), .op(n11937) );
  nand2_1 U11769 ( .ip1(n11941), .ip2(n11937), .op(n11946) );
  or2_1 U11770 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [16]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [17]), .op(n12014) );
  or4_1 U11771 ( .ip1(n11946), .ip2(n12014), .ip3(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [14]), .ip4(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [13]), .op(n9926) );
  nor4_1 U11772 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [23]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [22]), .ip3(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [20]), .ip4(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [21]), .op(n9924) );
  nor4_1 U11773 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [15]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [12]), .ip3(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [19]), .ip4(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [18]), .op(n9923) );
  nor3_1 U11774 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [9]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [10]), .ip3(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [8]), .op(n11973) );
  nor4_1 U11775 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [4]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [3]), .ip3(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [1]), .ip4(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [2]), .op(n9922) );
  nand4_1 U11776 ( .ip1(n9924), .ip2(n9923), .ip3(n11973), .ip4(n9922), .op(
        n9925) );
  nor4_1 U11777 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [11]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [7]), .ip3(n9926), .ip4(n9925), .op(
        n11908) );
  and4_1 U11778 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [0]), .ip2(
        \CORTEXM0DS_INST/u_logic/F2hvx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/S0hvx4 ), .ip4(n11908), .op(n2326) );
  inv_1 U11779 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [7]), .op(n3223) );
  nor2_1 U11780 ( .ip1(n9928), .ip2(n9927), .op(n9985) );
  nor3_1 U11781 ( .ip1(n11131), .ip2(n12118), .ip3(n11682), .op(n9931) );
  nor3_1 U11782 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n9929), .ip3(
        n11789), .op(n9930) );
  or2_1 U11783 ( .ip1(n9931), .ip2(n9930), .op(n9982) );
  nand2_1 U11784 ( .ip1(n10979), .ip2(n12588), .op(n10821) );
  inv_1 U11785 ( .ip(n10821), .op(n9932) );
  nor2_1 U11786 ( .ip1(n9933), .ip2(n9932), .op(n10844) );
  nor3_1 U11787 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/K79vx4 ), .op(n10499) );
  nor2_1 U11788 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n10623), .op(
        n9934) );
  or2_1 U11789 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n9934), .op(
        n9936) );
  nand2_1 U11790 ( .ip1(n11190), .ip2(n10841), .op(n10720) );
  or2_1 U11791 ( .ip1(n10720), .ip2(n9934), .op(n9935) );
  nand2_1 U11792 ( .ip1(n9936), .ip2(n9935), .op(n10503) );
  nor2_1 U11793 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(n10835), .op(
        n10205) );
  nand3_1 U11794 ( .ip1(n10503), .ip2(n10205), .ip3(n9937), .op(n9938) );
  not_ab_or_c_or_d U11795 ( .ip1(n10844), .ip2(n10499), .ip3(n9939), .ip4(
        n9938), .op(n9940) );
  not_ab_or_c_or_d U11796 ( .ip1(n11100), .ip2(n10492), .ip3(n9940), .ip4(
        n10842), .op(n9981) );
  inv_1 U11797 ( .ip(n11218), .op(n9942) );
  nor2_1 U11798 ( .ip1(n12118), .ip2(n11228), .op(n10202) );
  not_ab_or_c_or_d U11799 ( .ip1(n9942), .ip2(n9941), .ip3(n5420), .ip4(n10202), .op(n9979) );
  inv_1 U11800 ( .ip(n11136), .op(n9944) );
  nor2_1 U11801 ( .ip1(n12623), .ip2(n9943), .op(n10776) );
  not_ab_or_c_or_d U11802 ( .ip1(n9946), .ip2(n9945), .ip3(n9944), .ip4(n10776), .op(n9978) );
  nand2_1 U11803 ( .ip1(n10496), .ip2(n9947), .op(n9949) );
  not_ab_or_c_or_d U11804 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n9949), .ip3(n10820), .ip4(n9948), .op(n9951) );
  nand4_1 U11805 ( .ip1(\CORTEXM0DS_INST/u_logic/D69vx4 ), .ip2(n9951), .ip3(
        n9950), .ip4(n12571), .op(n9954) );
  nor2_1 U11806 ( .ip1(n9952), .ip2(n10646), .op(n9953) );
  not_ab_or_c_or_d U11807 ( .ip1(n9955), .ip2(n9954), .ip3(n10652), .ip4(n9953), .op(n9977) );
  nor2_1 U11808 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(n10988), .op(
        n10514) );
  nor2_1 U11809 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10988), .op(
        n9975) );
  or2_1 U11810 ( .ip1(n9956), .ip2(n9957), .op(n9959) );
  or2_1 U11811 ( .ip1(n10690), .ip2(n9957), .op(n9958) );
  nand2_1 U11812 ( .ip1(n9959), .ip2(n9958), .op(n9974) );
  inv_1 U11813 ( .ip(n11277), .op(n12134) );
  nor2_1 U11814 ( .ip1(n11223), .ip2(n10671), .op(n9961) );
  nor2_1 U11815 ( .ip1(n10610), .ip2(n10972), .op(n9960) );
  not_ab_or_c_or_d U11816 ( .ip1(n11213), .ip2(n12134), .ip3(n9961), .ip4(
        n9960), .op(n9972) );
  nand2_1 U11817 ( .ip1(n9962), .ip2(n10770), .op(n9971) );
  inv_1 U11818 ( .ip(n9963), .op(n10819) );
  nand2_1 U11819 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n10819), .op(
        n9966) );
  nand2_1 U11820 ( .ip1(n10636), .ip2(n10647), .op(n9964) );
  nand3_1 U11821 ( .ip1(n9966), .ip2(n9965), .ip3(n9964), .op(n9967) );
  nand2_1 U11822 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n9967), .op(
        n9970) );
  nand2_1 U11823 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n9968), .op(
        n9969) );
  nand4_1 U11824 ( .ip1(n9972), .ip2(n9971), .ip3(n9970), .ip4(n9969), .op(
        n9973) );
  nor4_1 U11825 ( .ip1(n10514), .ip2(n9975), .ip3(n9974), .ip4(n9973), .op(
        n9976) );
  nand4_1 U11826 ( .ip1(n9979), .ip2(n9978), .ip3(n9977), .ip4(n9976), .op(
        n9980) );
  not_ab_or_c_or_d U11827 ( .ip1(n10955), .ip2(n9982), .ip3(n9981), .ip4(n9980), .op(n9983) );
  not_ab_or_c_or_d U11828 ( .ip1(n5932), .ip2(n11693), .ip3(1'b0), .ip4(n9983), 
        .op(n9984) );
  or2_1 U11829 ( .ip1(n9985), .ip2(n9984), .op(
        \CORTEXM0DS_INST/u_logic/Qxhvx4 ) );
  inv_1 U11830 ( .ip(n9986), .op(n5913) );
  or2_1 U11831 ( .ip1(n5913), .ip2(n9987), .op(\interconnect_ip_inst/n6491 )
         );
  inv_1 U11832 ( .ip(\CORTEXM0DS_INST/vis_pc [30]), .op(n9989) );
  nor2_1 U11833 ( .ip1(n10457), .ip2(n9988), .op(n10030) );
  mux2_1 U11834 ( .ip1(n9989), .ip2(\CORTEXM0DS_INST/vis_pc [30]), .s(n10030), 
        .op(n5881) );
  nor2_1 U11835 ( .ip1(n12343), .ip2(n5881), .op(n9993) );
  nand2_1 U11836 ( .ip1(n10462), .ip2(n12352), .op(n9992) );
  nand2_1 U11837 ( .ip1(n12316), .ip2(n9990), .op(n9991) );
  nand2_1 U11838 ( .ip1(n9992), .ip2(n9991), .op(n10038) );
  nor2_1 U11839 ( .ip1(n9993), .ip2(n10038), .op(
        \CORTEXM0DS_INST/u_logic/N4518 ) );
  nand2_1 U11840 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(n12679), .op(
        n6175) );
  nor2_1 U11841 ( .ip1(n11705), .ip2(n6175), .op(n9994) );
  or2_1 U11842 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [5]), .ip2(n9994), .op(
        n9995) );
  nand2_1 U11843 ( .ip1(n9995), .ip2(n2683), .op(n9998) );
  nor2_1 U11844 ( .ip1(n11895), .ip2(n9996), .op(n9997) );
  nor2_1 U11845 ( .ip1(n9998), .ip2(n9997), .op(
        \CORTEXM0DS_INST/u_logic/K1ivx4 ) );
  nand2_1 U11846 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(n12675), .op(
        n6170) );
  nor2_1 U11847 ( .ip1(n11705), .ip2(n6170), .op(n9999) );
  or2_1 U11848 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [4]), .ip2(n9999), .op(
        n10000) );
  nand2_1 U11849 ( .ip1(n10000), .ip2(n2641), .op(n10003) );
  nor2_1 U11850 ( .ip1(n11895), .ip2(n10001), .op(n10002) );
  nor2_1 U11851 ( .ip1(n10003), .ip2(n10002), .op(
        \CORTEXM0DS_INST/u_logic/R1ivx4 ) );
  inv_1 U11852 ( .ip(\interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state [2]), 
        .op(n10005) );
  inv_1 U11853 ( .ip(\interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state [0]), 
        .op(n10015) );
  nand2_1 U11854 ( .ip1(n5933), .ip2(n10015), .op(n10004) );
  nand2_1 U11855 ( .ip1(n10005), .ip2(n10004), .op(
        \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_nextstate [2]) );
  or2_1 U11856 ( .ip1(\interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state [2]), 
        .ip2(n5934), .op(n10013) );
  nand3_1 U11857 ( .ip1(n10013), .ip2(
        \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state [0]), .ip3(
        \interconnect_ip_inst/i_apb_hready_resp ), .op(n10007) );
  or2_1 U11858 ( .ip1(\interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state [0]), 
        .ip2(\interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_nextstate [2]), .op(
        n10006) );
  nand2_1 U11859 ( .ip1(n10007), .ip2(n10006), .op(
        \interconnect_ip_inst/n4829 ) );
  inv_1 U11860 ( .ip(n5929), .op(n10009) );
  nand2_1 U11861 ( .ip1(n5932), .ip2(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [2]), .op(n10008) );
  nand2_1 U11862 ( .ip1(n10009), .ip2(n10008), .op(
        \interconnect_ip_inst/n4862 ) );
  nand2_1 U11863 ( .ip1(n5932), .ip2(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [3]), .op(n10010) );
  nand2_1 U11864 ( .ip1(n5928), .ip2(n10010), .op(\interconnect_ip_inst/n4863 ) );
  nand2_1 U11865 ( .ip1(n5932), .ip2(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [4]), .op(n10011) );
  nand2_1 U11866 ( .ip1(n5924), .ip2(n10011), .op(\interconnect_ip_inst/n4864 ) );
  inv_1 U11867 ( .ip(\interconnect_ip_inst/i_ahb_U_dfltslv_current_state ), 
        .op(n10012) );
  nand2_1 U11868 ( .ip1(n5921), .ip2(n10012), .op(
        \interconnect_ip_inst/i_ahb_U_dfltslv_N4 ) );
  or2_1 U11869 ( .ip1(n5917), .ip2(n10013), .op(n10014) );
  nand2_1 U11870 ( .ip1(n10015), .ip2(n10014), .op(
        \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_nextstate [0]) );
  nor2_1 U11871 ( .ip1(\interconnect_ip_inst/i_ahb_U_dfltslv_current_state ), 
        .ip2(n5921), .op(\interconnect_ip_inst/n10765 ) );
  inv_1 U11872 ( .ip(n10016), .op(n12323) );
  nand2_1 U11873 ( .ip1(n10017), .ip2(n12323), .op(
        \CORTEXM0DS_INST/u_logic/N4816 ) );
  nand3_1 U11874 ( .ip1(n12162), .ip2(\CORTEXM0DS_INST/vis_pc [8]), .ip3(
        \CORTEXM0DS_INST/vis_pc [9]), .op(n12186) );
  nor2_1 U11875 ( .ip1(n10193), .ip2(n12186), .op(n12195) );
  inv_1 U11876 ( .ip(n12195), .op(n10019) );
  nand2_1 U11877 ( .ip1(\CORTEXM0DS_INST/vis_pc [12]), .ip2(n12195), .op(
        n10024) );
  inv_1 U11878 ( .ip(n10024), .op(n10018) );
  not_ab_or_c_or_d U11879 ( .ip1(n10197), .ip2(n10019), .ip3(n10018), .ip4(
        n12343), .op(n10021) );
  nor2_1 U11880 ( .ip1(n10194), .ip2(n12311), .op(n10020) );
  not_ab_or_c_or_d U11881 ( .ip1(n12316), .ip2(n10022), .ip3(n10021), .ip4(
        n10020), .op(\CORTEXM0DS_INST/u_logic/N4767 ) );
  inv_1 U11882 ( .ip(n11006), .op(n10023) );
  not_ab_or_c_or_d U11883 ( .ip1(n10329), .ip2(n10024), .ip3(n10023), .ip4(
        n12343), .op(n10026) );
  nor2_1 U11884 ( .ip1(n10330), .ip2(n12311), .op(n10025) );
  not_ab_or_c_or_d U11885 ( .ip1(n12316), .ip2(n10027), .ip3(n10026), .ip4(
        n10025), .op(\CORTEXM0DS_INST/u_logic/N4751 ) );
  nand3_1 U11886 ( .ip1(n10028), .ip2(n1520), .ip3(n11201), .op(
        \CORTEXM0DS_INST/u_logic/N4674 ) );
  nor2_1 U11887 ( .ip1(n10029), .ip2(n12347), .op(n10032) );
  inv_1 U11888 ( .ip(\CORTEXM0DS_INST/vis_pc [29]), .op(n10601) );
  nand3_1 U11889 ( .ip1(\CORTEXM0DS_INST/vis_pc [27]), .ip2(
        \CORTEXM0DS_INST/vis_pc [28]), .ip3(n12308), .op(n10035) );
  not_ab_or_c_or_d U11890 ( .ip1(n10601), .ip2(n10035), .ip3(n10030), .ip4(
        n12343), .op(n10031) );
  not_ab_or_c_or_d U11891 ( .ip1(n12352), .ip2(n10608), .ip3(n10032), .ip4(
        n10031), .op(\CORTEXM0DS_INST/u_logic/N4439 ) );
  nand2_1 U11892 ( .ip1(n10033), .ip2(n12352), .op(n10039) );
  or2_1 U11893 ( .ip1(\CORTEXM0DS_INST/vis_pc [28]), .ip2(n10034), .op(n10036)
         );
  nand3_1 U11894 ( .ip1(n12605), .ip2(n10036), .ip3(n10035), .op(n10037) );
  nand2_1 U11895 ( .ip1(n10039), .ip2(n10037), .op(
        \CORTEXM0DS_INST/u_logic/E562z4 ) );
  or2_1 U11896 ( .ip1(n5885), .ip2(n10038), .op(n5886) );
  inv_1 U11897 ( .ip(n10039), .op(n5880) );
  nor2_1 U11898 ( .ip1(n10040), .ip2(n12347), .op(
        \CORTEXM0DS_INST/u_logic/Q462z4 ) );
  nor2_1 U11899 ( .ip1(n12605), .ip2(n10041), .op(
        \CORTEXM0DS_INST/u_logic/A362z4 ) );
  nor2_1 U11900 ( .ip1(n10949), .ip2(n10973), .op(n10786) );
  nor3_1 U11901 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Q5gvx4 ), .ip3(n10972), .op(n10042) );
  not_ab_or_c_or_d U11902 ( .ip1(n12617), .ip2(n10043), .ip3(n10786), .ip4(
        n10042), .op(n10057) );
  not_ab_or_c_or_d U11903 ( .ip1(n10953), .ip2(n12641), .ip3(n10045), .ip4(
        n10044), .op(n10056) );
  inv_1 U11904 ( .ip(n10983), .op(n10046) );
  or2_1 U11905 ( .ip1(n10046), .ip2(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .op(
        n10049) );
  nand2_1 U11906 ( .ip1(n11132), .ip2(n10992), .op(n10047) );
  or2_1 U11907 ( .ip1(n10047), .ip2(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .op(
        n10048) );
  nand2_1 U11908 ( .ip1(n10049), .ip2(n10048), .op(n10053) );
  nand3_1 U11909 ( .ip1(n11693), .ip2(n12656), .ip3(n11208), .op(n10051) );
  nand2_1 U11910 ( .ip1(n11782), .ip2(n5639), .op(n12625) );
  or2_1 U11911 ( .ip1(n10671), .ip2(n12625), .op(n10050) );
  nand2_1 U11912 ( .ip1(n10051), .ip2(n10050), .op(n10427) );
  and3_1 U11913 ( .ip1(n10057), .ip2(n10056), .ip3(n10055), .op(
        \CORTEXM0DS_INST/u_logic/N4396 ) );
  inv_1 U11914 ( .ip(n10058), .op(n11525) );
  nand2_1 U11915 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(n11525), .op(
        \CORTEXM0DS_INST/u_logic/N4359 ) );
  nand2_1 U11916 ( .ip1(n12664), .ip2(n11525), .op(n5998) );
  inv_1 U11917 ( .ip(n10076), .op(n10075) );
  inv_1 U11918 ( .ip(n12683), .op(n12684) );
  nor2_1 U11919 ( .ip1(n11455), .ip2(n12684), .op(n10060) );
  inv_1 U11920 ( .ip(n5998), .op(n10059) );
  not_ab_or_c_or_d U11921 ( .ip1(n10075), .ip2(n12661), .ip3(n10060), .ip4(
        n10059), .op(\CORTEXM0DS_INST/u_logic/N4282 ) );
  nand2_1 U11922 ( .ip1(n12664), .ip2(n12673), .op(n5996) );
  nor2_1 U11923 ( .ip1(n11462), .ip2(n12684), .op(n10062) );
  inv_1 U11924 ( .ip(n5996), .op(n10061) );
  not_ab_or_c_or_d U11925 ( .ip1(n10075), .ip2(n12662), .ip3(n10062), .ip4(
        n10061), .op(\CORTEXM0DS_INST/u_logic/N4227 ) );
  nand2_1 U11926 ( .ip1(n12664), .ip2(n12671), .op(n5994) );
  inv_1 U11927 ( .ip(n10063), .op(n12663) );
  nor2_1 U11928 ( .ip1(n11477), .ip2(n12684), .op(n10065) );
  inv_1 U11929 ( .ip(n5994), .op(n10064) );
  not_ab_or_c_or_d U11930 ( .ip1(n10075), .ip2(n12663), .ip3(n10065), .ip4(
        n10064), .op(\CORTEXM0DS_INST/u_logic/N4170 ) );
  nand2_1 U11931 ( .ip1(n12664), .ip2(n12677), .op(n5992) );
  inv_1 U11932 ( .ip(n10066), .op(n11484) );
  nor2_1 U11933 ( .ip1(n12665), .ip2(n10076), .op(n10068) );
  inv_1 U11934 ( .ip(n5992), .op(n10067) );
  not_ab_or_c_or_d U11935 ( .ip1(n12683), .ip2(n11484), .ip3(n10068), .ip4(
        n10067), .op(\CORTEXM0DS_INST/u_logic/N4116 ) );
  nand2_1 U11936 ( .ip1(n12664), .ip2(n12679), .op(n5988) );
  nor2_1 U11937 ( .ip1(n11330), .ip2(n10076), .op(n10070) );
  inv_1 U11938 ( .ip(n5988), .op(n10069) );
  not_ab_or_c_or_d U11939 ( .ip1(n12683), .ip2(n11488), .ip3(n10070), .ip4(
        n10069), .op(\CORTEXM0DS_INST/u_logic/N4005 ) );
  nand2_1 U11940 ( .ip1(n12664), .ip2(n12685), .op(n5986) );
  inv_1 U11941 ( .ip(n10071), .op(n12669) );
  nor2_1 U11942 ( .ip1(n10072), .ip2(n12684), .op(n10074) );
  inv_1 U11943 ( .ip(n5986), .op(n10073) );
  not_ab_or_c_or_d U11944 ( .ip1(n10075), .ip2(n12669), .ip3(n10074), .ip4(
        n10073), .op(\CORTEXM0DS_INST/u_logic/N3967 ) );
  nand2_1 U11945 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(n12677), .op(
        \CORTEXM0DS_INST/u_logic/N3966 ) );
  nand2_1 U11946 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(n12681), .op(
        \CORTEXM0DS_INST/u_logic/N3946 ) );
  inv_1 U11947 ( .ip(n11671), .op(n10080) );
  nor2_1 U11948 ( .ip1(n11340), .ip2(n10076), .op(n10079) );
  inv_1 U11949 ( .ip(n12664), .op(n12668) );
  nor2_1 U11950 ( .ip1(n10077), .ip2(n12668), .op(n10078) );
  not_ab_or_c_or_d U11951 ( .ip1(n12683), .ip2(n10080), .ip3(n10079), .ip4(
        n10078), .op(\CORTEXM0DS_INST/u_logic/N3783 ) );
  nand2_1 U11952 ( .ip1(n10916), .ip2(n11401), .op(n10158) );
  nand2_1 U11953 ( .ip1(\CORTEXM0DS_INST/vis_pc [17]), .ip2(
        \CORTEXM0DS_INST/vis_pc [18]), .op(n10082) );
  nand3_1 U11954 ( .ip1(n12113), .ip2(n10081), .ip3(n10327), .op(n10309) );
  nor2_1 U11955 ( .ip1(n10082), .ip2(n10309), .op(n10431) );
  inv_1 U11956 ( .ip(\CORTEXM0DS_INST/vis_pc [19]), .op(n12251) );
  nand2_1 U11957 ( .ip1(\CORTEXM0DS_INST/u_logic/Qsgvx4 ), .ip2(n10246), .op(
        n10085) );
  nand2_1 U11958 ( .ip1(n11853), .ip2(n10083), .op(n10084) );
  nand4_1 U11959 ( .ip1(n4092), .ip2(n10259), .ip3(n10085), .ip4(n10084), .op(
        n10392) );
  inv_1 U11960 ( .ip(n10086), .op(n10096) );
  nor2_1 U11961 ( .ip1(n10088), .ip2(n10087), .op(n10095) );
  and2_1 U11962 ( .ip1(n10271), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [4]), 
        .op(n10090) );
  inv_1 U11963 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [4]), .op(n11740) );
  nor2_1 U11964 ( .ip1(n11740), .ip2(n11830), .op(n10089) );
  not_ab_or_c_or_d U11965 ( .ip1(n11829), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [4]), .ip3(n10090), .ip4(n10089), .op(
        n10093) );
  nand2_1 U11966 ( .ip1(n10278), .ip2(\CORTEXM0DS_INST/u_logic/Vogvx4 ), .op(
        n10092) );
  nand2_1 U11967 ( .ip1(n10270), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [4]), 
        .op(n10091) );
  nand4_1 U11968 ( .ip1(n4097), .ip2(n10093), .ip3(n10092), .ip4(n10091), .op(
        n10094) );
  not_ab_or_c_or_d U11969 ( .ip1(n10285), .ip2(n10096), .ip3(n10095), .ip4(
        n10094), .op(n10393) );
  nor2_1 U11970 ( .ip1(n10393), .ip2(n10586), .op(n10154) );
  mux2_1 U11971 ( .ip1(n10098), .ip2(n10097), .s(n10256), .op(n10099) );
  nand2_1 U11972 ( .ip1(n11853), .ip2(n10099), .op(n10102) );
  nand2_1 U11973 ( .ip1(n10270), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [20]), 
        .op(n10101) );
  nand2_1 U11974 ( .ip1(n10271), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [20]), 
        .op(n10100) );
  nand4_1 U11975 ( .ip1(n4106), .ip2(n10102), .ip3(n10101), .ip4(n10100), .op(
        n10396) );
  nand2_1 U11976 ( .ip1(n10439), .ip2(n10396), .op(n10152) );
  inv_1 U11977 ( .ip(n10103), .op(n10137) );
  inv_1 U11978 ( .ip(n10104), .op(n10136) );
  nor2_1 U11979 ( .ip1(n10105), .ip2(n10108), .op(n10106) );
  not_ab_or_c_or_d U11980 ( .ip1(n10108), .ip2(n10107), .ip3(n10114), .ip4(
        n10106), .op(n10110) );
  not_ab_or_c_or_d U11981 ( .ip1(n10112), .ip2(n10111), .ip3(n10110), .ip4(
        n10109), .op(n10134) );
  nand3_1 U11982 ( .ip1(n10115), .ip2(n10114), .ip3(n10113), .op(n10133) );
  nand3_1 U11983 ( .ip1(n10117), .ip2(n10122), .ip3(n10116), .op(n10126) );
  nand3_1 U11984 ( .ip1(n10120), .ip2(n10119), .ip3(n10118), .op(n10125) );
  nand3_1 U11985 ( .ip1(n10123), .ip2(n10122), .ip3(n10121), .op(n10124) );
  nand3_1 U11986 ( .ip1(n10126), .ip2(n10125), .ip3(n10124), .op(n10127) );
  not_ab_or_c_or_d U11987 ( .ip1(n10130), .ip2(n10129), .ip3(n10128), .ip4(
        n10127), .op(n10132) );
  not_ab_or_c_or_d U11988 ( .ip1(n10134), .ip2(n10133), .ip3(n10132), .ip4(
        n10131), .op(n10135) );
  not_ab_or_c_or_d U11989 ( .ip1(n10138), .ip2(n10137), .ip3(n10136), .ip4(
        n10135), .op(n10139) );
  nor2_1 U11990 ( .ip1(\CORTEXM0DS_INST/u_logic/Krgvx4 ), .ip2(n10139), .op(
        n10140) );
  nor2_1 U11991 ( .ip1(\CORTEXM0DS_INST/u_logic/Eqgvx4 ), .ip2(n10140), .op(
        n12462) );
  nor3_1 U11992 ( .ip1(n10142), .ip2(n10141), .ip3(n11660), .op(n10150) );
  inv_1 U11993 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [12]), .op(n11707) );
  nor2_1 U11994 ( .ip1(n11707), .ip2(n11830), .op(n10143) );
  or2_1 U11995 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [12]), .ip2(n10143), 
        .op(n10145) );
  or2_1 U11996 ( .ip1(n10270), .ip2(n10143), .op(n10144) );
  nand2_1 U11997 ( .ip1(n10145), .ip2(n10144), .op(n10148) );
  nand2_1 U11998 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [12]), .ip2(n11829), 
        .op(n10147) );
  nand2_1 U11999 ( .ip1(n10271), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [12]), 
        .op(n10146) );
  nand4_1 U12000 ( .ip1(n4087), .ip2(n10148), .ip3(n10147), .ip4(n10146), .op(
        n10149) );
  not_ab_or_c_or_d U12001 ( .ip1(n10246), .ip2(n12462), .ip3(n10150), .ip4(
        n10149), .op(n10334) );
  inv_1 U12002 ( .ip(n10334), .op(n10390) );
  nand2_1 U12003 ( .ip1(n10437), .ip2(n10390), .op(n10151) );
  nand2_1 U12004 ( .ip1(n10152), .ip2(n10151), .op(n10153) );
  not_ab_or_c_or_d U12005 ( .ip1(n10392), .ip2(n10441), .ip3(n10154), .ip4(
        n10153), .op(n11404) );
  nor2_1 U12006 ( .ip1(n11404), .ip2(n10912), .op(n10156) );
  nor3_1 U12007 ( .ip1(n10431), .ip2(n10901), .ip3(n12251), .op(n10155) );
  not_ab_or_c_or_d U12008 ( .ip1(n10431), .ip2(n12251), .ip3(n10156), .ip4(
        n10155), .op(n10157) );
  nand3_1 U12009 ( .ip1(n10158), .ip2(n10157), .ip3(n10322), .op(
        \CORTEXM0DS_INST/u_logic/Ldhvx4 ) );
  inv_1 U12010 ( .ip(n4130), .op(n10448) );
  nand2_1 U12011 ( .ip1(n10448), .ip2(n10364), .op(n10161) );
  inv_1 U12012 ( .ip(n4149), .op(n10171) );
  nand2_1 U12013 ( .ip1(n10171), .ip2(n10361), .op(n10160) );
  nand2_1 U12014 ( .ip1(n10454), .ip2(n10370), .op(n10159) );
  nand3_1 U12015 ( .ip1(n10161), .ip2(n10160), .ip3(n10159), .op(n10162) );
  not_ab_or_c_or_d U12016 ( .ip1(n10451), .ip2(n10362), .ip3(n10369), .ip4(
        n10162), .op(n11595) );
  nor2_1 U12017 ( .ip1(n11595), .ip2(n10912), .op(n10166) );
  not_ab_or_c_or_d U12018 ( .ip1(n11005), .ip2(n10164), .ip3(n10163), .ip4(
        n10901), .op(n10165) );
  not_ab_or_c_or_d U12019 ( .ip1(n10916), .ip2(n11579), .ip3(n10166), .ip4(
        n10165), .op(n10167) );
  nand2_1 U12020 ( .ip1(n10167), .ip2(n10917), .op(
        \CORTEXM0DS_INST/u_logic/Sdhvx4 ) );
  nand3_1 U12021 ( .ip1(n12113), .ip2(n10168), .ip3(n10327), .op(n10465) );
  inv_1 U12022 ( .ip(n10465), .op(n10289) );
  not_ab_or_c_or_d U12023 ( .ip1(n12144), .ip2(n10169), .ip3(n10289), .ip4(
        n10901), .op(n10170) );
  inv_1 U12024 ( .ip(n10322), .op(n10433) );
  not_ab_or_c_or_d U12025 ( .ip1(n10916), .ip2(n12148), .ip3(n10170), .ip4(
        n10433), .op(n10177) );
  nand2_1 U12026 ( .ip1(n10448), .ip2(n10441), .op(n10175) );
  nand2_1 U12027 ( .ip1(n10452), .ip2(n10171), .op(n10174) );
  nand2_1 U12028 ( .ip1(n10454), .ip2(n10439), .op(n10173) );
  nand2_1 U12029 ( .ip1(n10451), .ip2(n10437), .op(n10172) );
  nand4_1 U12030 ( .ip1(n10175), .ip2(n10174), .ip3(n10173), .ip4(n10172), 
        .op(n11573) );
  nand2_1 U12031 ( .ip1(n10475), .ip2(n11573), .op(n10176) );
  nand2_1 U12032 ( .ip1(n10177), .ip2(n10176), .op(
        \CORTEXM0DS_INST/u_logic/Zdhvx4 ) );
  nor2_1 U12033 ( .ip1(\CORTEXM0DS_INST/vis_pc [20]), .ip2(n10179), .op(n10178) );
  not_ab_or_c_or_d U12034 ( .ip1(\CORTEXM0DS_INST/vis_pc [20]), .ip2(n10179), 
        .ip3(n10178), .ip4(n10901), .op(n10186) );
  inv_1 U12035 ( .ip(n10187), .op(n10378) );
  nor2_1 U12036 ( .ip1(n10375), .ip2(n10314), .op(n10183) );
  nand2_1 U12037 ( .ip1(n10439), .ip2(n10379), .op(n10181) );
  nand2_1 U12038 ( .ip1(n10441), .ip2(n10374), .op(n10180) );
  nand2_1 U12039 ( .ip1(n10181), .ip2(n10180), .op(n10182) );
  not_ab_or_c_or_d U12040 ( .ip1(n10452), .ip2(n10378), .ip3(n10183), .ip4(
        n10182), .op(n11417) );
  nor2_1 U12041 ( .ip1(n11417), .ip2(n10912), .op(n10185) );
  nor2_1 U12042 ( .ip1(n12263), .ip2(n10383), .op(n10184) );
  or4_1 U12043 ( .ip1(n10186), .ip2(n10185), .ip3(n10184), .ip4(n10433), .op(
        \CORTEXM0DS_INST/u_logic/Gehvx4 ) );
  nand2_1 U12044 ( .ip1(n10364), .ip2(n10374), .op(n10191) );
  nor2_1 U12045 ( .ip1(n10187), .ip2(n10350), .op(n10189) );
  nor2_1 U12046 ( .ip1(n10375), .ip2(n10351), .op(n10188) );
  not_ab_or_c_or_d U12047 ( .ip1(n10379), .ip2(n10370), .ip3(n10189), .ip4(
        n10188), .op(n10190) );
  inv_1 U12048 ( .ip(n10369), .op(n10354) );
  nand3_1 U12049 ( .ip1(n10191), .ip2(n10190), .ip3(n10354), .op(n11335) );
  nand2_1 U12050 ( .ip1(n10475), .ip2(n11335), .op(n10199) );
  nor2_1 U12051 ( .ip1(n10193), .ip2(n10192), .op(n10339) );
  nor2_1 U12052 ( .ip1(n10194), .ip2(n10383), .op(n10196) );
  nor3_1 U12053 ( .ip1(n10339), .ip2(n10901), .ip3(n10197), .op(n10195) );
  not_ab_or_c_or_d U12054 ( .ip1(n10339), .ip2(n10197), .ip3(n10196), .ip4(
        n10195), .op(n10198) );
  nand3_1 U12055 ( .ip1(n10199), .ip2(n10198), .ip3(n10917), .op(
        \CORTEXM0DS_INST/u_logic/Nehvx4 ) );
  nand2_1 U12056 ( .ip1(n10200), .ip2(n11786), .op(n10585) );
  nand2_1 U12057 ( .ip1(n10585), .ip2(n10201), .op(n11081) );
  not_ab_or_c_or_d U12058 ( .ip1(n10203), .ip2(n11782), .ip3(n10202), .ip4(
        n11081), .op(n12106) );
  nor2_1 U12059 ( .ip1(n12106), .ip2(n10204), .op(n10217) );
  inv_1 U12060 ( .ip(n10205), .op(n10626) );
  nand2_1 U12061 ( .ip1(n10647), .ip2(n10818), .op(n12090) );
  mux2_1 U12062 ( .ip1(n10218), .ip2(n12090), .s(n10206), .op(n11106) );
  inv_1 U12063 ( .ip(n11106), .op(n10207) );
  not_ab_or_c_or_d U12064 ( .ip1(n11181), .ip2(n10626), .ip3(n10732), .ip4(
        n10207), .op(n10219) );
  or2_1 U12065 ( .ip1(n10219), .ip2(n12571), .op(n10210) );
  nand3_1 U12066 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n10818), .ip3(
        n11090), .op(n10208) );
  or2_1 U12067 ( .ip1(n10208), .ip2(n12571), .op(n10209) );
  nand2_1 U12068 ( .ip1(n10210), .ip2(n10209), .op(n10212) );
  or2_1 U12069 ( .ip1(\CORTEXM0DS_INST/u_logic/K79vx4 ), .ip2(n10212), .op(
        n10214) );
  nand2_1 U12070 ( .ip1(n11101), .ip2(n11146), .op(n10211) );
  nand2_1 U12071 ( .ip1(n10572), .ip2(n10211), .op(n12094) );
  or2_1 U12072 ( .ip1(n12094), .ip2(n10212), .op(n10213) );
  nand2_1 U12073 ( .ip1(n10214), .ip2(n10213), .op(n10215) );
  nor2_1 U12074 ( .ip1(n10215), .ip2(n5772), .op(n10216) );
  ab_or_c_or_d U12075 ( .ip1(n5772), .ip2(\CORTEXM0DS_INST/u_logic/Ks9vx4 ), 
        .ip3(n10217), .ip4(n10216), .op(\CORTEXM0DS_INST/u_logic/Wfhvx4 ) );
  nand2_1 U12076 ( .ip1(n10219), .ip2(n10218), .op(n12101) );
  nand2_1 U12077 ( .ip1(\CORTEXM0DS_INST/u_logic/K79vx4 ), .ip2(n12101), .op(
        n10220) );
  or2_1 U12078 ( .ip1(n10220), .ip2(n5772), .op(n10223) );
  nand2_1 U12079 ( .ip1(\CORTEXM0DS_INST/u_logic/D69vx4 ), .ip2(n12094), .op(
        n10221) );
  or2_1 U12080 ( .ip1(n10221), .ip2(n5772), .op(n10222) );
  nand2_1 U12081 ( .ip1(n10223), .ip2(n10222), .op(n10226) );
  nor2_1 U12082 ( .ip1(n12106), .ip2(n10224), .op(n10225) );
  ab_or_c_or_d U12083 ( .ip1(n5772), .ip2(\CORTEXM0DS_INST/u_logic/Gr9vx4 ), 
        .ip3(n10226), .ip4(n10225), .op(\CORTEXM0DS_INST/u_logic/Dghvx4 ) );
  nor2_1 U12084 ( .ip1(n10589), .ip2(n10393), .op(n10228) );
  nor2_1 U12085 ( .ip1(n10334), .ip2(n10586), .op(n10227) );
  ab_or_c_or_d U12086 ( .ip1(n10593), .ip2(n10396), .ip3(n10228), .ip4(n10227), 
        .op(n10229) );
  not_ab_or_c_or_d U12087 ( .ip1(n10597), .ip2(n10392), .ip3(n10595), .ip4(
        n10229), .op(n11511) );
  nor2_1 U12088 ( .ip1(n11511), .ip2(n10912), .op(n10235) );
  not_ab_or_c_or_d U12089 ( .ip1(n10231), .ip2(n10240), .ip3(n10230), .ip4(
        n10901), .op(n10234) );
  nor2_1 U12090 ( .ip1(n10232), .ip2(n10383), .op(n10233) );
  or4_1 U12091 ( .ip1(n10467), .ip2(n10235), .ip3(n10234), .ip4(n10233), .op(
        \CORTEXM0DS_INST/u_logic/Thhvx4 ) );
  nor2_1 U12092 ( .ip1(n10589), .ip2(n10435), .op(n10239) );
  nand2_1 U12093 ( .ip1(n10436), .ip2(n10452), .op(n10237) );
  nand2_1 U12094 ( .ip1(n10593), .ip2(n10438), .op(n10236) );
  inv_1 U12095 ( .ip(n10595), .op(n10472) );
  nand3_1 U12096 ( .ip1(n10237), .ip2(n10236), .ip3(n10472), .op(n10238) );
  not_ab_or_c_or_d U12097 ( .ip1(n10597), .ip2(n10440), .ip3(n10239), .ip4(
        n10238), .op(n11487) );
  nor2_1 U12098 ( .ip1(n11487), .ip2(n10912), .op(n10245) );
  inv_1 U12099 ( .ip(n10290), .op(n10242) );
  inv_1 U12100 ( .ip(n10240), .op(n10241) );
  not_ab_or_c_or_d U12101 ( .ip1(n12309), .ip2(n10242), .ip3(n10241), .ip4(
        n10901), .op(n10244) );
  nor2_1 U12102 ( .ip1(n12312), .ip2(n10383), .op(n10243) );
  or4_1 U12103 ( .ip1(n10467), .ip2(n10245), .ip3(n10244), .ip4(n10243), .op(
        \CORTEXM0DS_INST/u_logic/Aihvx4 ) );
  nand2_1 U12104 ( .ip1(\CORTEXM0DS_INST/u_logic/R3hvx4 ), .ip2(n10246), .op(
        n10252) );
  nand2_1 U12105 ( .ip1(n10248), .ip2(n10247), .op(n10251) );
  nand2_1 U12106 ( .ip1(n10249), .ip2(n11853), .op(n10250) );
  nand4_1 U12107 ( .ip1(n4227), .ip2(n10252), .ip3(n10251), .ip4(n10250), .op(
        n10405) );
  nor2_1 U12108 ( .ip1(n10253), .ip2(n10256), .op(n10254) );
  not_ab_or_c_or_d U12109 ( .ip1(n10256), .ip2(n10255), .ip3(n10254), .ip4(
        n11660), .op(n10257) );
  not_ab_or_c_or_d U12110 ( .ip1(n10270), .ip2(
        \CORTEXM0DS_INST/u_logic/Czh2z4 [18]), .ip3(n4241), .ip4(n10257), .op(
        n10260) );
  nand2_1 U12111 ( .ip1(n10271), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [18]), 
        .op(n10258) );
  nand4_1 U12112 ( .ip1(n4243), .ip2(n10260), .ip3(n10259), .ip4(n10258), .op(
        n10411) );
  nand2_1 U12113 ( .ip1(n11829), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [10]), 
        .op(n10262) );
  nand2_1 U12114 ( .ip1(n10272), .ip2(\CORTEXM0DS_INST/u_logic/T1i2z4 [10]), 
        .op(n10261) );
  nand2_1 U12115 ( .ip1(n10262), .ip2(n10261), .op(n10268) );
  nand2_1 U12116 ( .ip1(n10285), .ip2(n10263), .op(n10266) );
  nand2_1 U12117 ( .ip1(n10271), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [10]), 
        .op(n10265) );
  nand2_1 U12118 ( .ip1(n10270), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [10]), 
        .op(n10264) );
  nand4_1 U12119 ( .ip1(n4237), .ip2(n10266), .ip3(n10265), .ip4(n10264), .op(
        n10267) );
  not_ab_or_c_or_d U12120 ( .ip1(n11645), .ip2(n10269), .ip3(n10268), .ip4(
        n10267), .op(n10406) );
  nor2_1 U12121 ( .ip1(n10406), .ip2(n10586), .op(n10287) );
  nand2_1 U12122 ( .ip1(n10270), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [2]), 
        .op(n10276) );
  nand2_1 U12123 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [2]), .ip2(n11829), 
        .op(n10275) );
  nand2_1 U12124 ( .ip1(n10271), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [2]), 
        .op(n10274) );
  nand2_1 U12125 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [2]), .ip2(n10272), 
        .op(n10273) );
  nand4_1 U12126 ( .ip1(n10276), .ip2(n10275), .ip3(n10274), .ip4(n10273), 
        .op(n10283) );
  nand2_1 U12127 ( .ip1(n11645), .ip2(n10277), .op(n10280) );
  nand2_1 U12128 ( .ip1(n10278), .ip2(\CORTEXM0DS_INST/u_logic/Nngvx4 ), .op(
        n10279) );
  nand4_1 U12129 ( .ip1(n4263), .ip2(n10281), .ip3(n10280), .ip4(n10279), .op(
        n10282) );
  not_ab_or_c_or_d U12130 ( .ip1(n10285), .ip2(n10284), .ip3(n10283), .ip4(
        n10282), .op(n10407) );
  nor2_1 U12131 ( .ip1(n10589), .ip2(n10407), .op(n10286) );
  ab_or_c_or_d U12132 ( .ip1(n10593), .ip2(n10411), .ip3(n10287), .ip4(n10286), 
        .op(n10288) );
  not_ab_or_c_or_d U12133 ( .ip1(n10597), .ip2(n10405), .ip3(n10595), .ip4(
        n10288), .op(n11482) );
  nor2_1 U12134 ( .ip1(n11482), .ip2(n10912), .op(n10295) );
  inv_1 U12135 ( .ip(\CORTEXM0DS_INST/vis_pc [25]), .op(n10292) );
  nand3_1 U12136 ( .ip1(\CORTEXM0DS_INST/vis_pc [23]), .ip2(
        \CORTEXM0DS_INST/vis_pc [24]), .ip3(n10289), .op(n10291) );
  not_ab_or_c_or_d U12137 ( .ip1(n10292), .ip2(n10291), .ip3(n10290), .ip4(
        n10901), .op(n10294) );
  nor2_1 U12138 ( .ip1(n12301), .ip2(n10383), .op(n10293) );
  or4_1 U12139 ( .ip1(n10467), .ip2(n10295), .ip3(n10294), .ip4(n10293), .op(
        \CORTEXM0DS_INST/u_logic/Hihvx4 ) );
  nor2_1 U12140 ( .ip1(n12345), .ip2(n10465), .op(n10464) );
  inv_1 U12141 ( .ip(\CORTEXM0DS_INST/vis_pc [24]), .op(n12289) );
  inv_1 U12142 ( .ip(n10589), .op(n10469) );
  nor2_1 U12143 ( .ip1(n10903), .ip2(n10586), .op(n10299) );
  nand2_1 U12144 ( .ip1(n10597), .ip2(n10905), .op(n10297) );
  nand2_1 U12145 ( .ip1(n10593), .ip2(n10911), .op(n10296) );
  nand3_1 U12146 ( .ip1(n10297), .ip2(n10296), .ip3(n10472), .op(n10298) );
  not_ab_or_c_or_d U12147 ( .ip1(n10469), .ip2(n10904), .ip3(n10299), .ip4(
        n10298), .op(n11469) );
  nor2_1 U12148 ( .ip1(n11469), .ip2(n10912), .op(n10301) );
  nor3_1 U12149 ( .ip1(n10464), .ip2(n10901), .ip3(n12289), .op(n10300) );
  not_ab_or_c_or_d U12150 ( .ip1(n10464), .ip2(n12289), .ip3(n10301), .ip4(
        n10300), .op(n10303) );
  or2_1 U12151 ( .ip1(n10383), .ip2(n12291), .op(n10302) );
  nand3_1 U12152 ( .ip1(n10303), .ip2(n10302), .ip3(n10917), .op(
        \CORTEXM0DS_INST/u_logic/Oihvx4 ) );
  nor2_1 U12153 ( .ip1(n10407), .ip2(n10586), .op(n10305) );
  nor2_1 U12154 ( .ip1(n10314), .ip2(n10406), .op(n10304) );
  not_ab_or_c_or_d U12155 ( .ip1(n10441), .ip2(n10405), .ip3(n10305), .ip4(
        n10304), .op(n10307) );
  nand2_1 U12156 ( .ip1(n10439), .ip2(n10411), .op(n10306) );
  nand2_1 U12157 ( .ip1(n10307), .ip2(n10306), .op(n11377) );
  nor2_1 U12158 ( .ip1(n12232), .ip2(n10383), .op(n10308) );
  not_ab_or_c_or_d U12159 ( .ip1(n10475), .ip2(n11377), .ip3(n10308), .ip4(
        n10433), .op(n10312) );
  inv_1 U12160 ( .ip(\CORTEXM0DS_INST/vis_pc [17]), .op(n12231) );
  inv_1 U12161 ( .ip(n10309), .op(n10430) );
  nand2_1 U12162 ( .ip1(n12231), .ip2(n10430), .op(n10311) );
  nand3_1 U12163 ( .ip1(\CORTEXM0DS_INST/vis_pc [17]), .ip2(n10309), .ip3(
        n12113), .op(n10310) );
  nand3_1 U12164 ( .ip1(n10312), .ip2(n10311), .ip3(n10310), .op(
        \CORTEXM0DS_INST/u_logic/Cjhvx4 ) );
  not_ab_or_c_or_d U12165 ( .ip1(n12220), .ip2(n10313), .ip3(n10430), .ip4(
        n10901), .op(n10320) );
  nor2_1 U12166 ( .ip1(n10314), .ip2(n10903), .op(n10318) );
  nand2_1 U12167 ( .ip1(n10911), .ip2(n10439), .op(n10316) );
  nand2_1 U12168 ( .ip1(n10452), .ip2(n10904), .op(n10315) );
  nand2_1 U12169 ( .ip1(n10316), .ip2(n10315), .op(n10317) );
  not_ab_or_c_or_d U12170 ( .ip1(n10441), .ip2(n10905), .ip3(n10318), .ip4(
        n10317), .op(n11372) );
  nor2_1 U12171 ( .ip1(n11372), .ip2(n10912), .op(n10319) );
  not_ab_or_c_or_d U12172 ( .ip1(n10916), .ip2(n11370), .ip3(n10320), .ip4(
        n10319), .op(n10321) );
  nand2_1 U12173 ( .ip1(n10322), .ip2(n10321), .op(
        \CORTEXM0DS_INST/u_logic/Jjhvx4 ) );
  nand2_1 U12174 ( .ip1(n10364), .ip2(n10596), .op(n10326) );
  nor2_1 U12175 ( .ip1(n10588), .ip2(n10350), .op(n10324) );
  nor2_1 U12176 ( .ip1(n10587), .ip2(n10351), .op(n10323) );
  not_ab_or_c_or_d U12177 ( .ip1(n10592), .ip2(n10370), .ip3(n10324), .ip4(
        n10323), .op(n10325) );
  nand3_1 U12178 ( .ip1(n10326), .ip2(n10325), .ip3(n10354), .op(n11345) );
  nand2_1 U12179 ( .ip1(\CORTEXM0DS_INST/vis_pc [12]), .ip2(n10339), .op(
        n10328) );
  not_ab_or_c_or_d U12180 ( .ip1(n10329), .ip2(n10328), .ip3(n10327), .ip4(
        n10901), .op(n10332) );
  nor2_1 U12181 ( .ip1(n10330), .ip2(n10383), .op(n10331) );
  not_ab_or_c_or_d U12182 ( .ip1(n10475), .ip2(n11345), .ip3(n10332), .ip4(
        n10331), .op(n10333) );
  nand2_1 U12183 ( .ip1(n10333), .ip2(n10917), .op(
        \CORTEXM0DS_INST/u_logic/Xjhvx4 ) );
  nor2_1 U12184 ( .ip1(n10393), .ip2(n10350), .op(n10336) );
  nor2_1 U12185 ( .ip1(n10334), .ip2(n10351), .op(n10335) );
  ab_or_c_or_d U12186 ( .ip1(n10396), .ip2(n10370), .ip3(n10336), .ip4(n10335), 
        .op(n10337) );
  not_ab_or_c_or_d U12187 ( .ip1(n10392), .ip2(n10364), .ip3(n10369), .ip4(
        n10337), .op(n11329) );
  nor2_1 U12188 ( .ip1(n11329), .ip2(n10912), .op(n10342) );
  inv_1 U12189 ( .ip(\CORTEXM0DS_INST/vis_pc [11]), .op(n12197) );
  nand2_1 U12190 ( .ip1(\CORTEXM0DS_INST/vis_pc [10]), .ip2(n10338), .op(
        n10340) );
  not_ab_or_c_or_d U12191 ( .ip1(n12197), .ip2(n10340), .ip3(n10339), .ip4(
        n10901), .op(n10341) );
  not_ab_or_c_or_d U12192 ( .ip1(n10916), .ip2(n11326), .ip3(n10342), .ip4(
        n10341), .op(n10343) );
  nand2_1 U12193 ( .ip1(n10343), .ip2(n10917), .op(
        \CORTEXM0DS_INST/u_logic/Ekhvx4 ) );
  inv_1 U12194 ( .ip(\CORTEXM0DS_INST/vis_pc [9]), .op(n12176) );
  or2_1 U12195 ( .ip1(n12176), .ip2(n10345), .op(n10348) );
  inv_1 U12196 ( .ip(n10344), .op(n10359) );
  nand2_1 U12197 ( .ip1(\CORTEXM0DS_INST/vis_pc [8]), .ip2(n10359), .op(n10346) );
  or2_1 U12198 ( .ip1(n10346), .ip2(n10345), .op(n10347) );
  nand2_1 U12199 ( .ip1(n10348), .ip2(n10347), .op(n10349) );
  not_ab_or_c_or_d U12200 ( .ip1(n12180), .ip2(n10916), .ip3(n10467), .ip4(
        n10349), .op(n10358) );
  nand2_1 U12201 ( .ip1(n10405), .ip2(n10364), .op(n10356) );
  nor2_1 U12202 ( .ip1(n10350), .ip2(n10407), .op(n10353) );
  nor2_1 U12203 ( .ip1(n10351), .ip2(n10406), .op(n10352) );
  not_ab_or_c_or_d U12204 ( .ip1(n10370), .ip2(n10411), .ip3(n10353), .ip4(
        n10352), .op(n10355) );
  nand3_1 U12205 ( .ip1(n10356), .ip2(n10355), .ip3(n10354), .op(n11302) );
  nand2_1 U12206 ( .ip1(n10475), .ip2(n11302), .op(n10357) );
  nand2_1 U12207 ( .ip1(n10358), .ip2(n10357), .op(
        \CORTEXM0DS_INST/u_logic/Lkhvx4 ) );
  inv_1 U12208 ( .ip(n12155), .op(n11556) );
  not_ab_or_c_or_d U12209 ( .ip1(n12154), .ip2(n10360), .ip3(n10359), .ip4(
        n10901), .op(n10372) );
  nand2_1 U12210 ( .ip1(n11044), .ip2(n10361), .op(n10367) );
  nand2_1 U12211 ( .ip1(n10363), .ip2(n10362), .op(n10366) );
  nand2_1 U12212 ( .ip1(n10468), .ip2(n10364), .op(n10365) );
  nand3_1 U12213 ( .ip1(n10367), .ip2(n10366), .ip3(n10365), .op(n10368) );
  not_ab_or_c_or_d U12214 ( .ip1(n11036), .ip2(n10370), .ip3(n10369), .ip4(
        n10368), .op(n11567) );
  nor2_1 U12215 ( .ip1(n11567), .ip2(n10912), .op(n10371) );
  not_ab_or_c_or_d U12216 ( .ip1(n10916), .ip2(n11556), .ip3(n10372), .ip4(
        n10371), .op(n10373) );
  nand2_1 U12217 ( .ip1(n10373), .ip2(n10917), .op(
        \CORTEXM0DS_INST/u_logic/Skhvx4 ) );
  nand2_1 U12218 ( .ip1(n10906), .ip2(n10374), .op(n10382) );
  nor2_1 U12219 ( .ip1(n10375), .ip2(n11038), .op(n10377) );
  not_ab_or_c_or_d U12220 ( .ip1(n10378), .ip2(n11043), .ip3(n10377), .ip4(
        n10376), .op(n10381) );
  nand2_1 U12221 ( .ip1(n10379), .ip2(n11037), .op(n10380) );
  nand3_1 U12222 ( .ip1(n10382), .ip2(n10381), .ip3(n10380), .op(n11442) );
  nor2_1 U12223 ( .ip1(n10384), .ip2(n10383), .op(n10388) );
  nor2_1 U12224 ( .ip1(n10401), .ip2(n10400), .op(n10399) );
  nor2_1 U12225 ( .ip1(\CORTEXM0DS_INST/vis_pc [4]), .ip2(n10399), .op(n10386)
         );
  nor3_1 U12226 ( .ip1(n10386), .ip2(n10385), .ip3(n10901), .op(n10387) );
  not_ab_or_c_or_d U12227 ( .ip1(n10475), .ip2(n11442), .ip3(n10388), .ip4(
        n10387), .op(n10389) );
  nand2_1 U12228 ( .ip1(n10389), .ip2(n10917), .op(
        \CORTEXM0DS_INST/u_logic/Nlhvx4 ) );
  nand2_1 U12229 ( .ip1(n10391), .ip2(n10390), .op(n10398) );
  and2_1 U12230 ( .ip1(n10392), .ip2(n10906), .op(n10395) );
  nor2_1 U12231 ( .ip1(n10393), .ip2(n10408), .op(n10394) );
  not_ab_or_c_or_d U12232 ( .ip1(n10396), .ip2(n11037), .ip3(n10395), .ip4(
        n10394), .op(n10397) );
  nand3_1 U12233 ( .ip1(n10398), .ip2(n10397), .ip3(n11045), .op(n11435) );
  not_ab_or_c_or_d U12234 ( .ip1(n10401), .ip2(n10400), .ip3(n10399), .ip4(
        n10901), .op(n10402) );
  not_ab_or_c_or_d U12235 ( .ip1(n10475), .ip2(n11435), .ip3(n10467), .ip4(
        n10402), .op(n10404) );
  nand2_1 U12236 ( .ip1(n11437), .ip2(n10916), .op(n10403) );
  nand2_1 U12237 ( .ip1(n10404), .ip2(n10403), .op(
        \CORTEXM0DS_INST/u_logic/Ulhvx4 ) );
  nand2_1 U12238 ( .ip1(n10405), .ip2(n10906), .op(n10413) );
  nor2_1 U12239 ( .ip1(n11038), .ip2(n10406), .op(n10410) );
  nor2_1 U12240 ( .ip1(n10408), .ip2(n10407), .op(n10409) );
  not_ab_or_c_or_d U12241 ( .ip1(n11037), .ip2(n10411), .ip3(n10410), .ip4(
        n10409), .op(n10412) );
  nand3_1 U12242 ( .ip1(n10413), .ip2(n10412), .ip3(n11045), .op(n11298) );
  nand2_1 U12243 ( .ip1(\CORTEXM0DS_INST/vis_pc [0]), .ip2(n10414), .op(n10416) );
  not_ab_or_c_or_d U12244 ( .ip1(n12401), .ip2(n10416), .ip3(n10415), .ip4(
        n10901), .op(n10417) );
  not_ab_or_c_or_d U12245 ( .ip1(n10475), .ip2(n11298), .ip3(n10467), .ip4(
        n10417), .op(n10420) );
  nand2_1 U12246 ( .ip1(n10418), .ip2(n10916), .op(n10419) );
  nand2_1 U12247 ( .ip1(n10420), .ip2(n10419), .op(
        \CORTEXM0DS_INST/u_logic/Imhvx4 ) );
  nor2_1 U12248 ( .ip1(n12609), .ip2(n11693), .op(n10429) );
  inv_1 U12249 ( .ip(n10740), .op(n12612) );
  nand3_1 U12250 ( .ip1(n12619), .ip2(n10421), .ip3(n12612), .op(n12615) );
  inv_1 U12251 ( .ip(n12615), .op(n10428) );
  nand3_1 U12252 ( .ip1(n11267), .ip2(n12624), .ip3(n12623), .op(n10564) );
  nand2_1 U12253 ( .ip1(n12610), .ip2(n12612), .op(n10423) );
  ab_or_c_or_d U12254 ( .ip1(n12118), .ip2(n10423), .ip3(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip4(n10422), .op(n10424) );
  nand3_1 U12255 ( .ip1(n10425), .ip2(n10564), .ip3(n10424), .op(n10426) );
  not_ab_or_c_or_d U12256 ( .ip1(n10429), .ip2(n10428), .ip3(n10427), .ip4(
        n10426), .op(\CORTEXM0DS_INST/u_logic/N2678 ) );
  inv_1 U12257 ( .ip(\CORTEXM0DS_INST/vis_pc [18]), .op(n12243) );
  nand2_1 U12258 ( .ip1(\CORTEXM0DS_INST/vis_pc [17]), .ip2(n10430), .op(
        n10432) );
  not_ab_or_c_or_d U12259 ( .ip1(n12243), .ip2(n10432), .ip3(n10431), .ip4(
        n10901), .op(n10434) );
  not_ab_or_c_or_d U12260 ( .ip1(n10916), .ip2(n12246), .ip3(n10434), .ip4(
        n10433), .op(n10447) );
  or2_1 U12261 ( .ip1(n10586), .ip2(n10435), .op(n10445) );
  nand2_1 U12262 ( .ip1(n10437), .ip2(n10436), .op(n10444) );
  nand2_1 U12263 ( .ip1(n10439), .ip2(n10438), .op(n10443) );
  nand2_1 U12264 ( .ip1(n10441), .ip2(n10440), .op(n10442) );
  nand4_1 U12265 ( .ip1(n10445), .ip2(n10444), .ip3(n10443), .ip4(n10442), 
        .op(n11391) );
  nand2_1 U12266 ( .ip1(n10475), .ip2(n11391), .op(n10446) );
  nand2_1 U12267 ( .ip1(n10447), .ip2(n10446), .op(
        \CORTEXM0DS_INST/u_logic/Ithvx4 ) );
  and2_1 U12268 ( .ip1(n10448), .ip2(n10597), .op(n10450) );
  nor2_1 U12269 ( .ip1(n4149), .ip2(n10589), .op(n10449) );
  ab_or_c_or_d U12270 ( .ip1(n10452), .ip2(n10451), .ip3(n10450), .ip4(n10449), 
        .op(n10453) );
  not_ab_or_c_or_d U12271 ( .ip1(n10454), .ip2(n10593), .ip3(n10595), .ip4(
        n10453), .op(n11662) );
  nor2_1 U12272 ( .ip1(n11662), .ip2(n10912), .op(n10461) );
  nor4_1 U12273 ( .ip1(n10457), .ip2(n12309), .ip3(n10456), .ip4(n10455), .op(
        n10598) );
  nor2_1 U12274 ( .ip1(n10598), .ip2(\CORTEXM0DS_INST/vis_pc [30]), .op(n10458) );
  not_ab_or_c_or_d U12275 ( .ip1(n10598), .ip2(\CORTEXM0DS_INST/vis_pc [30]), 
        .ip3(n10458), .ip4(n10901), .op(n10459) );
  mux2_1 U12276 ( .ip1(n10459), .ip2(\CORTEXM0DS_INST/vis_pc [30]), .s(n5814), 
        .op(n10460) );
  not_ab_or_c_or_d U12277 ( .ip1(n10462), .ip2(n10916), .ip3(n10461), .ip4(
        n10460), .op(n10463) );
  nand2_1 U12278 ( .ip1(n10463), .ip2(n10917), .op(
        \CORTEXM0DS_INST/u_logic/Wthvx4 ) );
  not_ab_or_c_or_d U12279 ( .ip1(n12345), .ip2(n10465), .ip3(n10464), .ip4(
        n10901), .op(n10466) );
  not_ab_or_c_or_d U12280 ( .ip1(n12351), .ip2(n10916), .ip3(n10467), .ip4(
        n10466), .op(n10477) );
  nand2_1 U12281 ( .ip1(n10468), .ip2(n10597), .op(n10474) );
  nor2_1 U12282 ( .ip1(n4286), .ip2(n10586), .op(n10471) );
  and2_1 U12283 ( .ip1(n10469), .ip2(n11044), .op(n10470) );
  not_ab_or_c_or_d U12284 ( .ip1(n10593), .ip2(n11036), .ip3(n10471), .ip4(
        n10470), .op(n10473) );
  nand3_1 U12285 ( .ip1(n10474), .ip2(n10473), .ip3(n10472), .op(n11456) );
  nand2_1 U12286 ( .ip1(n10475), .ip2(n11456), .op(n10476) );
  nand2_1 U12287 ( .ip1(n10477), .ip2(n10476), .op(
        \CORTEXM0DS_INST/u_logic/Duhvx4 ) );
  nor2_1 U12288 ( .ip1(n5932), .ip2(n12118), .op(n12651) );
  nand3_1 U12289 ( .ip1(n11693), .ip2(n12651), .ip3(n10478), .op(n10529) );
  nand2_1 U12290 ( .ip1(n5932), .ip2(n11796), .op(n10527) );
  nor3_1 U12291 ( .ip1(n11011), .ip2(n12623), .ip3(n12117), .op(n10480) );
  nor2_1 U12292 ( .ip1(n10479), .ip2(n10779), .op(n10708) );
  nor3_1 U12293 ( .ip1(n11686), .ip2(n10480), .ip3(n10708), .op(n10525) );
  inv_1 U12294 ( .ip(n10481), .op(n10836) );
  nand2_1 U12295 ( .ip1(n10836), .ip2(n11102), .op(n10483) );
  nand2_1 U12296 ( .ip1(n10635), .ip2(n12583), .op(n10482) );
  not_ab_or_c_or_d U12297 ( .ip1(n10483), .ip2(n10482), .ip3(n12321), .ip4(
        n10542), .op(n10485) );
  nor2_1 U12298 ( .ip1(n10484), .ip2(n11788), .op(n12622) );
  not_ab_or_c_or_d U12299 ( .ip1(n10651), .ip2(n10635), .ip3(n10485), .ip4(
        n12622), .op(n10509) );
  nor3_1 U12300 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n12321), .ip3(
        n10486), .op(n10489) );
  nor2_1 U12301 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n10487), .op(
        n10488) );
  not_ab_or_c_or_d U12302 ( .ip1(n10490), .ip2(n10636), .ip3(n10489), .ip4(
        n10488), .op(n10508) );
  or2_1 U12303 ( .ip1(n10491), .ip2(n10542), .op(n10498) );
  nand3_1 U12304 ( .ip1(n10869), .ip2(n11107), .ip3(n10492), .op(n10723) );
  nor4_1 U12305 ( .ip1(\CORTEXM0DS_INST/u_logic/K79vx4 ), .ip2(n10494), .ip3(
        n12599), .ip4(n10493), .op(n10495) );
  nand3_1 U12306 ( .ip1(n10496), .ip2(n10651), .ip3(n10495), .op(n10497) );
  nand3_1 U12307 ( .ip1(n10498), .ip2(n10723), .ip3(n10497), .op(n10506) );
  not_ab_or_c_or_d U12308 ( .ip1(n10500), .ip2(n10979), .ip3(n10499), .ip4(
        n10492), .op(n10502) );
  nand2_1 U12309 ( .ip1(n10635), .ip2(n10551), .op(n10501) );
  not_ab_or_c_or_d U12310 ( .ip1(n10503), .ip2(n10502), .ip3(
        \CORTEXM0DS_INST/u_logic/Ho8vx4 ), .ip4(n10501), .op(n10505) );
  nor3_1 U12311 ( .ip1(n10892), .ip2(n10851), .ip3(n10671), .op(n10504) );
  not_ab_or_c_or_d U12312 ( .ip1(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip2(
        n10506), .ip3(n10505), .ip4(n10504), .op(n10507) );
  nand3_1 U12313 ( .ip1(n10509), .ip2(n10508), .ip3(n10507), .op(n10521) );
  nand4_1 U12314 ( .ip1(n12132), .ip2(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip3(
        n11796), .ip4(n10955), .op(n10669) );
  or2_1 U12315 ( .ip1(n10669), .ip2(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .op(
        n10511) );
  nand2_1 U12316 ( .ip1(\CORTEXM0DS_INST/u_logic/Ki8vx4 ), .ip2(n10863), .op(
        n10510) );
  nand2_1 U12317 ( .ip1(n10511), .ip2(n10510), .op(n10520) );
  nor4_1 U12318 ( .ip1(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip2(n10512), .ip3(
        n10706), .ip4(n10842), .op(n10513) );
  nor4_1 U12319 ( .ip1(n10516), .ip2(n10515), .ip3(n10514), .ip4(n10513), .op(
        n10518) );
  inv_1 U12320 ( .ip(n11802), .op(n10517) );
  nand4_1 U12321 ( .ip1(n10752), .ip2(n10518), .ip3(n10564), .ip4(n10517), 
        .op(n10519) );
  not_ab_or_c_or_d U12322 ( .ip1(n5639), .ip2(n10521), .ip3(n10520), .ip4(
        n10519), .op(n10524) );
  nand3_1 U12323 ( .ip1(n10764), .ip2(n12117), .ip3(n11786), .op(n10522) );
  nand4_1 U12324 ( .ip1(n10525), .ip2(n10524), .ip3(n10523), .ip4(n10522), 
        .op(n10526) );
  nand2_1 U12325 ( .ip1(n10527), .ip2(n10526), .op(n10528) );
  nand2_1 U12326 ( .ip1(n10529), .ip2(n10528), .op(
        \CORTEXM0DS_INST/u_logic/Yuhvx4 ) );
  nor3_1 U12327 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n12623), .ip3(
        n11228), .op(n10804) );
  nor2_1 U12328 ( .ip1(n10530), .ip2(n11786), .op(n10688) );
  inv_1 U12329 ( .ip(n10688), .op(n10560) );
  or2_1 U12330 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n10531), .op(
        n10532) );
  or2_1 U12331 ( .ip1(n10532), .ip2(n11277), .op(n10644) );
  or2_1 U12332 ( .ip1(n10533), .ip2(n11228), .op(n10534) );
  or2_1 U12333 ( .ip1(n10534), .ip2(n11277), .op(n10535) );
  nand2_1 U12334 ( .ip1(n10644), .ip2(n10535), .op(n10559) );
  nand2_1 U12335 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n10884), .op(
        n10537) );
  nand3_1 U12336 ( .ip1(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip2(n12583), .ip3(
        n12122), .op(n10536) );
  not_ab_or_c_or_d U12337 ( .ip1(n10537), .ip2(n10536), .ip3(n12592), .ip4(
        n9807), .op(n10538) );
  nor4_1 U12338 ( .ip1(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip3(n9807), .ip4(n11100), .op(
        n10874) );
  not_ab_or_c_or_d U12339 ( .ip1(n10933), .ip2(n10539), .ip3(n10538), .ip4(
        n10874), .op(n10554) );
  nand3_1 U12340 ( .ip1(n10492), .ip2(n10551), .ip3(
        \CORTEXM0DS_INST/u_logic/Kg9vx4 ), .op(n10541) );
  nand2_1 U12341 ( .ip1(n10541), .ip2(n10540), .op(n10545) );
  nor2_1 U12342 ( .ip1(n10542), .ip2(n12321), .op(n10544) );
  nor2_1 U12343 ( .ip1(n12538), .ip2(n10492), .op(n10622) );
  nor2_1 U12344 ( .ip1(n10622), .ip2(n11088), .op(n10543) );
  not_ab_or_c_or_d U12345 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(
        n10545), .ip3(n10544), .ip4(n10543), .op(n10553) );
  nand4_1 U12346 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/R89vx4 ), .ip3(n12588), .ip4(n10546), .op(
        n10549) );
  nand2_1 U12347 ( .ip1(n10713), .ip2(n12567), .op(n10548) );
  nand2_1 U12348 ( .ip1(n12588), .ip2(n10837), .op(n10719) );
  nand3_1 U12349 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n10719), .ip3(
        n10623), .op(n10547) );
  nand4_1 U12350 ( .ip1(n10635), .ip2(n10549), .ip3(n10548), .ip4(n10547), 
        .op(n10550) );
  nand4_1 U12351 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n10551), .ip3(
        n12122), .ip4(n10550), .op(n10552) );
  nand3_1 U12352 ( .ip1(n10554), .ip2(n10553), .ip3(n10552), .op(n10557) );
  ab_or_c_or_d U12353 ( .ip1(n5639), .ip2(n10557), .ip3(n10556), .ip4(n10555), 
        .op(n10558) );
  not_ab_or_c_or_d U12354 ( .ip1(n10804), .ip2(n10560), .ip3(n10559), .ip4(
        n10558), .op(n10561) );
  nor2_1 U12355 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n10561), .op(
        n10582) );
  nor4_1 U12356 ( .ip1(n10892), .ip2(n11786), .ip3(n10563), .ip4(n10562), .op(
        n10581) );
  nor3_1 U12357 ( .ip1(n10955), .ip2(n12627), .ip3(n10564), .op(n10580) );
  nor3_1 U12358 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip3(n11080), .op(n11757) );
  nand2_1 U12359 ( .ip1(n10786), .ip2(n11796), .op(n10934) );
  nor2_1 U12360 ( .ip1(n11243), .ip2(n10934), .op(n10565) );
  or2_1 U12361 ( .ip1(n11757), .ip2(n10565), .op(n10567) );
  or2_1 U12362 ( .ip1(n11250), .ip2(n10565), .op(n10566) );
  nand2_1 U12363 ( .ip1(n10567), .ip2(n10566), .op(n10578) );
  nor4_1 U12364 ( .ip1(n12126), .ip2(n11228), .ip3(n11231), .ip4(n10949), .op(
        n10951) );
  nor2_1 U12365 ( .ip1(n12609), .ip2(n10885), .op(n10816) );
  inv_1 U12366 ( .ip(n10816), .op(n10568) );
  or2_1 U12367 ( .ip1(n10568), .ip2(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .op(
        n10571) );
  or2_1 U12368 ( .ip1(n10569), .ip2(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .op(
        n10570) );
  nand2_1 U12369 ( .ip1(n10571), .ip2(n10570), .op(n10574) );
  not_ab_or_c_or_d U12370 ( .ip1(n10572), .ip2(n11105), .ip3(
        \CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip4(n12592), .op(n10573) );
  not_ab_or_c_or_d U12371 ( .ip1(n10951), .ip2(n11248), .ip3(n10574), .ip4(
        n10573), .op(n10577) );
  nor2_1 U12372 ( .ip1(n10610), .ip2(n10949), .op(n10731) );
  nand3_1 U12373 ( .ip1(n11250), .ip2(n10731), .ip3(n11796), .op(n10576) );
  nand2_1 U12374 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n11076), .op(
        n10575) );
  nand4_1 U12375 ( .ip1(n10578), .ip2(n10577), .ip3(n10576), .ip4(n10575), 
        .op(n10579) );
  nor4_1 U12376 ( .ip1(n10582), .ip2(n10581), .ip3(n10580), .ip4(n10579), .op(
        n10583) );
  inv_1 U12377 ( .ip(n5932), .op(n12648) );
  mux2_1 U12378 ( .ip1(n12609), .ip2(n10583), .s(n12648), .op(n10584) );
  nand2_1 U12379 ( .ip1(n10585), .ip2(n10584), .op(
        \CORTEXM0DS_INST/u_logic/Mvhvx4 ) );
  nor2_1 U12380 ( .ip1(n10587), .ip2(n10586), .op(n10591) );
  nor2_1 U12381 ( .ip1(n10589), .ip2(n10588), .op(n10590) );
  ab_or_c_or_d U12382 ( .ip1(n10593), .ip2(n10592), .ip3(n10591), .ip4(n10590), 
        .op(n10594) );
  not_ab_or_c_or_d U12383 ( .ip1(n10597), .ip2(n10596), .ip3(n10595), .ip4(
        n10594), .op(n11672) );
  nor2_1 U12384 ( .ip1(n11672), .ip2(n10912), .op(n10607) );
  inv_1 U12385 ( .ip(n10598), .op(n10599) );
  or2_1 U12386 ( .ip1(n10599), .ip2(n5814), .op(n10600) );
  nand2_1 U12387 ( .ip1(n12113), .ip2(n10600), .op(n10602) );
  or2_1 U12388 ( .ip1(n10601), .ip2(n10602), .op(n10605) );
  or2_1 U12389 ( .ip1(n10603), .ip2(n10602), .op(n10604) );
  nand2_1 U12390 ( .ip1(n10605), .ip2(n10604), .op(n10606) );
  not_ab_or_c_or_d U12391 ( .ip1(n10916), .ip2(n10608), .ip3(n10607), .ip4(
        n10606), .op(n10609) );
  nand2_1 U12392 ( .ip1(n10609), .ip2(n10917), .op(
        \CORTEXM0DS_INST/u_logic/Tvhvx4 ) );
  nand2_1 U12393 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n10610), .op(
        n11251) );
  and2_1 U12394 ( .ip1(n10611), .ip2(n11757), .op(n10618) );
  inv_1 U12395 ( .ip(n10612), .op(n11266) );
  not_ab_or_c_or_d U12396 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n5639), .ip3(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip4(n11789), .op(n10615) );
  nor2_1 U12397 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Q5gvx4 ), .op(n10613) );
  nor3_1 U12398 ( .ip1(n10613), .ip2(n11223), .ip3(n11796), .op(n10614) );
  not_ab_or_c_or_d U12399 ( .ip1(n11099), .ip2(n11266), .ip3(n10615), .ip4(
        n10614), .op(n10616) );
  nor2_1 U12400 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10616), .op(
        n10617) );
  not_ab_or_c_or_d U12401 ( .ip1(n10619), .ip2(n11251), .ip3(n10618), .ip4(
        n10617), .op(n10681) );
  not_ab_or_c_or_d U12402 ( .ip1(n10622), .ip2(n10621), .ip3(
        \CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip4(n10620), .op(n10630) );
  or3_1 U12403 ( .ip1(n12567), .ip2(n10624), .ip3(n10623), .op(n10629) );
  or2_1 U12404 ( .ip1(n10626), .ip2(n10625), .op(n10628) );
  nand3_1 U12405 ( .ip1(n10932), .ip2(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip3(
        n11100), .op(n10627) );
  nand4_1 U12406 ( .ip1(n10630), .ip2(n10629), .ip3(n10628), .ip4(n10627), 
        .op(n10640) );
  or2_1 U12407 ( .ip1(n12628), .ip2(n5639), .op(n10773) );
  or2_1 U12408 ( .ip1(n10773), .ip2(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .op(
        n10634) );
  nand3_1 U12409 ( .ip1(n10632), .ip2(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip3(
        n10631), .op(n10633) );
  nand2_1 U12410 ( .ip1(n10634), .ip2(n10633), .op(n10639) );
  nor2_1 U12411 ( .ip1(\CORTEXM0DS_INST/u_logic/R89vx4 ), .ip2(n12583), .op(
        n10859) );
  not_ab_or_c_or_d U12412 ( .ip1(n10859), .ip2(n12567), .ip3(n10636), .ip4(
        n10635), .op(n10637) );
  nor2_1 U12413 ( .ip1(n10637), .ip2(n12321), .op(n10638) );
  not_ab_or_c_or_d U12414 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(
        n10640), .ip3(n10639), .ip4(n10638), .op(n10668) );
  nor3_1 U12415 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(n12138), .ip3(
        n11228), .op(n10641) );
  not_ab_or_c_or_d U12416 ( .ip1(n10892), .ip2(n10642), .ip3(n11250), .ip4(
        n10641), .op(n10643) );
  nor3_1 U12417 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip3(n10643), .op(n10661) );
  or2_1 U12418 ( .ip1(n10971), .ip2(n11277), .op(n10645) );
  nand2_1 U12419 ( .ip1(n10645), .ip2(n10644), .op(n10660) );
  nor2_1 U12420 ( .ip1(n12599), .ip2(n10646), .op(n10769) );
  not_ab_or_c_or_d U12421 ( .ip1(n10647), .ip2(n10836), .ip3(n11107), .ip4(
        n10769), .op(n10648) );
  nor2_1 U12422 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(n10648), .op(
        n10659) );
  nor3_1 U12423 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n11100), .ip3(
        n10842), .op(n10649) );
  not_ab_or_c_or_d U12424 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(
        n11146), .ip3(n10650), .ip4(n10649), .op(n10657) );
  nand3_1 U12425 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n10651), .ip3(
        n12588), .op(n10656) );
  nor2_1 U12426 ( .ip1(n10932), .ip2(n10859), .op(n10721) );
  nand4_1 U12427 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip4(n10721), .op(n10655) );
  nand2_1 U12428 ( .ip1(n10653), .ip2(n10652), .op(n10654) );
  nand4_1 U12429 ( .ip1(n10657), .ip2(n10656), .ip3(n10655), .ip4(n10654), 
        .op(n10658) );
  nor4_1 U12430 ( .ip1(n10661), .ip2(n10660), .ip3(n10659), .ip4(n10658), .op(
        n10667) );
  nand3_1 U12431 ( .ip1(n10892), .ip2(n11256), .ip3(n10662), .op(n10666) );
  nand2_1 U12432 ( .ip1(n5092), .ip2(n10806), .op(n10663) );
  nand2_1 U12433 ( .ip1(n10664), .ip2(n10663), .op(n10665) );
  nand4_1 U12434 ( .ip1(n10668), .ip2(n10667), .ip3(n10666), .ip4(n10665), 
        .op(n10676) );
  nor2_1 U12435 ( .ip1(n11239), .ip2(n10669), .op(n10675) );
  inv_1 U12436 ( .ip(n10670), .op(n10672) );
  nor4_1 U12437 ( .ip1(n10851), .ip2(n10673), .ip3(n10672), .ip4(n10671), .op(
        n10674) );
  not_ab_or_c_or_d U12438 ( .ip1(n12125), .ip2(n10676), .ip3(n10675), .ip4(
        n10674), .op(n10680) );
  nand2_1 U12439 ( .ip1(n10677), .ip2(n10764), .op(n10678) );
  nand4_1 U12440 ( .ip1(n10681), .ip2(n10680), .ip3(n10679), .ip4(n10678), 
        .op(n10682) );
  mux2_1 U12441 ( .ip1(n10682), .ip2(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .s(
        n5932), .op(\CORTEXM0DS_INST/u_logic/Hwhvx4 ) );
  nor3_1 U12442 ( .ip1(\CORTEXM0DS_INST/u_logic/K79vx4 ), .ip2(n10683), .ip3(
        n10926), .op(n10686) );
  nor3_1 U12443 ( .ip1(n12592), .ip2(n12567), .ip3(n10978), .op(n10685) );
  nor2_1 U12444 ( .ip1(\CORTEXM0DS_INST/u_logic/R89vx4 ), .ip2(n10978), .op(
        n10684) );
  ab_or_c_or_d U12445 ( .ip1(n10686), .ip2(n12571), .ip3(n10685), .ip4(n10684), 
        .op(n10792) );
  nor2_1 U12446 ( .ip1(n12138), .ip2(n10687), .op(n10694) );
  not_ab_or_c_or_d U12447 ( .ip1(n10689), .ip2(n11703), .ip3(n10688), .ip4(
        n12625), .op(n10693) );
  nor2_1 U12448 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n10690), .op(
        n10692) );
  nor3_1 U12449 ( .ip1(n11796), .ip2(n11793), .ip3(n10782), .op(n10691) );
  nor4_1 U12450 ( .ip1(n10694), .ip2(n10693), .ip3(n10692), .ip4(n10691), .op(
        n10695) );
  or2_1 U12451 ( .ip1(n10695), .ip2(n10865), .op(n10704) );
  nor3_1 U12452 ( .ip1(n10698), .ip2(n10697), .ip3(n10696), .op(n10699) );
  or2_1 U12453 ( .ip1(n10699), .ip2(n10743), .op(n10700) );
  nand3_1 U12454 ( .ip1(n10701), .ip2(n10818), .ip3(n10700), .op(n10702) );
  or2_1 U12455 ( .ip1(n10702), .ip2(n10865), .op(n10703) );
  nand2_1 U12456 ( .ip1(n10704), .ip2(n10703), .op(n10791) );
  nor2_1 U12457 ( .ip1(n10706), .ip2(n10705), .op(n10707) );
  not_ab_or_c_or_d U12458 ( .ip1(n10804), .ip2(n11786), .ip3(n10708), .ip4(
        n10707), .op(n10709) );
  or2_1 U12459 ( .ip1(n10709), .ip2(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .op(
        n10712) );
  nand2_1 U12460 ( .ip1(n11249), .ip2(n12134), .op(n10710) );
  or2_1 U12461 ( .ip1(n10710), .ip2(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .op(
        n10711) );
  nand2_1 U12462 ( .ip1(n10712), .ip2(n10711), .op(n10757) );
  nand2_1 U12463 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n10713), .op(
        n10714) );
  nand2_1 U12464 ( .ip1(n10715), .ip2(n10714), .op(n10716) );
  nand2_1 U12465 ( .ip1(n10884), .ip2(n10716), .op(n10717) );
  nor3_1 U12466 ( .ip1(n10717), .ip2(n10740), .ip3(n11088), .op(n10756) );
  nand3_1 U12467 ( .ip1(n10720), .ip2(n10719), .ip3(n10718), .op(n10925) );
  nor3_1 U12468 ( .ip1(n10721), .ip2(n10925), .ip3(n10921), .op(n10755) );
  nor3_1 U12469 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip3(n10722), .op(n11014) );
  or2_1 U12470 ( .ip1(n10723), .ip2(n10740), .op(n10729) );
  nand2_1 U12471 ( .ip1(n10933), .ip2(n10724), .op(n10725) );
  nand2_1 U12472 ( .ip1(n10848), .ip2(n10725), .op(n10726) );
  nand2_1 U12473 ( .ip1(n10869), .ip2(n10726), .op(n10727) );
  or2_1 U12474 ( .ip1(n10727), .ip2(n10740), .op(n10728) );
  nand2_1 U12475 ( .ip1(n10729), .ip2(n10728), .op(n10730) );
  nor4_1 U12476 ( .ip1(n11014), .ip2(n10731), .ip3(n10730), .ip4(n10816), .op(
        n10753) );
  nor2_1 U12477 ( .ip1(n10949), .ip2(n11788), .op(n10733) );
  or2_1 U12478 ( .ip1(n10732), .ip2(n10733), .op(n10736) );
  or2_1 U12479 ( .ip1(n10734), .ip2(n10733), .op(n10735) );
  nand2_1 U12480 ( .ip1(n10736), .ip2(n10735), .op(n10738) );
  nor2_1 U12481 ( .ip1(n10738), .ip2(n10737), .op(n10749) );
  nor4_1 U12482 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n11786), .ip3(
        n10740), .ip4(n10739), .op(n10742) );
  or2_1 U12483 ( .ip1(n10741), .ip2(n10742), .op(n10745) );
  or2_1 U12484 ( .ip1(n10743), .ip2(n10742), .op(n10744) );
  nand2_1 U12485 ( .ip1(n10745), .ip2(n10744), .op(n10746) );
  nor2_1 U12486 ( .ip1(n10746), .ip2(n11682), .op(n10748) );
  nor2_1 U12487 ( .ip1(n12126), .ip2(n11789), .op(n10854) );
  nor2_1 U12488 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(n12070), .op(
        n10747) );
  nor4_1 U12489 ( .ip1(n10749), .ip2(n10748), .ip3(n10854), .ip4(n10747), .op(
        n10751) );
  nand4_1 U12490 ( .ip1(n12612), .ip2(n12320), .ip3(n10492), .ip4(n12122), 
        .op(n10750) );
  nand4_1 U12491 ( .ip1(n10753), .ip2(n10752), .ip3(n10751), .ip4(n10750), 
        .op(n10754) );
  nor4_1 U12492 ( .ip1(n10757), .ip2(n10756), .ip3(n10755), .ip4(n10754), .op(
        n10789) );
  or2_1 U12493 ( .ip1(n12624), .ip2(n10758), .op(n10760) );
  or2_1 U12494 ( .ip1(n11275), .ip2(n10758), .op(n10759) );
  nand2_1 U12495 ( .ip1(n10760), .ip2(n10759), .op(n10761) );
  nor2_1 U12496 ( .ip1(n10761), .ip2(n11693), .op(n10768) );
  inv_1 U12497 ( .ip(n10762), .op(n10763) );
  or2_1 U12498 ( .ip1(n10763), .ip2(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(
        n10766) );
  nand2_1 U12499 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n10764), .op(
        n10809) );
  or2_1 U12500 ( .ip1(n10809), .ip2(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(
        n10765) );
  nand2_1 U12501 ( .ip1(n10766), .ip2(n10765), .op(n10767) );
  not_ab_or_c_or_d U12502 ( .ip1(n10991), .ip2(n10769), .ip3(n10768), .ip4(
        n10767), .op(n10788) );
  nand2_1 U12503 ( .ip1(n11099), .ip2(n10770), .op(n10771) );
  nand2_1 U12504 ( .ip1(n10949), .ip2(n10771), .op(n10961) );
  nor2_1 U12505 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n10865), .op(
        n10775) );
  or2_1 U12506 ( .ip1(n11218), .ip2(n5639), .op(n10772) );
  nand2_1 U12507 ( .ip1(n10773), .ip2(n10772), .op(n10774) );
  not_ab_or_c_or_d U12508 ( .ip1(n10777), .ip2(n10776), .ip3(n10775), .ip4(
        n10774), .op(n10778) );
  nor2_1 U12509 ( .ip1(\CORTEXM0DS_INST/u_logic/Rkgvx4 ), .ip2(n10778), .op(
        n10781) );
  nor2_1 U12510 ( .ip1(n10779), .ip2(\CORTEXM0DS_INST/u_logic/P39vx4 ), .op(
        n10780) );
  nor2_1 U12511 ( .ip1(n10781), .ip2(n10780), .op(n10783) );
  nor2_1 U12512 ( .ip1(n10783), .ip2(n10782), .op(n10785) );
  and3_1 U12513 ( .ip1(n10955), .ip2(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip3(
        n10953), .op(n10784) );
  not_ab_or_c_or_d U12514 ( .ip1(n12116), .ip2(n10961), .ip3(n10785), .ip4(
        n10784), .op(n10787) );
  nand2_1 U12515 ( .ip1(n12641), .ip2(n10786), .op(n10995) );
  nand4_1 U12516 ( .ip1(n10789), .ip2(n10788), .ip3(n10787), .ip4(n10995), 
        .op(n10790) );
  not_ab_or_c_or_d U12517 ( .ip1(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip2(
        n10792), .ip3(n10791), .ip4(n10790), .op(n10793) );
  not_ab_or_c_or_d U12518 ( .ip1(n5932), .ip2(n12117), .ip3(1'b0), .ip4(n10793), .op(\CORTEXM0DS_INST/u_logic/Owhvx4 ) );
  nor4_1 U12519 ( .ip1(n12623), .ip2(n10795), .ip3(n10794), .ip4(
        \CORTEXM0DS_INST/u_logic/Ho8vx4 ), .op(n10800) );
  nand2_1 U12520 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(n10797) );
  not_ab_or_c_or_d U12521 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Ho8vx4 ), .ip3(n10797), .ip4(n10796), .op(
        n10799) );
  nor4_1 U12522 ( .ip1(n12389), .ip2(n10800), .ip3(n10799), .ip4(n10798), .op(
        n10899) );
  inv_1 U12523 ( .ip(n11184), .op(n10982) );
  nand2_1 U12524 ( .ip1(n10982), .ip2(n11228), .op(n10937) );
  inv_1 U12525 ( .ip(n10937), .op(n10802) );
  nor3_1 U12526 ( .ip1(n11755), .ip2(n11080), .ip3(n11680), .op(n10801) );
  not_ab_or_c_or_d U12527 ( .ip1(n11779), .ip2(n12138), .ip3(n10802), .ip4(
        n10801), .op(n10898) );
  not_ab_or_c_or_d U12528 ( .ip1(\CORTEXM0DS_INST/u_logic/P39vx4 ), .ip2(
        n10804), .ip3(n11146), .ip4(n10803), .op(n10808) );
  nand2_1 U12529 ( .ip1(n10805), .ip2(n11100), .op(n10807) );
  nand4_1 U12530 ( .ip1(n10808), .ip2(n10807), .ip3(n5092), .ip4(n10806), .op(
        n10817) );
  nor2_1 U12531 ( .ip1(n11693), .ip2(n10809), .op(n10812) );
  nor2_1 U12532 ( .ip1(n11796), .ip2(n10810), .op(n10811) );
  or4_1 U12533 ( .ip1(n10814), .ip2(n10813), .ip3(n10812), .ip4(n10811), .op(
        n10815) );
  not_ab_or_c_or_d U12534 ( .ip1(n10818), .ip2(n10817), .ip3(n10816), .ip4(
        n10815), .op(n10897) );
  nand2_1 U12535 ( .ip1(n10819), .ip2(n12583), .op(n10823) );
  nand2_1 U12536 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n10820), .op(
        n10822) );
  nand4_1 U12537 ( .ip1(n10824), .ip2(n10823), .ip3(n10822), .ip4(n10821), 
        .op(n10831) );
  or2_1 U12538 ( .ip1(n10825), .ip2(n12538), .op(n10829) );
  nand2_1 U12539 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n10826), .op(
        n10827) );
  or2_1 U12540 ( .ip1(n10827), .ip2(n12538), .op(n10828) );
  nand2_1 U12541 ( .ip1(n10829), .ip2(n10828), .op(n10830) );
  or2_1 U12542 ( .ip1(n10831), .ip2(n10830), .op(n10832) );
  nand2_1 U12543 ( .ip1(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip2(n10832), .op(
        n10834) );
  nor2_1 U12544 ( .ip1(n10834), .ip2(n10833), .op(n10882) );
  nor3_1 U12545 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n10835), .ip3(
        n12321), .op(n10846) );
  nor2_1 U12546 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(n12571), .op(
        n10858) );
  or2_1 U12547 ( .ip1(n10836), .ip2(n11190), .op(n10839) );
  or2_1 U12548 ( .ip1(n10837), .ip2(n11190), .op(n10838) );
  nand2_1 U12549 ( .ip1(n10839), .ip2(n10838), .op(n10840) );
  not_ab_or_c_or_d U12550 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(
        n10841), .ip3(n10858), .ip4(n10840), .op(n10843) );
  not_ab_or_c_or_d U12551 ( .ip1(n10844), .ip2(n10843), .ip3(
        \CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip4(n10842), .op(n10845) );
  not_ab_or_c_or_d U12552 ( .ip1(n12320), .ip2(n10932), .ip3(n10846), .ip4(
        n10845), .op(n10847) );
  or2_1 U12553 ( .ip1(n10847), .ip2(\CORTEXM0DS_INST/u_logic/Ho8vx4 ), .op(
        n10850) );
  or2_1 U12554 ( .ip1(n10848), .ip2(\CORTEXM0DS_INST/u_logic/Ho8vx4 ), .op(
        n10849) );
  nand2_1 U12555 ( .ip1(n10850), .ip2(n10849), .op(n10881) );
  nor2_1 U12556 ( .ip1(n10852), .ip2(n10851), .op(n10853) );
  or2_1 U12557 ( .ip1(n11131), .ip2(n10853), .op(n10856) );
  or2_1 U12558 ( .ip1(n10854), .ip2(n10853), .op(n10855) );
  nand2_1 U12559 ( .ip1(n10856), .ip2(n10855), .op(n10857) );
  nor2_1 U12560 ( .ip1(n10892), .ip2(n10857), .op(n10880) );
  nor2_1 U12561 ( .ip1(\CORTEXM0DS_INST/u_logic/Ki8vx4 ), .ip2(n12117), .op(
        n10943) );
  nor3_1 U12562 ( .ip1(n10859), .ip2(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip3(
        n10858), .op(n10860) );
  nor2_1 U12563 ( .ip1(n10860), .ip2(n11088), .op(n10861) );
  not_ab_or_c_or_d U12564 ( .ip1(n10943), .ip2(n10863), .ip3(n10862), .ip4(
        n10861), .op(n10878) );
  or2_1 U12565 ( .ip1(n10864), .ip2(n10865), .op(n10868) );
  nand3_1 U12566 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n11224), .ip3(
        n12117), .op(n10866) );
  or2_1 U12567 ( .ip1(n10866), .ip2(n10865), .op(n10867) );
  nand2_1 U12568 ( .ip1(n10868), .ip2(n10867), .op(n10871) );
  and2_1 U12569 ( .ip1(n10869), .ip2(n11107), .op(n10870) );
  not_ab_or_c_or_d U12570 ( .ip1(n10872), .ip2(n12124), .ip3(n10871), .ip4(
        n10870), .op(n10877) );
  nand3_1 U12571 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n11256), .ip3(
        n10873), .op(n10876) );
  nand2_1 U12572 ( .ip1(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip2(n10874), .op(
        n10875) );
  nand4_1 U12573 ( .ip1(n10878), .ip2(n10877), .ip3(n10876), .ip4(n10875), 
        .op(n10879) );
  or4_1 U12574 ( .ip1(n10882), .ip2(n10881), .ip3(n10880), .ip4(n10879), .op(
        n10895) );
  and3_1 U12575 ( .ip1(n11786), .ip2(n11703), .ip3(
        \CORTEXM0DS_INST/u_logic/Rkgvx4 ), .op(n10883) );
  not_ab_or_c_or_d U12576 ( .ip1(n10884), .ip2(n8424), .ip3(
        \CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip4(n10883), .op(n10886) );
  nor2_1 U12577 ( .ip1(n10886), .ip2(n10885), .op(n10894) );
  nor2_1 U12578 ( .ip1(n12126), .ip2(n10949), .op(n10887) );
  or2_1 U12579 ( .ip1(n11248), .ip2(n10887), .op(n10890) );
  or2_1 U12580 ( .ip1(n10888), .ip2(n10887), .op(n10889) );
  nand2_1 U12581 ( .ip1(n10890), .ip2(n10889), .op(n10891) );
  nor2_1 U12582 ( .ip1(n10892), .ip2(n10891), .op(n10893) );
  not_ab_or_c_or_d U12583 ( .ip1(n12125), .ip2(n10895), .ip3(n10894), .ip4(
        n10893), .op(n10896) );
  nand4_1 U12584 ( .ip1(n10899), .ip2(n10898), .ip3(n10897), .ip4(n10896), 
        .op(n10900) );
  mux2_1 U12585 ( .ip1(n10900), .ip2(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .s(
        n5932), .op(\CORTEXM0DS_INST/u_logic/Vwhvx4 ) );
  nor2_1 U12586 ( .ip1(n5814), .ip2(n10901), .op(n10902) );
  mux2_1 U12587 ( .ip1(n10902), .ip2(n5814), .s(\CORTEXM0DS_INST/vis_pc [0]), 
        .op(n10914) );
  nor2_1 U12588 ( .ip1(n11038), .ip2(n10903), .op(n10910) );
  nand2_1 U12589 ( .ip1(n11043), .ip2(n10904), .op(n10908) );
  nand2_1 U12590 ( .ip1(n10906), .ip2(n10905), .op(n10907) );
  nand3_1 U12591 ( .ip1(n10908), .ip2(n10907), .ip3(n11045), .op(n10909) );
  not_ab_or_c_or_d U12592 ( .ip1(n11037), .ip2(n10911), .ip3(n10910), .ip4(
        n10909), .op(n11534) );
  nor2_1 U12593 ( .ip1(n11534), .ip2(n10912), .op(n10913) );
  not_ab_or_c_or_d U12594 ( .ip1(n10916), .ip2(n10915), .ip3(n10914), .ip4(
        n10913), .op(n10918) );
  nand2_1 U12595 ( .ip1(n10918), .ip2(n10917), .op(
        \CORTEXM0DS_INST/u_logic/Cxhvx4 ) );
  or2_1 U12596 ( .ip1(n5639), .ip2(n10919), .op(n5013) );
  nor3_1 U12597 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n12623), .ip3(
        n5639), .op(n10920) );
  nor2_1 U12598 ( .ip1(n11802), .ip2(n10920), .op(n5014) );
  inv_1 U12599 ( .ip(n10921), .op(n10977) );
  nor2_1 U12600 ( .ip1(n11240), .ip2(n12072), .op(n10924) );
  and3_1 U12601 ( .ip1(n10922), .ip2(\CORTEXM0DS_INST/u_logic/Ih8vx4 ), .ip3(
        n11693), .op(n10923) );
  not_ab_or_c_or_d U12602 ( .ip1(n10977), .ip2(n10925), .ip3(n10924), .ip4(
        n10923), .op(n10969) );
  nor3_1 U12603 ( .ip1(\CORTEXM0DS_INST/u_logic/R89vx4 ), .ip2(n12562), .ip3(
        \CORTEXM0DS_INST/u_logic/K79vx4 ), .op(n10927) );
  nor2_1 U12604 ( .ip1(n10927), .ip2(n10926), .op(n10941) );
  inv_1 U12605 ( .ip(n10928), .op(n10929) );
  nor4_1 U12606 ( .ip1(n10932), .ip2(n10931), .ip3(n10930), .ip4(n10929), .op(
        n10940) );
  nand2_1 U12607 ( .ip1(n10991), .ip2(n10933), .op(n10935) );
  nand4_1 U12608 ( .ip1(n10937), .ip2(n10936), .ip3(n10935), .ip4(n10934), 
        .op(n10938) );
  nor4_1 U12609 ( .ip1(n10941), .ip2(n10940), .ip3(n10939), .ip4(n10938), .op(
        n10968) );
  nor3_1 U12610 ( .ip1(n10942), .ip2(n11084), .ip3(n11154), .op(n12084) );
  and3_1 U12611 ( .ip1(n12118), .ip2(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip3(
        n12084), .op(n12087) );
  nor2_1 U12612 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n10943), .op(
        n10947) );
  nor2_1 U12613 ( .ip1(n10945), .ip2(n10944), .op(n10946) );
  not_ab_or_c_or_d U12614 ( .ip1(n12087), .ip2(n11228), .ip3(n10947), .ip4(
        n10946), .op(n10948) );
  nand2_1 U12615 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n12623), .op(
        n11234) );
  not_ab_or_c_or_d U12616 ( .ip1(n10948), .ip2(n11234), .ip3(n10949), .ip4(
        n8424), .op(n10960) );
  not_ab_or_c_or_d U12617 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(
        n10950), .ip3(n11796), .ip4(n10949), .op(n10952) );
  not_ab_or_c_or_d U12618 ( .ip1(n10953), .ip2(n11228), .ip3(n10952), .ip4(
        n10951), .op(n10954) );
  or2_1 U12619 ( .ip1(n10954), .ip2(n10955), .op(n10958) );
  or2_1 U12620 ( .ip1(n10956), .ip2(n10955), .op(n10957) );
  nand2_1 U12621 ( .ip1(n10958), .ip2(n10957), .op(n10959) );
  not_ab_or_c_or_d U12622 ( .ip1(n10962), .ip2(n10961), .ip3(n10960), .ip4(
        n10959), .op(n10967) );
  nand4_1 U12623 ( .ip1(n10965), .ip2(n5639), .ip3(n10964), .ip4(n10963), .op(
        n10966) );
  nand4_1 U12624 ( .ip1(n10969), .ip2(n10968), .ip3(n10967), .ip4(n10966), 
        .op(n10970) );
  mux2_1 U12625 ( .ip1(n10970), .ip2(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .s(
        n5932), .op(\CORTEXM0DS_INST/u_logic/Xxhvx4 ) );
  nor2_1 U12626 ( .ip1(n11693), .ip2(n10971), .op(n11221) );
  and3_1 U12627 ( .ip1(n12121), .ip2(n11221), .ip3(n12117), .op(n10975) );
  nor4_1 U12628 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Q5gvx4 ), .ip3(n10973), .ip4(n10972), .op(
        n10974) );
  not_ab_or_c_or_d U12629 ( .ip1(n10977), .ip2(n10976), .ip3(n10975), .ip4(
        n10974), .op(n11002) );
  not_ab_or_c_or_d U12630 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(
        n10979), .ip3(n12599), .ip4(n10978), .op(n10980) );
  not_ab_or_c_or_d U12631 ( .ip1(n10982), .ip2(n8424), .ip3(n10981), .ip4(
        n10980), .op(n11001) );
  or2_1 U12632 ( .ip1(n10983), .ip2(n10984), .op(n10986) );
  or2_1 U12633 ( .ip1(n12118), .ip2(n10984), .op(n10985) );
  nand2_1 U12634 ( .ip1(n10986), .ip2(n10985), .op(n11185) );
  nand2_1 U12635 ( .ip1(n11185), .ip2(n10987), .op(n10999) );
  nor3_1 U12636 ( .ip1(n10989), .ip2(n10988), .ip3(n12627), .op(n10998) );
  nand3_1 U12637 ( .ip1(n10991), .ip2(n10492), .ip3(n10990), .op(n10994) );
  nand3_1 U12638 ( .ip1(n11267), .ip2(n11266), .ip3(n10992), .op(n10993) );
  nand4_1 U12639 ( .ip1(n10996), .ip2(n10995), .ip3(n10994), .ip4(n10993), 
        .op(n10997) );
  not_ab_or_c_or_d U12640 ( .ip1(n11786), .ip2(n10999), .ip3(n10998), .ip4(
        n10997), .op(n11000) );
  nand3_1 U12641 ( .ip1(n11002), .ip2(n11001), .ip3(n11000), .op(n11003) );
  mux2_1 U12642 ( .ip1(n11003), .ip2(\CORTEXM0DS_INST/u_logic/Dw8vx4 ), .s(
        n5932), .op(\CORTEXM0DS_INST/u_logic/Lyhvx4 ) );
  inv_1 U12643 ( .ip(n11004), .op(n11585) );
  not_ab_or_c_or_d U12644 ( .ip1(n11006), .ip2(n11005), .ip3(n12209), .ip4(
        n12343), .op(n11009) );
  nor2_1 U12645 ( .ip1(n11007), .ip2(n12311), .op(n11008) );
  not_ab_or_c_or_d U12646 ( .ip1(n12316), .ip2(n11585), .ip3(n11009), .ip4(
        n11008), .op(\CORTEXM0DS_INST/u_logic/N1447 ) );
  nand2_1 U12647 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [3]), .ip2(n4823), .op(
        n11019) );
  nor2_1 U12648 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n11764), .op(
        n11013) );
  nor4_1 U12649 ( .ip1(n11011), .ip2(n12623), .ip3(n12117), .ip4(n11010), .op(
        n11012) );
  or4_1 U12650 ( .ip1(n11014), .ip2(n11262), .ip3(n11013), .ip4(n11012), .op(
        n11687) );
  nand3_1 U12651 ( .ip1(n12648), .ip2(n11687), .ip3(n11051), .op(n11031) );
  inv_1 U12652 ( .ip(n11031), .op(n11073) );
  nand2_1 U12653 ( .ip1(n11073), .ip2(n11430), .op(n11018) );
  inv_1 U12654 ( .ip(n4823), .op(n12400) );
  nand2_1 U12655 ( .ip1(n11016), .ip2(n11015), .op(n12065) );
  nand2_1 U12656 ( .ip1(n12400), .ip2(n12065), .op(n12063) );
  nor2_1 U12657 ( .ip1(n12453), .ip2(n12063), .op(n11035) );
  nand2_1 U12658 ( .ip1(\CORTEXM0DS_INST/u_logic/Lrevx4 ), .ip2(n11035), .op(
        n11017) );
  nand3_1 U12659 ( .ip1(n11019), .ip2(n11018), .ip3(n11017), .op(
        \CORTEXM0DS_INST/u_logic/L8mvx4 ) );
  nand2_1 U12660 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [2]), .ip2(n4823), .op(
        n11022) );
  nand2_1 U12661 ( .ip1(n11073), .ip2(n11298), .op(n11021) );
  nand2_1 U12662 ( .ip1(\CORTEXM0DS_INST/u_logic/Bqevx4 ), .ip2(n11035), .op(
        n11020) );
  nand3_1 U12663 ( .ip1(n11022), .ip2(n11021), .ip3(n11020), .op(
        \CORTEXM0DS_INST/u_logic/U9mvx4 ) );
  nor2_1 U12664 ( .ip1(n11023), .ip2(n12400), .op(n11025) );
  nand2_1 U12665 ( .ip1(\CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Vsevx4 ), .op(n12456) );
  nor2_1 U12666 ( .ip1(n12456), .ip2(n12063), .op(n11024) );
  ab_or_c_or_d U12667 ( .ip1(n11073), .ip2(n11435), .ip3(n11025), .ip4(n11024), 
        .op(\CORTEXM0DS_INST/u_logic/Pamvx4 ) );
  nand2_1 U12668 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [5]), .ip2(n4823), .op(
        n11028) );
  nand2_1 U12669 ( .ip1(n11073), .ip2(n11442), .op(n11027) );
  nand2_1 U12670 ( .ip1(\CORTEXM0DS_INST/u_logic/Fuevx4 ), .ip2(n11035), .op(
        n11026) );
  nand3_1 U12671 ( .ip1(n11028), .ip2(n11027), .ip3(n11026), .op(
        \CORTEXM0DS_INST/u_logic/Wamvx4 ) );
  nand2_1 U12672 ( .ip1(\CORTEXM0DS_INST/u_logic/G8fvx4 ), .ip2(n11029), .op(
        n11030) );
  nand3_1 U12673 ( .ip1(n11030), .ip2(n4808), .ip3(n12062), .op(
        \CORTEXM0DS_INST/u_logic/G8nvx4 ) );
  nor2_1 U12674 ( .ip1(n11534), .ip2(n11031), .op(n11034) );
  nor2_1 U12675 ( .ip1(n11032), .ip2(n12400), .op(n11033) );
  ab_or_c_or_d U12676 ( .ip1(n11035), .ip2(\CORTEXM0DS_INST/u_logic/Roevx4 ), 
        .ip3(n11034), .ip4(n11033), .op(\CORTEXM0DS_INST/u_logic/Acnvx4 ) );
  nand2_1 U12677 ( .ip1(n11037), .ip2(n11036), .op(n11047) );
  nor2_1 U12678 ( .ip1(n4286), .ip2(n11038), .op(n11042) );
  nor2_1 U12679 ( .ip1(n11040), .ip2(n11039), .op(n11041) );
  not_ab_or_c_or_d U12680 ( .ip1(n11044), .ip2(n11043), .ip3(n11042), .ip4(
        n11041), .op(n11046) );
  nand3_1 U12681 ( .ip1(n11047), .ip2(n11046), .ip3(n11045), .op(n11526) );
  nor2_1 U12682 ( .ip1(n11048), .ip2(n12400), .op(n11050) );
  nand2_1 U12683 ( .ip1(\CORTEXM0DS_INST/u_logic/Hnevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Xlevx4 ), .op(n12459) );
  nor2_1 U12684 ( .ip1(n12459), .ip2(n12063), .op(n11049) );
  ab_or_c_or_d U12685 ( .ip1(n11073), .ip2(n11526), .ip3(n11050), .ip4(n11049), 
        .op(\CORTEXM0DS_INST/u_logic/Ocnvx4 ) );
  nor3_1 U12686 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip3(n11812), .op(n11668) );
  inv_1 U12687 ( .ip(n11668), .op(n11818) );
  nand2_1 U12688 ( .ip1(n11687), .ip2(n11051), .op(n11820) );
  nand2_1 U12689 ( .ip1(n11818), .ip2(n11820), .op(n11663) );
  inv_1 U12690 ( .ip(n11663), .op(n11825) );
  nor2_1 U12691 ( .ip1(n11511), .ip2(n11820), .op(n11054) );
  nor2_1 U12692 ( .ip1(n11052), .ip2(n11818), .op(n11053) );
  ab_or_c_or_d U12693 ( .ip1(n11825), .ip2(n11055), .ip3(n11054), .ip4(n11053), 
        .op(n11058) );
  not_ab_or_c_or_d U12694 ( .ip1(n11056), .ip2(n11825), .ip3(1'b0), .ip4(n5932), .op(n11057) );
  mux2_1 U12695 ( .ip1(\CORTEXM0DS_INST/vis_apsr [0]), .ip2(n11058), .s(n11057), .op(\CORTEXM0DS_INST/u_logic/Rhnvx4 ) );
  nor2_1 U12696 ( .ip1(n11060), .ip2(n11059), .op(n11062) );
  or2_1 U12697 ( .ip1(n11061), .ip2(n11062), .op(n11064) );
  or2_1 U12698 ( .ip1(n11526), .ip2(n11062), .op(n11063) );
  nand2_1 U12699 ( .ip1(n11064), .ip2(n11063), .op(n11072) );
  not_ab_or_c_or_d U12700 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(
        n11067), .ip3(n11066), .ip4(n11065), .op(n11068) );
  nor3_1 U12701 ( .ip1(n11068), .ip2(LOCKUP_top_out), .ip3(n12113), .op(n11069) );
  nor2_1 U12702 ( .ip1(n11073), .ip2(n11069), .op(n11070) );
  mux2_1 U12703 ( .ip1(n11072), .ip2(n11071), .s(n11070), .op(n11075) );
  nand2_1 U12704 ( .ip1(n11073), .ip2(n11456), .op(n11074) );
  nand2_1 U12705 ( .ip1(n11075), .ip2(n11074), .op(
        \CORTEXM0DS_INST/u_logic/Ojnvx4 ) );
  nor2_1 U12706 ( .ip1(n11856), .ip2(n12687), .op(n4705) );
  mux2_1 U12707 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [31]), .ip2(n12644), 
        .s(n4705), .op(\CORTEXM0DS_INST/u_logic/Vkmvx4 ) );
  inv_1 U12708 ( .ip(n3226), .op(n4704) );
  mux2_1 U12709 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [29]), .ip2(n4704), .s(
        n4705), .op(\CORTEXM0DS_INST/u_logic/Jlmvx4 ) );
  nand2_1 U12710 ( .ip1(n11863), .ip2(\CORTEXM0DS_INST/u_logic/Mf8vx4 ), .op(
        n4701) );
  mux2_1 U12711 ( .ip1(n12644), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [23]), 
        .s(n4701), .op(\CORTEXM0DS_INST/u_logic/Rimvx4 ) );
  mux2_1 U12712 ( .ip1(n4704), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [21]), .s(
        n4701), .op(\CORTEXM0DS_INST/u_logic/Fjmvx4 ) );
  and2_1 U12713 ( .ip1(n11864), .ip2(\CORTEXM0DS_INST/u_logic/Mf8vx4 ), .op(
        n4699) );
  mux2_1 U12714 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [15]), .ip2(n12644), 
        .s(n4699), .op(\CORTEXM0DS_INST/u_logic/Ngmvx4 ) );
  mux2_1 U12715 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [13]), .ip2(n4704), .s(
        n4699), .op(\CORTEXM0DS_INST/u_logic/Bhmvx4 ) );
  nand2_1 U12716 ( .ip1(n11841), .ip2(\CORTEXM0DS_INST/u_logic/Mf8vx4 ), .op(
        n4697) );
  mux2_1 U12717 ( .ip1(n12644), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [7]), .s(
        n4697), .op(\CORTEXM0DS_INST/u_logic/Jemvx4 ) );
  mux2_1 U12718 ( .ip1(n4704), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [5]), .s(
        n4697), .op(\CORTEXM0DS_INST/u_logic/Xemvx4 ) );
  or2_1 U12719 ( .ip1(n12624), .ip2(n11076), .op(n11078) );
  or2_1 U12720 ( .ip1(n11683), .ip2(n11076), .op(n11077) );
  nand2_1 U12721 ( .ip1(n11078), .ip2(n11077), .op(n11182) );
  nor2_1 U12722 ( .ip1(n11182), .ip2(n12453), .op(n11087) );
  nand2_1 U12723 ( .ip1(\CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip2(n11079), .op(
        n11083) );
  nor2_1 U12724 ( .ip1(n11080), .ip2(n11680), .op(n11082) );
  not_ab_or_c_or_d U12725 ( .ip1(n11099), .ip2(n12610), .ip3(n11082), .ip4(
        n11081), .op(n12086) );
  not_ab_or_c_or_d U12726 ( .ip1(n11084), .ip2(n11083), .ip3(n12086), .ip4(
        n12084), .op(n11086) );
  nor3_1 U12727 ( .ip1(n12132), .ip2(n12624), .ip3(n11782), .op(n11085) );
  not_ab_or_c_or_d U12728 ( .ip1(n11087), .ip2(
        \CORTEXM0DS_INST/u_logic/Lrevx4 ), .ip3(n11086), .ip4(n11085), .op(
        n11130) );
  not_ab_or_c_or_d U12729 ( .ip1(n11089), .ip2(n11088), .ip3(
        \CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip4(n10492), .op(n11164) );
  or2_1 U12730 ( .ip1(n11096), .ip2(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .op(
        n11092) );
  nand2_1 U12731 ( .ip1(n11101), .ip2(n11090), .op(n12089) );
  or2_1 U12732 ( .ip1(n12089), .ip2(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .op(
        n11091) );
  nand2_1 U12733 ( .ip1(n11092), .ip2(n11091), .op(n11148) );
  or2_1 U12734 ( .ip1(n11093), .ip2(n11148), .op(n11094) );
  nor2_1 U12735 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Aj9vx4 ), .op(n11145) );
  nand2_1 U12736 ( .ip1(n11094), .ip2(n11145), .op(n11095) );
  nor2_1 U12737 ( .ip1(n11095), .ip2(n12583), .op(n11098) );
  nor2_1 U12738 ( .ip1(n11100), .ip2(n11096), .op(n12093) );
  inv_1 U12739 ( .ip(n12093), .op(n12074) );
  nor2_1 U12740 ( .ip1(n11190), .ip2(n12074), .op(n11097) );
  not_ab_or_c_or_d U12741 ( .ip1(\CORTEXM0DS_INST/u_logic/I29vx4 ), .ip2(
        n11164), .ip3(n11098), .ip4(n11097), .op(n11129) );
  nand2_1 U12742 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n11099), .op(
        n11104) );
  nand4_1 U12743 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n11102), .ip3(
        n11101), .ip4(n11100), .op(n11103) );
  nand4_1 U12744 ( .ip1(n11106), .ip2(n11105), .ip3(n11104), .ip4(n11103), 
        .op(n11189) );
  nand2_1 U12745 ( .ip1(\CORTEXM0DS_INST/u_logic/P39vx4 ), .ip2(n11189), .op(
        n11128) );
  nand2_1 U12746 ( .ip1(n11108), .ip2(n11107), .op(n11109) );
  nand2_1 U12747 ( .ip1(n11110), .ip2(n11109), .op(n11193) );
  inv_1 U12748 ( .ip(n11111), .op(n11114) );
  mux2_1 U12749 ( .ip1(n11114), .ip2(n11111), .s(n11113), .op(n11118) );
  nand2_1 U12750 ( .ip1(\CORTEXM0DS_INST/u_logic/R89vx4 ), .ip2(n11118), .op(
        n11167) );
  fulladder U12751 ( .a(\CORTEXM0DS_INST/u_logic/B19vx4 ), .b(
        \CORTEXM0DS_INST/u_logic/I29vx4 ), .ci(
        \CORTEXM0DS_INST/u_logic/Uz8vx4 ), .co(n11121), .s(n11112) );
  fulladder U12752 ( .a(\CORTEXM0DS_INST/u_logic/W49vx4 ), .b(
        \CORTEXM0DS_INST/u_logic/P39vx4 ), .ci(n11112), .co(n11120), .s(n11113) );
  nand2_1 U12753 ( .ip1(\CORTEXM0DS_INST/u_logic/K79vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/D69vx4 ), .op(n11116) );
  nand2_1 U12754 ( .ip1(n11114), .ip2(n11113), .op(n11115) );
  nand2_1 U12755 ( .ip1(n11116), .ip2(n11115), .op(n11119) );
  inv_1 U12756 ( .ip(n11117), .op(n11166) );
  nor2_1 U12757 ( .ip1(n11167), .ip2(n11166), .op(n11122) );
  nand3_1 U12758 ( .ip1(n11122), .ip2(n11120), .ip3(n11121), .op(n11125) );
  mux2_1 U12759 ( .ip1(\CORTEXM0DS_INST/u_logic/R89vx4 ), .ip2(n12571), .s(
        n11118), .op(n11192) );
  nand3_1 U12760 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip3(n11192), .op(n11195) );
  nor2_1 U12761 ( .ip1(n11166), .ip2(n11195), .op(n11165) );
  nand2_1 U12762 ( .ip1(n11121), .ip2(n11120), .op(n11124) );
  fulladder U12763 ( .a(n11121), .b(n11120), .ci(n11119), .co(n11123), .s(
        n11117) );
  inv_1 U12764 ( .ip(n11122), .op(n11170) );
  mux2_1 U12765 ( .ip1(n11124), .ip2(n11123), .s(n11170), .op(n11142) );
  nand2_1 U12766 ( .ip1(n11165), .ip2(n11142), .op(n11144) );
  nand2_1 U12767 ( .ip1(n11125), .ip2(n11144), .op(n11126) );
  nand2_1 U12768 ( .ip1(n11193), .ip2(n11126), .op(n11127) );
  nand4_1 U12769 ( .ip1(n11130), .ip2(n11129), .ip3(n11128), .ip4(n11127), 
        .op(n11135) );
  inv_1 U12770 ( .ip(n11131), .op(n11133) );
  nand3_1 U12771 ( .ip1(n11133), .ip2(n12651), .ip3(n11132), .op(n11134) );
  nand2_1 U12772 ( .ip1(n4620), .ip2(n11134), .op(n11199) );
  mux2_1 U12773 ( .ip1(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .ip2(n11135), .s(
        n11199), .op(\CORTEXM0DS_INST/u_logic/N2mvx4 ) );
  or2_1 U12774 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n11136), .op(
        n11138) );
  or2_1 U12775 ( .ip1(n12552), .ip2(n11136), .op(n11137) );
  nand2_1 U12776 ( .ip1(n11138), .ip2(n11137), .op(n11179) );
  nor3_1 U12777 ( .ip1(\CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip2(n12086), .ip3(
        n11154), .op(n11139) );
  not_ab_or_c_or_d U12778 ( .ip1(n12093), .ip2(
        \CORTEXM0DS_INST/u_logic/R89vx4 ), .ip3(n11179), .ip4(n11139), .op(
        n11152) );
  inv_1 U12779 ( .ip(\CORTEXM0DS_INST/u_logic/Bqevx4 ), .op(n12553) );
  nor3_1 U12780 ( .ip1(n11182), .ip2(n12553), .ip3(n12453), .op(n11141) );
  and2_1 U12781 ( .ip1(n11189), .ip2(\CORTEXM0DS_INST/u_logic/I29vx4 ), .op(
        n11140) );
  not_ab_or_c_or_d U12782 ( .ip1(\CORTEXM0DS_INST/u_logic/B19vx4 ), .ip2(
        n11164), .ip3(n11141), .ip4(n11140), .op(n11151) );
  or2_1 U12783 ( .ip1(n11165), .ip2(n11142), .op(n11143) );
  nand3_1 U12784 ( .ip1(n11144), .ip2(n11143), .ip3(n11193), .op(n11150) );
  and2_1 U12785 ( .ip1(n11146), .ip2(n11145), .op(n11147) );
  nor2_1 U12786 ( .ip1(n11148), .ip2(n11147), .op(n11161) );
  inv_1 U12787 ( .ip(n11161), .op(n11183) );
  nand2_1 U12788 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n11183), .op(
        n11149) );
  nand4_1 U12789 ( .ip1(n11152), .ip2(n11151), .ip3(n11150), .ip4(n11149), 
        .op(n11153) );
  nand2_1 U12790 ( .ip1(n11153), .ip2(n11199), .op(n11157) );
  inv_1 U12791 ( .ip(n12086), .op(n11159) );
  nand2_1 U12792 ( .ip1(n11154), .ip2(n11159), .op(n11155) );
  nand2_1 U12793 ( .ip1(n11199), .ip2(n11155), .op(n11176) );
  nand2_1 U12794 ( .ip1(\CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip2(n11176), .op(
        n11156) );
  nand2_1 U12795 ( .ip1(n11157), .ip2(n11156), .op(
        \CORTEXM0DS_INST/u_logic/U2mvx4 ) );
  inv_1 U12796 ( .ip(\CORTEXM0DS_INST/u_logic/Roevx4 ), .op(n12547) );
  nor3_1 U12797 ( .ip1(n11182), .ip2(n12547), .ip3(n12453), .op(n11158) );
  not_ab_or_c_or_d U12798 ( .ip1(n11160), .ip2(n11159), .ip3(n11179), .ip4(
        n11158), .op(n11174) );
  nor2_1 U12799 ( .ip1(n11161), .ip2(n12571), .op(n11163) );
  nor2_1 U12800 ( .ip1(n12567), .ip2(n12074), .op(n11162) );
  not_ab_or_c_or_d U12801 ( .ip1(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), .ip2(
        n11164), .ip3(n11163), .ip4(n11162), .op(n11173) );
  inv_1 U12802 ( .ip(n11165), .op(n11169) );
  nand3_1 U12803 ( .ip1(n11167), .ip2(n11166), .ip3(n11195), .op(n11168) );
  nand4_1 U12804 ( .ip1(n11193), .ip2(n11170), .ip3(n11169), .ip4(n11168), 
        .op(n11172) );
  nand2_1 U12805 ( .ip1(\CORTEXM0DS_INST/u_logic/B19vx4 ), .ip2(n11189), .op(
        n11171) );
  nand4_1 U12806 ( .ip1(n11174), .ip2(n11173), .ip3(n11172), .ip4(n11171), 
        .op(n11175) );
  nand2_1 U12807 ( .ip1(n11199), .ip2(n11175), .op(n11178) );
  nand2_1 U12808 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n11176), .op(
        n11177) );
  nand2_1 U12809 ( .ip1(n11178), .ip2(n11177), .op(
        \CORTEXM0DS_INST/u_logic/Jdnvx4 ) );
  nor2_1 U12810 ( .ip1(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip2(n12086), .op(
        n11180) );
  not_ab_or_c_or_d U12811 ( .ip1(n11181), .ip2(n12592), .ip3(n11180), .ip4(
        n11179), .op(n11198) );
  nor2_1 U12812 ( .ip1(n11182), .ip2(n12459), .op(n11188) );
  nand2_1 U12813 ( .ip1(\CORTEXM0DS_INST/u_logic/K79vx4 ), .ip2(n11183), .op(
        n11186) );
  nand3_1 U12814 ( .ip1(n11186), .ip2(n11185), .ip3(n11184), .op(n11187) );
  not_ab_or_c_or_d U12815 ( .ip1(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), .ip2(
        n11189), .ip3(n11188), .ip4(n11187), .op(n11197) );
  nor2_1 U12816 ( .ip1(n11190), .ip2(n12599), .op(n11191) );
  or2_1 U12817 ( .ip1(n11192), .ip2(n11191), .op(n11194) );
  nand3_1 U12818 ( .ip1(n11195), .ip2(n11194), .ip3(n11193), .op(n11196) );
  nand4_1 U12819 ( .ip1(n11198), .ip2(n11197), .ip3(n11765), .ip4(n11196), 
        .op(n11200) );
  mux2_1 U12820 ( .ip1(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip2(n11200), .s(
        n11199), .op(\CORTEXM0DS_INST/u_logic/Tinvx4 ) );
  mux2_1 U12821 ( .ip1(n11201), .ip2(\CORTEXM0DS_INST/u_logic/Zph2z4 [1]), .s(
        n4578), .op(\CORTEXM0DS_INST/u_logic/X9kvx4 ) );
  mux2_1 U12822 ( .ip1(n12323), .ip2(\CORTEXM0DS_INST/u_logic/Zph2z4 [0]), .s(
        n4578), .op(\CORTEXM0DS_INST/u_logic/Ufnvx4 ) );
  not_ab_or_c_or_d U12823 ( .ip1(n11594), .ip2(n12662), .ip3(n11202), .ip4(
        n11761), .op(n11203) );
  nand2_1 U12824 ( .ip1(n11204), .ip2(n11203), .op(n11622) );
  nor2_1 U12825 ( .ip1(n11285), .ip2(n11205), .op(n11280) );
  nor2_1 U12826 ( .ip1(n11284), .ip2(n11206), .op(n11279) );
  nor2_1 U12827 ( .ip1(n11283), .ip2(n11207), .op(n11278) );
  or2_1 U12828 ( .ip1(n11208), .ip2(n11209), .op(n11211) );
  or2_1 U12829 ( .ip1(n5639), .ip2(n11209), .op(n11210) );
  nand2_1 U12830 ( .ip1(n11211), .ip2(n11210), .op(n11212) );
  or2_1 U12831 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n11212), .op(
        n11215) );
  nand4_1 U12832 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip3(n11782), .ip4(n11213), .op(
        n11214) );
  nand3_1 U12833 ( .ip1(n11216), .ip2(n11215), .ip3(n11214), .op(n11274) );
  not_ab_or_c_or_d U12834 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        n11218), .ip3(n11217), .ip4(n12610), .op(n11220) );
  nor3_1 U12835 ( .ip1(n11221), .ip2(n11220), .ip3(n11219), .op(n11222) );
  nor2_1 U12836 ( .ip1(n11222), .ip2(n12124), .op(n11273) );
  nor4_1 U12837 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n11228), .ip3(
        n12609), .ip4(n11763), .op(n11238) );
  nor2_1 U12838 ( .ip1(n11223), .ip2(n11680), .op(n11225) );
  or2_1 U12839 ( .ip1(n11224), .ip2(n11225), .op(n11227) );
  or2_1 U12840 ( .ip1(n12369), .ip2(n11225), .op(n11226) );
  nand2_1 U12841 ( .ip1(n11227), .ip2(n11226), .op(n11229) );
  nor2_1 U12842 ( .ip1(n11229), .ip2(n11228), .op(n11237) );
  inv_1 U12843 ( .ip(n11230), .op(n11233) );
  nor4_1 U12844 ( .ip1(n12125), .ip2(n11233), .ip3(n11232), .ip4(n11231), .op(
        n11236) );
  nor2_1 U12845 ( .ip1(n11765), .ip2(n11234), .op(n11235) );
  nor4_1 U12846 ( .ip1(n11238), .ip2(n11237), .ip3(n11236), .ip4(n11235), .op(
        n11271) );
  nor3_1 U12847 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(n11228), .ip3(
        n11239), .op(n11246) );
  nor4_1 U12848 ( .ip1(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip2(n11693), .ip3(
        n11241), .ip4(n11240), .op(n11245) );
  nor3_1 U12849 ( .ip1(n12117), .ip2(n11243), .ip3(n11242), .op(n11244) );
  nor4_1 U12850 ( .ip1(n11247), .ip2(n11246), .ip3(n11245), .ip4(n11244), .op(
        n11270) );
  nand3_1 U12851 ( .ip1(n11250), .ip2(n11249), .ip3(n11248), .op(n11255) );
  nand3_1 U12852 ( .ip1(n11253), .ip2(n11252), .ip3(n11251), .op(n11254) );
  nand2_1 U12853 ( .ip1(n11255), .ip2(n11254), .op(n11265) );
  nand3_1 U12854 ( .ip1(n11256), .ip2(n12656), .ip3(n8424), .op(n11261) );
  nand2_1 U12855 ( .ip1(n11257), .ip2(n12623), .op(n11260) );
  nand2_1 U12856 ( .ip1(n12133), .ip2(n11258), .op(n11259) );
  nand4_1 U12857 ( .ip1(n11796), .ip2(n11261), .ip3(n11260), .ip4(n11259), 
        .op(n11264) );
  not_ab_or_c_or_d U12858 ( .ip1(n11265), .ip2(n11264), .ip3(n11263), .ip4(
        n11262), .op(n11269) );
  nand3_1 U12859 ( .ip1(n11267), .ip2(n11266), .ip3(n12623), .op(n11268) );
  nand4_1 U12860 ( .ip1(n11271), .ip2(n11270), .ip3(n11269), .ip4(n11268), 
        .op(n11272) );
  not_ab_or_c_or_d U12861 ( .ip1(n11275), .ip2(n11274), .ip3(n11273), .ip4(
        n11272), .op(n11276) );
  nor2_1 U12862 ( .ip1(n5932), .ip2(n11276), .op(n11281) );
  nand2_1 U12863 ( .ip1(n11281), .ip2(n11277), .op(n11296) );
  nor4_1 U12864 ( .ip1(n11280), .ip2(n11279), .ip3(n11278), .ip4(n11296), .op(
        n11542) );
  nand2_1 U12865 ( .ip1(n11281), .ip2(n11601), .op(n11536) );
  nor2_1 U12866 ( .ip1(n11542), .ip2(n11536), .op(n11540) );
  inv_1 U12867 ( .ip(n11282), .op(n11295) );
  inv_1 U12868 ( .ip(n11283), .op(n11290) );
  nand2_1 U12869 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [2]), .ip2(n11290), 
        .op(n11288) );
  inv_1 U12870 ( .ip(n11284), .op(n11289) );
  nand2_1 U12871 ( .ip1(\CORTEXM0DS_INST/u_logic/Wv9vx4 ), .ip2(n11289), .op(
        n11287) );
  inv_1 U12872 ( .ip(n11285), .op(n11291) );
  nand2_1 U12873 ( .ip1(\CORTEXM0DS_INST/u_logic/Nt8vx4 ), .ip2(n11291), .op(
        n11286) );
  nand4_1 U12874 ( .ip1(n11295), .ip2(n11288), .ip3(n11287), .ip4(n11286), 
        .op(n11537) );
  nor2_1 U12875 ( .ip1(n11296), .ip2(n11537), .op(n11549) );
  nand2_1 U12876 ( .ip1(\CORTEXM0DS_INST/u_logic/Bx9vx4 ), .ip2(n11289), .op(
        n11294) );
  nand2_1 U12877 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [3]), .ip2(n11290), 
        .op(n11293) );
  nand2_1 U12878 ( .ip1(\CORTEXM0DS_INST/u_logic/Vu8vx4 ), .ip2(n11291), .op(
        n11292) );
  nand4_1 U12879 ( .ip1(n11295), .ip2(n11294), .ip3(n11293), .ip4(n11292), 
        .op(n11547) );
  nor2_1 U12880 ( .ip1(n11296), .ip2(n11547), .op(n11538) );
  nor2_1 U12881 ( .ip1(n11549), .ip2(n11538), .op(n11602) );
  nand2_1 U12882 ( .ip1(n11540), .ip2(n11602), .op(n11570) );
  nor2_1 U12883 ( .ip1(\CORTEXM0DS_INST/u_logic/O7evx4 ), .ip2(n11570), .op(
        n11506) );
  mux2_1 U12884 ( .ip1(\CORTEXM0DS_INST/vis_msp [7]), .ip2(n11622), .s(n11506), 
        .op(\CORTEXM0DS_INST/u_logic/Plivx4 ) );
  nor2_1 U12885 ( .ip1(n11297), .ip2(n11494), .op(n11300) );
  or4_1 U12886 ( .ip1(n11301), .ip2(n11300), .ip3(n11299), .ip4(n11298), .op(
        n11623) );
  buf_1 U12887 ( .ip(n11506), .op(n11599) );
  mux2_1 U12888 ( .ip1(\CORTEXM0DS_INST/vis_msp [0]), .ip2(n11623), .s(n11599), 
        .op(\CORTEXM0DS_INST/u_logic/Eqivx4 ) );
  not_ab_or_c_or_d U12889 ( .ip1(n11594), .ip2(n12663), .ip3(n11593), .ip4(
        n11302), .op(n11305) );
  nand3_1 U12890 ( .ip1(n11305), .ip2(n11304), .ip3(n11303), .op(n11624) );
  mux2_1 U12891 ( .ip1(\CORTEXM0DS_INST/vis_msp [8]), .ip2(n11624), .s(n11506), 
        .op(\CORTEXM0DS_INST/u_logic/Tuivx4 ) );
  nor2_1 U12892 ( .ip1(n12665), .ip2(n11494), .op(n11306) );
  not_ab_or_c_or_d U12893 ( .ip1(n11308), .ip2(n11558), .ip3(n11307), .ip4(
        n11306), .op(n11314) );
  nor2_1 U12894 ( .ip1(n11501), .ip2(n11309), .op(n11311) );
  not_ab_or_c_or_d U12895 ( .ip1(n11312), .ip2(n11578), .ip3(n11311), .ip4(
        n11310), .op(n11313) );
  nand3_1 U12896 ( .ip1(n11314), .ip2(n11313), .ip3(n11438), .op(n11625) );
  mux2_1 U12897 ( .ip1(\CORTEXM0DS_INST/vis_msp [9]), .ip2(n11625), .s(n11599), 
        .op(\CORTEXM0DS_INST/u_logic/Izivx4 ) );
  inv_1 U12898 ( .ip(n11315), .op(n12666) );
  or2_1 U12899 ( .ip1(n11581), .ip2(n11316), .op(n11317) );
  nand2_1 U12900 ( .ip1(n11322), .ip2(n11317), .op(n11319) );
  or2_1 U12901 ( .ip1(n11583), .ip2(n11319), .op(n11321) );
  inv_1 U12902 ( .ip(n11318), .op(n12201) );
  or2_1 U12903 ( .ip1(n12201), .ip2(n11319), .op(n11320) );
  nand2_1 U12904 ( .ip1(n11321), .ip2(n11320), .op(n11324) );
  nor2_1 U12905 ( .ip1(n11322), .ip2(n11588), .op(n11323) );
  nor2_1 U12906 ( .ip1(n11324), .ip2(n11323), .op(n11325) );
  not_ab_or_c_or_d U12907 ( .ip1(n11594), .ip2(n12666), .ip3(n11593), .ip4(
        n11325), .op(n11328) );
  nand2_1 U12908 ( .ip1(n11326), .ip2(n11578), .op(n11327) );
  nand3_1 U12909 ( .ip1(n11329), .ip2(n11328), .ip3(n11327), .op(n11626) );
  mux2_1 U12910 ( .ip1(\CORTEXM0DS_INST/vis_msp [10]), .ip2(n11626), .s(n11506), .op(\CORTEXM0DS_INST/u_logic/X3jvx4 ) );
  inv_1 U12911 ( .ip(n11330), .op(n12667) );
  nor2_1 U12912 ( .ip1(n11581), .ip2(n11331), .op(n11332) );
  not_ab_or_c_or_d U12913 ( .ip1(n11594), .ip2(n12667), .ip3(n11333), .ip4(
        n11332), .op(n11339) );
  nor2_1 U12914 ( .ip1(n11501), .ip2(n11334), .op(n11336) );
  not_ab_or_c_or_d U12915 ( .ip1(n11337), .ip2(n11578), .ip3(n11336), .ip4(
        n11335), .op(n11338) );
  nand3_1 U12916 ( .ip1(n11339), .ip2(n11338), .ip3(n11438), .op(n11627) );
  mux2_1 U12917 ( .ip1(\CORTEXM0DS_INST/vis_msp [11]), .ip2(n11627), .s(n11599), .op(\CORTEXM0DS_INST/u_logic/M8jvx4 ) );
  nor2_1 U12918 ( .ip1(n11340), .ip2(n11494), .op(n11341) );
  not_ab_or_c_or_d U12919 ( .ip1(n11343), .ip2(n11558), .ip3(n11342), .ip4(
        n11341), .op(n11349) );
  nor2_1 U12920 ( .ip1(n11501), .ip2(n11344), .op(n11346) );
  not_ab_or_c_or_d U12921 ( .ip1(n11347), .ip2(n11578), .ip3(n11346), .ip4(
        n11345), .op(n11348) );
  nand3_1 U12922 ( .ip1(n11349), .ip2(n11348), .ip3(n11438), .op(n11628) );
  mux2_1 U12923 ( .ip1(\CORTEXM0DS_INST/vis_msp [12]), .ip2(n11628), .s(n11506), .op(\CORTEXM0DS_INST/u_logic/Bdjvx4 ) );
  inv_1 U12924 ( .ip(n11350), .op(n11354) );
  nor2_1 U12925 ( .ip1(n11501), .ip2(n11351), .op(n11352) );
  not_ab_or_c_or_d U12926 ( .ip1(n11558), .ip2(n11354), .ip3(n11353), .ip4(
        n11352), .op(n11360) );
  nor2_1 U12927 ( .ip1(n11593), .ip2(n11355), .op(n11577) );
  inv_1 U12928 ( .ip(n11577), .op(n11420) );
  not_ab_or_c_or_d U12929 ( .ip1(n11357), .ip2(n11578), .ip3(n11420), .ip4(
        n11356), .op(n11359) );
  nand3_1 U12930 ( .ip1(n11360), .ip2(n11359), .ip3(n11358), .op(n11629) );
  mux2_1 U12931 ( .ip1(\CORTEXM0DS_INST/vis_msp [14]), .ip2(n11629), .s(n11599), .op(\CORTEXM0DS_INST/u_logic/Qhjvx4 ) );
  nor2_1 U12932 ( .ip1(n12672), .ip2(n11494), .op(n11369) );
  nor2_1 U12933 ( .ip1(n11588), .ip2(n11361), .op(n11366) );
  or2_1 U12934 ( .ip1(n11558), .ip2(n12225), .op(n11364) );
  or2_1 U12935 ( .ip1(n11362), .ip2(n12225), .op(n11363) );
  nand2_1 U12936 ( .ip1(n11364), .ip2(n11363), .op(n11365) );
  not_ab_or_c_or_d U12937 ( .ip1(n11367), .ip2(n11564), .ip3(n11366), .ip4(
        n11365), .op(n11368) );
  not_ab_or_c_or_d U12938 ( .ip1(n11370), .ip2(n11578), .ip3(n11369), .ip4(
        n11368), .op(n11371) );
  nand3_1 U12939 ( .ip1(n11577), .ip2(n11372), .ip3(n11371), .op(n11630) );
  mux2_1 U12940 ( .ip1(\CORTEXM0DS_INST/vis_msp [15]), .ip2(n11630), .s(n11506), .op(\CORTEXM0DS_INST/u_logic/Fmjvx4 ) );
  nor2_1 U12941 ( .ip1(n11501), .ip2(n11373), .op(n11375) );
  nor2_1 U12942 ( .ip1(n12670), .ip2(n11494), .op(n11374) );
  not_ab_or_c_or_d U12943 ( .ip1(n11376), .ip2(n11558), .ip3(n11375), .ip4(
        n11374), .op(n11381) );
  inv_1 U12944 ( .ip(n12232), .op(n11378) );
  not_ab_or_c_or_d U12945 ( .ip1(n11378), .ip2(n11578), .ip3(n11420), .ip4(
        n11377), .op(n11380) );
  nand3_1 U12946 ( .ip1(n11381), .ip2(n11380), .ip3(n11379), .op(n11631) );
  mux2_1 U12947 ( .ip1(\CORTEXM0DS_INST/vis_msp [16]), .ip2(n11631), .s(n11599), .op(\CORTEXM0DS_INST/u_logic/Uqjvx4 ) );
  inv_1 U12948 ( .ip(n11382), .op(n12676) );
  nor2_1 U12949 ( .ip1(n11588), .ip2(n11383), .op(n11389) );
  or2_1 U12950 ( .ip1(n11558), .ip2(n11384), .op(n11387) );
  or2_1 U12951 ( .ip1(n11385), .ip2(n11384), .op(n11386) );
  nand2_1 U12952 ( .ip1(n11387), .ip2(n11386), .op(n11388) );
  not_ab_or_c_or_d U12953 ( .ip1(n11390), .ip2(n11564), .ip3(n11389), .ip4(
        n11388), .op(n11392) );
  not_ab_or_c_or_d U12954 ( .ip1(n11594), .ip2(n12676), .ip3(n11392), .ip4(
        n11391), .op(n11394) );
  nand3_1 U12955 ( .ip1(n11577), .ip2(n11394), .ip3(n11393), .op(n11632) );
  mux2_1 U12956 ( .ip1(\CORTEXM0DS_INST/vis_msp [17]), .ip2(n11632), .s(n11506), .op(\CORTEXM0DS_INST/u_logic/Jvjvx4 ) );
  nor2_1 U12957 ( .ip1(n11501), .ip2(n11395), .op(n11399) );
  nor2_1 U12958 ( .ip1(n12674), .ip2(n11494), .op(n11398) );
  nor2_1 U12959 ( .ip1(n11581), .ip2(n11396), .op(n11397) );
  nor4_1 U12960 ( .ip1(n11400), .ip2(n11399), .ip3(n11398), .ip4(n11397), .op(
        n11403) );
  nand2_1 U12961 ( .ip1(n11401), .ip2(n11578), .op(n11402) );
  nand4_1 U12962 ( .ip1(n11404), .ip2(n11577), .ip3(n11403), .ip4(n11402), 
        .op(n11633) );
  mux2_1 U12963 ( .ip1(\CORTEXM0DS_INST/vis_msp [18]), .ip2(n11633), .s(n11599), .op(\CORTEXM0DS_INST/u_logic/Yzjvx4 ) );
  or2_1 U12964 ( .ip1(n11405), .ip2(n11406), .op(n11409) );
  nand2_1 U12965 ( .ip1(n11501), .ip2(n12266), .op(n11407) );
  or2_1 U12966 ( .ip1(n11407), .ip2(n11406), .op(n11408) );
  nand2_1 U12967 ( .ip1(n11409), .ip2(n11408), .op(n11411) );
  or2_1 U12968 ( .ip1(n11410), .ip2(n11411), .op(n11413) );
  or2_1 U12969 ( .ip1(n11581), .ip2(n11411), .op(n11412) );
  nand2_1 U12970 ( .ip1(n11413), .ip2(n11412), .op(n11414) );
  not_ab_or_c_or_d U12971 ( .ip1(n11594), .ip2(n12678), .ip3(n11415), .ip4(
        n11414), .op(n11416) );
  nand3_1 U12972 ( .ip1(n11577), .ip2(n11417), .ip3(n11416), .op(n11634) );
  mux2_1 U12973 ( .ip1(\CORTEXM0DS_INST/vis_msp [19]), .ip2(n11634), .s(n11506), .op(\CORTEXM0DS_INST/u_logic/N4kvx4 ) );
  nand2_1 U12974 ( .ip1(n11418), .ip2(n11558), .op(n11426) );
  not_ab_or_c_or_d U12975 ( .ip1(n12276), .ip2(n11578), .ip3(n11420), .ip4(
        n11419), .op(n11425) );
  nor2_1 U12976 ( .ip1(n11501), .ip2(n11421), .op(n11422) );
  not_ab_or_c_or_d U12977 ( .ip1(n11594), .ip2(n12680), .ip3(n11423), .ip4(
        n11422), .op(n11424) );
  nand3_1 U12978 ( .ip1(n11426), .ip2(n11425), .ip3(n11424), .op(n11635) );
  mux2_1 U12979 ( .ip1(\CORTEXM0DS_INST/vis_msp [20]), .ip2(n11635), .s(n11506), .op(\CORTEXM0DS_INST/u_logic/C9kvx4 ) );
  nor2_1 U12980 ( .ip1(n11438), .ip2(n11811), .op(n11429) );
  and2_1 U12981 ( .ip1(n11427), .ip2(\CORTEXM0DS_INST/vis_ipsr [3]), .op(
        n11428) );
  not_ab_or_c_or_d U12982 ( .ip1(n11594), .ip2(n12677), .ip3(n11429), .ip4(
        n11428), .op(n11434) );
  not_ab_or_c_or_d U12983 ( .ip1(n11432), .ip2(n11578), .ip3(n11431), .ip4(
        n11430), .op(n11433) );
  nand2_1 U12984 ( .ip1(n11434), .ip2(n11433), .op(n11636) );
  mux2_1 U12985 ( .ip1(\CORTEXM0DS_INST/vis_msp [1]), .ip2(n11636), .s(n11506), 
        .op(\CORTEXM0DS_INST/u_logic/Ydkvx4 ) );
  not_ab_or_c_or_d U12986 ( .ip1(n11437), .ip2(n11578), .ip3(n11436), .ip4(
        n11435), .op(n11439) );
  nand3_1 U12987 ( .ip1(n11440), .ip2(n11439), .ip3(n11438), .op(n11637) );
  mux2_1 U12988 ( .ip1(\CORTEXM0DS_INST/vis_msp [2]), .ip2(n11637), .s(n11506), 
        .op(\CORTEXM0DS_INST/u_logic/Nikvx4 ) );
  inv_1 U12989 ( .ip(n11441), .op(n11443) );
  or4_1 U12990 ( .ip1(n11445), .ip2(n11444), .ip3(n11443), .ip4(n11442), .op(
        n11638) );
  mux2_1 U12991 ( .ip1(\CORTEXM0DS_INST/vis_msp [3]), .ip2(n11638), .s(n11506), 
        .op(\CORTEXM0DS_INST/u_logic/Cnkvx4 ) );
  nor2_1 U12992 ( .ip1(n11581), .ip2(n11446), .op(n11447) );
  not_ab_or_c_or_d U12993 ( .ip1(n11594), .ip2(n12681), .ip3(n11593), .ip4(
        n11447), .op(n11454) );
  nor2_1 U12994 ( .ip1(n11501), .ip2(n11448), .op(n11450) );
  not_ab_or_c_or_d U12995 ( .ip1(n11451), .ip2(n11578), .ip3(n11450), .ip4(
        n11449), .op(n11453) );
  nand3_1 U12996 ( .ip1(n11454), .ip2(n11453), .ip3(n11452), .op(n11639) );
  mux2_1 U12997 ( .ip1(\CORTEXM0DS_INST/vis_msp [4]), .ip2(n11639), .s(n11599), 
        .op(\CORTEXM0DS_INST/u_logic/Rrkvx4 ) );
  nand2_1 U12998 ( .ip1(n12351), .ip2(n11578), .op(n11460) );
  inv_1 U12999 ( .ip(n11455), .op(n11457) );
  not_ab_or_c_or_d U13000 ( .ip1(n11594), .ip2(n11457), .ip3(n11593), .ip4(
        n11456), .op(n11459) );
  nand3_1 U13001 ( .ip1(n11460), .ip2(n11459), .ip3(n11458), .op(n11640) );
  mux2_1 U13002 ( .ip1(\CORTEXM0DS_INST/vis_msp [22]), .ip2(n11640), .s(n11506), .op(\CORTEXM0DS_INST/u_logic/Gwkvx4 ) );
  nor2_1 U13003 ( .ip1(n11581), .ip2(n11461), .op(n11464) );
  nor2_1 U13004 ( .ip1(n11462), .ip2(n11494), .op(n11463) );
  nor4_1 U13005 ( .ip1(n11593), .ip2(n11465), .ip3(n11464), .ip4(n11463), .op(
        n11468) );
  inv_1 U13006 ( .ip(n11466), .op(n11467) );
  nand3_1 U13007 ( .ip1(n11469), .ip2(n11468), .ip3(n11467), .op(n11641) );
  mux2_1 U13008 ( .ip1(\CORTEXM0DS_INST/vis_msp [23]), .ip2(n11641), .s(n11599), .op(\CORTEXM0DS_INST/u_logic/O0lvx4 ) );
  nor2_1 U13009 ( .ip1(n11470), .ip2(n11588), .op(n11475) );
  or2_1 U13010 ( .ip1(n11558), .ip2(n12304), .op(n11473) );
  or2_1 U13011 ( .ip1(n11471), .ip2(n12304), .op(n11472) );
  nand2_1 U13012 ( .ip1(n11473), .ip2(n11472), .op(n11474) );
  not_ab_or_c_or_d U13013 ( .ip1(n11564), .ip2(n11476), .ip3(n11475), .ip4(
        n11474), .op(n11479) );
  nor2_1 U13014 ( .ip1(n11477), .ip2(n11494), .op(n11478) );
  nor4_1 U13015 ( .ip1(n11593), .ip2(n11480), .ip3(n11479), .ip4(n11478), .op(
        n11481) );
  nand2_1 U13016 ( .ip1(n11482), .ip2(n11481), .op(n11642) );
  mux2_1 U13017 ( .ip1(\CORTEXM0DS_INST/vis_msp [24]), .ip2(n11642), .s(n11506), .op(\CORTEXM0DS_INST/u_logic/D5lvx4 ) );
  not_ab_or_c_or_d U13018 ( .ip1(n11594), .ip2(n11484), .ip3(n11593), .ip4(
        n11483), .op(n11486) );
  nand3_1 U13019 ( .ip1(n11487), .ip2(n11486), .ip3(n11485), .op(n11644) );
  mux2_1 U13020 ( .ip1(\CORTEXM0DS_INST/vis_msp [25]), .ip2(n11644), .s(n11599), .op(\CORTEXM0DS_INST/u_logic/S9lvx4 ) );
  or2_1 U13021 ( .ip1(n11594), .ip2(n11593), .op(n11490) );
  or2_1 U13022 ( .ip1(n11488), .ip2(n11593), .op(n11489) );
  nand2_1 U13023 ( .ip1(n11490), .ip2(n11489), .op(n11492) );
  nand4_1 U13024 ( .ip1(n11493), .ip2(n11821), .ip3(n11492), .ip4(n11491), 
        .op(n11647) );
  mux2_1 U13025 ( .ip1(\CORTEXM0DS_INST/vis_msp [27]), .ip2(n11647), .s(n11506), .op(\CORTEXM0DS_INST/u_logic/Helvx4 ) );
  nor2_1 U13026 ( .ip1(n11671), .ip2(n11494), .op(n11495) );
  ab_or_c_or_d U13027 ( .ip1(n11496), .ip2(\CORTEXM0DS_INST/vis_apsr [2]), 
        .ip3(n11593), .ip4(n11495), .op(n11497) );
  not_ab_or_c_or_d U13028 ( .ip1(n11499), .ip2(n11558), .ip3(n11498), .ip4(
        n11497), .op(n11504) );
  or2_1 U13029 ( .ip1(n11501), .ip2(n11500), .op(n11502) );
  nand4_1 U13030 ( .ip1(n11672), .ip2(n11504), .ip3(n11503), .ip4(n11502), 
        .op(n11648) );
  mux2_1 U13031 ( .ip1(\CORTEXM0DS_INST/vis_msp [28]), .ip2(n11648), .s(n11599), .op(\CORTEXM0DS_INST/u_logic/Djlvx4 ) );
  nand2_1 U13032 ( .ip1(n11505), .ip2(n11662), .op(n11654) );
  mux2_1 U13033 ( .ip1(\CORTEXM0DS_INST/vis_msp [29]), .ip2(n11654), .s(n11506), .op(\CORTEXM0DS_INST/u_logic/Rjlvx4 ) );
  inv_1 U13034 ( .ip(n11507), .op(n11510) );
  nand2_1 U13035 ( .ip1(n11594), .ip2(n11508), .op(n11509) );
  nand4_1 U13036 ( .ip1(n11512), .ip2(n11511), .ip3(n11510), .ip4(n11509), 
        .op(n11652) );
  mux2_1 U13037 ( .ip1(\CORTEXM0DS_INST/vis_msp [26]), .ip2(n11652), .s(n11599), .op(\CORTEXM0DS_INST/u_logic/Yjlvx4 ) );
  or2_1 U13038 ( .ip1(n11514), .ip2(n11513), .op(n11651) );
  mux2_1 U13039 ( .ip1(\CORTEXM0DS_INST/vis_msp [5]), .ip2(n11651), .s(n11599), 
        .op(\CORTEXM0DS_INST/u_logic/Fklvx4 ) );
  nand3_1 U13040 ( .ip1(n11542), .ip2(n11601), .ip3(n11602), .op(n11531) );
  mux2_1 U13041 ( .ip1(n11622), .ip2(\CORTEXM0DS_INST/cm0_r12 [9]), .s(n11531), 
        .op(\CORTEXM0DS_INST/u_logic/Blivx4 ) );
  buf_1 U13042 ( .ip(n11531), .op(n11605) );
  mux2_1 U13043 ( .ip1(n11623), .ip2(\CORTEXM0DS_INST/cm0_r12 [2]), .s(n11605), 
        .op(\CORTEXM0DS_INST/u_logic/Qpivx4 ) );
  mux2_1 U13044 ( .ip1(n11624), .ip2(\CORTEXM0DS_INST/cm0_r12 [10]), .s(n11531), .op(\CORTEXM0DS_INST/u_logic/Fuivx4 ) );
  mux2_1 U13045 ( .ip1(n11625), .ip2(\CORTEXM0DS_INST/cm0_r12 [11]), .s(n11605), .op(\CORTEXM0DS_INST/u_logic/Uyivx4 ) );
  mux2_1 U13046 ( .ip1(n11626), .ip2(\CORTEXM0DS_INST/cm0_r12 [12]), .s(n11531), .op(\CORTEXM0DS_INST/u_logic/J3jvx4 ) );
  mux2_1 U13047 ( .ip1(n11627), .ip2(\CORTEXM0DS_INST/cm0_r12 [13]), .s(n11605), .op(\CORTEXM0DS_INST/u_logic/Y7jvx4 ) );
  mux2_1 U13048 ( .ip1(n11628), .ip2(\CORTEXM0DS_INST/cm0_r12 [14]), .s(n11531), .op(\CORTEXM0DS_INST/u_logic/Ncjvx4 ) );
  mux2_1 U13049 ( .ip1(n11629), .ip2(\CORTEXM0DS_INST/cm0_r12 [16]), .s(n11605), .op(\CORTEXM0DS_INST/u_logic/Chjvx4 ) );
  mux2_1 U13050 ( .ip1(n11630), .ip2(\CORTEXM0DS_INST/cm0_r12 [17]), .s(n11531), .op(\CORTEXM0DS_INST/u_logic/Rljvx4 ) );
  mux2_1 U13051 ( .ip1(n11631), .ip2(\CORTEXM0DS_INST/cm0_r12 [18]), .s(n11605), .op(\CORTEXM0DS_INST/u_logic/Gqjvx4 ) );
  mux2_1 U13052 ( .ip1(n11632), .ip2(\CORTEXM0DS_INST/cm0_r12 [19]), .s(n11531), .op(\CORTEXM0DS_INST/u_logic/Vujvx4 ) );
  mux2_1 U13053 ( .ip1(n11633), .ip2(\CORTEXM0DS_INST/cm0_r12 [20]), .s(n11605), .op(\CORTEXM0DS_INST/u_logic/Kzjvx4 ) );
  mux2_1 U13054 ( .ip1(n11634), .ip2(\CORTEXM0DS_INST/cm0_r12 [21]), .s(n11531), .op(\CORTEXM0DS_INST/u_logic/Z3kvx4 ) );
  mux2_1 U13055 ( .ip1(n11635), .ip2(\CORTEXM0DS_INST/cm0_r12 [22]), .s(n11531), .op(\CORTEXM0DS_INST/u_logic/O8kvx4 ) );
  mux2_1 U13056 ( .ip1(n11636), .ip2(\CORTEXM0DS_INST/cm0_r12 [3]), .s(n11531), 
        .op(\CORTEXM0DS_INST/u_logic/Kdkvx4 ) );
  mux2_1 U13057 ( .ip1(n11637), .ip2(\CORTEXM0DS_INST/cm0_r12 [4]), .s(n11531), 
        .op(\CORTEXM0DS_INST/u_logic/Zhkvx4 ) );
  mux2_1 U13058 ( .ip1(n11638), .ip2(\CORTEXM0DS_INST/cm0_r12 [5]), .s(n11531), 
        .op(\CORTEXM0DS_INST/u_logic/Omkvx4 ) );
  mux2_1 U13059 ( .ip1(n11639), .ip2(\CORTEXM0DS_INST/cm0_r12 [6]), .s(n11531), 
        .op(\CORTEXM0DS_INST/u_logic/Drkvx4 ) );
  mux2_1 U13060 ( .ip1(n11640), .ip2(\CORTEXM0DS_INST/cm0_r12 [24]), .s(n11531), .op(\CORTEXM0DS_INST/u_logic/Svkvx4 ) );
  mux2_1 U13061 ( .ip1(n11641), .ip2(\CORTEXM0DS_INST/cm0_r12 [25]), .s(n11605), .op(\CORTEXM0DS_INST/u_logic/A0lvx4 ) );
  mux2_1 U13062 ( .ip1(n11642), .ip2(\CORTEXM0DS_INST/cm0_r12 [26]), .s(n11531), .op(\CORTEXM0DS_INST/u_logic/P4lvx4 ) );
  mux2_1 U13063 ( .ip1(n11644), .ip2(\CORTEXM0DS_INST/cm0_r12 [27]), .s(n11605), .op(\CORTEXM0DS_INST/u_logic/E9lvx4 ) );
  mux2_1 U13064 ( .ip1(n11647), .ip2(\CORTEXM0DS_INST/cm0_r12 [29]), .s(n11531), .op(\CORTEXM0DS_INST/u_logic/Tdlvx4 ) );
  mux2_1 U13065 ( .ip1(n11648), .ip2(\CORTEXM0DS_INST/cm0_r12 [30]), .s(n11605), .op(\CORTEXM0DS_INST/u_logic/Pilvx4 ) );
  nor2_1 U13066 ( .ip1(n11516), .ip2(n11515), .op(n11518) );
  or2_1 U13067 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [0]), .ip2(n11518), .op(n11521) );
  nor2_1 U13068 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(n11517), .op(
        n11519) );
  or2_1 U13069 ( .ip1(n11519), .ip2(n11518), .op(n11520) );
  nand2_1 U13070 ( .ip1(n11521), .ip2(n11520), .op(n11523) );
  nor2_1 U13071 ( .ip1(n11523), .ip2(n11522), .op(n11524) );
  not_ab_or_c_or_d U13072 ( .ip1(n11594), .ip2(n11525), .ip3(n11524), .ip4(
        n11593), .op(n11530) );
  not_ab_or_c_or_d U13073 ( .ip1(n11528), .ip2(n11578), .ip3(n11527), .ip4(
        n11526), .op(n11529) );
  nand2_1 U13074 ( .ip1(n11530), .ip2(n11529), .op(n11649) );
  mux2_1 U13075 ( .ip1(n11649), .ip2(\CORTEXM0DS_INST/cm0_r12 [0]), .s(n11531), 
        .op(\CORTEXM0DS_INST/u_logic/Mrlvx4 ) );
  nand2_1 U13076 ( .ip1(n11594), .ip2(n12673), .op(n11532) );
  nand4_1 U13077 ( .ip1(n11535), .ip2(n11534), .ip3(n11533), .ip4(n11532), 
        .op(n11650) );
  mux2_1 U13078 ( .ip1(n11650), .ip2(\CORTEXM0DS_INST/cm0_r12 [1]), .s(n11605), 
        .op(\CORTEXM0DS_INST/u_logic/Trlvx4 ) );
  mux2_1 U13079 ( .ip1(n11651), .ip2(\CORTEXM0DS_INST/cm0_r12 [7]), .s(n11605), 
        .op(\CORTEXM0DS_INST/u_logic/Aslvx4 ) );
  mux2_1 U13080 ( .ip1(n11652), .ip2(\CORTEXM0DS_INST/cm0_r12 [28]), .s(n11605), .op(\CORTEXM0DS_INST/u_logic/Hslvx4 ) );
  mux2_1 U13081 ( .ip1(n11654), .ip2(\CORTEXM0DS_INST/cm0_r12 [31]), .s(n11605), .op(\CORTEXM0DS_INST/u_logic/Oslvx4 ) );
  inv_1 U13082 ( .ip(n11542), .op(n11600) );
  nand2_1 U13083 ( .ip1(n11600), .ip2(n11536), .op(n11550) );
  nand2_1 U13084 ( .ip1(n11538), .ip2(n11537), .op(n11608) );
  nor2_1 U13085 ( .ip1(n11550), .ip2(n11608), .op(n11539) );
  mux2_1 U13086 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [9]), .ip2(n11622), .s(n11539), 
        .op(\CORTEXM0DS_INST/u_logic/Ukivx4 ) );
  buf_1 U13087 ( .ip(n11539), .op(n11606) );
  mux2_1 U13088 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [2]), .ip2(n11623), .s(n11606), 
        .op(\CORTEXM0DS_INST/u_logic/Jpivx4 ) );
  mux2_1 U13089 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [10]), .ip2(n11624), .s(n11539), .op(\CORTEXM0DS_INST/u_logic/Ytivx4 ) );
  mux2_1 U13090 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [11]), .ip2(n11625), .s(n11606), .op(\CORTEXM0DS_INST/u_logic/Nyivx4 ) );
  mux2_1 U13091 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [12]), .ip2(n11626), .s(n11539), .op(\CORTEXM0DS_INST/u_logic/C3jvx4 ) );
  mux2_1 U13092 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [13]), .ip2(n11627), .s(n11606), .op(\CORTEXM0DS_INST/u_logic/R7jvx4 ) );
  mux2_1 U13093 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [14]), .ip2(n11628), .s(n11539), .op(\CORTEXM0DS_INST/u_logic/Gcjvx4 ) );
  mux2_1 U13094 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [16]), .ip2(n11629), .s(n11606), .op(\CORTEXM0DS_INST/u_logic/Vgjvx4 ) );
  mux2_1 U13095 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [17]), .ip2(n11630), .s(n11539), .op(\CORTEXM0DS_INST/u_logic/Kljvx4 ) );
  mux2_1 U13096 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [18]), .ip2(n11631), .s(n11606), .op(\CORTEXM0DS_INST/u_logic/Zpjvx4 ) );
  mux2_1 U13097 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [19]), .ip2(n11632), .s(n11539), .op(\CORTEXM0DS_INST/u_logic/Oujvx4 ) );
  mux2_1 U13098 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [20]), .ip2(n11633), .s(n11606), .op(\CORTEXM0DS_INST/u_logic/Dzjvx4 ) );
  mux2_1 U13099 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [21]), .ip2(n11634), .s(n11539), .op(\CORTEXM0DS_INST/u_logic/S3kvx4 ) );
  mux2_1 U13100 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [22]), .ip2(n11635), .s(n11539), .op(\CORTEXM0DS_INST/u_logic/H8kvx4 ) );
  mux2_1 U13101 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [3]), .ip2(n11636), .s(n11539), 
        .op(\CORTEXM0DS_INST/u_logic/Ddkvx4 ) );
  mux2_1 U13102 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [4]), .ip2(n11637), .s(n11539), 
        .op(\CORTEXM0DS_INST/u_logic/Shkvx4 ) );
  mux2_1 U13103 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [5]), .ip2(n11638), .s(n11539), 
        .op(\CORTEXM0DS_INST/u_logic/Hmkvx4 ) );
  mux2_1 U13104 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [6]), .ip2(n11639), .s(n11539), 
        .op(\CORTEXM0DS_INST/u_logic/Wqkvx4 ) );
  mux2_1 U13105 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [24]), .ip2(n11640), .s(n11539), .op(\CORTEXM0DS_INST/u_logic/Lvkvx4 ) );
  mux2_1 U13106 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [25]), .ip2(n11641), .s(n11606), .op(\CORTEXM0DS_INST/u_logic/Tzkvx4 ) );
  mux2_1 U13107 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [26]), .ip2(n11642), .s(n11539), .op(\CORTEXM0DS_INST/u_logic/I4lvx4 ) );
  mux2_1 U13108 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [27]), .ip2(n11644), .s(n11606), .op(\CORTEXM0DS_INST/u_logic/X8lvx4 ) );
  mux2_1 U13109 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [29]), .ip2(n11647), .s(n11539), .op(\CORTEXM0DS_INST/u_logic/Mdlvx4 ) );
  mux2_1 U13110 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [30]), .ip2(n11648), .s(n11606), .op(\CORTEXM0DS_INST/u_logic/Iilvx4 ) );
  mux2_1 U13111 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [0]), .ip2(n11649), .s(n11539), 
        .op(\CORTEXM0DS_INST/u_logic/Dqlvx4 ) );
  mux2_1 U13112 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [1]), .ip2(n11650), .s(n11606), 
        .op(\CORTEXM0DS_INST/u_logic/Kqlvx4 ) );
  mux2_1 U13113 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [7]), .ip2(n11651), .s(n11606), 
        .op(\CORTEXM0DS_INST/u_logic/Rqlvx4 ) );
  mux2_1 U13114 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [28]), .ip2(n11652), .s(n11606), .op(\CORTEXM0DS_INST/u_logic/Yqlvx4 ) );
  mux2_1 U13115 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [31]), .ip2(n11654), .s(n11606), .op(\CORTEXM0DS_INST/u_logic/Frlvx4 ) );
  inv_1 U13116 ( .ip(n11540), .op(n11552) );
  nor2_1 U13117 ( .ip1(n11552), .ip2(n11608), .op(n11541) );
  mux2_1 U13118 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [9]), .ip2(n11622), .s(n11541), 
        .op(\CORTEXM0DS_INST/u_logic/Gkivx4 ) );
  buf_1 U13119 ( .ip(n11541), .op(n11611) );
  mux2_1 U13120 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [2]), .ip2(n11623), .s(n11611), 
        .op(\CORTEXM0DS_INST/u_logic/Voivx4 ) );
  mux2_1 U13121 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [10]), .ip2(n11624), .s(n11541), .op(\CORTEXM0DS_INST/u_logic/Ktivx4 ) );
  mux2_1 U13122 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [11]), .ip2(n11625), .s(n11611), .op(\CORTEXM0DS_INST/u_logic/Zxivx4 ) );
  mux2_1 U13123 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [12]), .ip2(n11626), .s(n11541), .op(\CORTEXM0DS_INST/u_logic/O2jvx4 ) );
  mux2_1 U13124 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [13]), .ip2(n11627), .s(n11611), .op(\CORTEXM0DS_INST/u_logic/D7jvx4 ) );
  mux2_1 U13125 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [14]), .ip2(n11628), .s(n11541), .op(\CORTEXM0DS_INST/u_logic/Sbjvx4 ) );
  mux2_1 U13126 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [16]), .ip2(n11629), .s(n11611), .op(\CORTEXM0DS_INST/u_logic/Hgjvx4 ) );
  mux2_1 U13127 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [17]), .ip2(n11630), .s(n11541), .op(\CORTEXM0DS_INST/u_logic/Wkjvx4 ) );
  mux2_1 U13128 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [18]), .ip2(n11631), .s(n11611), .op(\CORTEXM0DS_INST/u_logic/Lpjvx4 ) );
  mux2_1 U13129 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [19]), .ip2(n11632), .s(n11541), .op(\CORTEXM0DS_INST/u_logic/Aujvx4 ) );
  mux2_1 U13130 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [20]), .ip2(n11633), .s(n11611), .op(\CORTEXM0DS_INST/u_logic/Pyjvx4 ) );
  mux2_1 U13131 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [21]), .ip2(n11634), .s(n11541), .op(\CORTEXM0DS_INST/u_logic/E3kvx4 ) );
  mux2_1 U13132 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [22]), .ip2(n11635), .s(n11541), .op(\CORTEXM0DS_INST/u_logic/T7kvx4 ) );
  mux2_1 U13133 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [3]), .ip2(n11636), .s(n11541), 
        .op(\CORTEXM0DS_INST/u_logic/Pckvx4 ) );
  mux2_1 U13134 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [4]), .ip2(n11637), .s(n11541), 
        .op(\CORTEXM0DS_INST/u_logic/Ehkvx4 ) );
  mux2_1 U13135 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [5]), .ip2(n11638), .s(n11541), 
        .op(\CORTEXM0DS_INST/u_logic/Tlkvx4 ) );
  mux2_1 U13136 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [6]), .ip2(n11639), .s(n11541), 
        .op(\CORTEXM0DS_INST/u_logic/Iqkvx4 ) );
  mux2_1 U13137 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [24]), .ip2(n11640), .s(n11541), .op(\CORTEXM0DS_INST/u_logic/Xukvx4 ) );
  mux2_1 U13138 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [25]), .ip2(n11641), .s(n11611), .op(\CORTEXM0DS_INST/u_logic/Fzkvx4 ) );
  mux2_1 U13139 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [26]), .ip2(n11642), .s(n11541), .op(\CORTEXM0DS_INST/u_logic/U3lvx4 ) );
  mux2_1 U13140 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [27]), .ip2(n11644), .s(n11611), .op(\CORTEXM0DS_INST/u_logic/J8lvx4 ) );
  mux2_1 U13141 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [29]), .ip2(n11647), .s(n11541), .op(\CORTEXM0DS_INST/u_logic/Yclvx4 ) );
  mux2_1 U13142 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [30]), .ip2(n11648), .s(n11611), .op(\CORTEXM0DS_INST/u_logic/Uhlvx4 ) );
  mux2_1 U13143 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [0]), .ip2(n11649), .s(n11541), 
        .op(\CORTEXM0DS_INST/u_logic/Lnlvx4 ) );
  mux2_1 U13144 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [1]), .ip2(n11650), .s(n11611), 
        .op(\CORTEXM0DS_INST/u_logic/Snlvx4 ) );
  mux2_1 U13145 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [7]), .ip2(n11651), .s(n11611), 
        .op(\CORTEXM0DS_INST/u_logic/Znlvx4 ) );
  mux2_1 U13146 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [28]), .ip2(n11652), .s(n11611), .op(\CORTEXM0DS_INST/u_logic/Golvx4 ) );
  mux2_1 U13147 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [31]), .ip2(n11654), .s(n11611), .op(\CORTEXM0DS_INST/u_logic/Nolvx4 ) );
  nand2_1 U13148 ( .ip1(n11542), .ip2(n11601), .op(n11554) );
  nor2_1 U13149 ( .ip1(n11554), .ip2(n11608), .op(n11543) );
  mux2_1 U13150 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [9]), .ip2(n11622), .s(n11543), 
        .op(\CORTEXM0DS_INST/u_logic/Zjivx4 ) );
  buf_1 U13151 ( .ip(n11543), .op(n11612) );
  mux2_1 U13152 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [2]), .ip2(n11623), .s(n11612), 
        .op(\CORTEXM0DS_INST/u_logic/Ooivx4 ) );
  mux2_1 U13153 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [10]), .ip2(n11624), .s(n11543), .op(\CORTEXM0DS_INST/u_logic/Dtivx4 ) );
  mux2_1 U13154 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [11]), .ip2(n11625), .s(n11612), .op(\CORTEXM0DS_INST/u_logic/Sxivx4 ) );
  mux2_1 U13155 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [12]), .ip2(n11626), .s(n11543), .op(\CORTEXM0DS_INST/u_logic/H2jvx4 ) );
  mux2_1 U13156 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [13]), .ip2(n11627), .s(n11612), .op(\CORTEXM0DS_INST/u_logic/W6jvx4 ) );
  mux2_1 U13157 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [14]), .ip2(n11628), .s(n11543), .op(\CORTEXM0DS_INST/u_logic/Lbjvx4 ) );
  mux2_1 U13158 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [16]), .ip2(n11629), .s(n11612), .op(\CORTEXM0DS_INST/u_logic/Agjvx4 ) );
  mux2_1 U13159 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [17]), .ip2(n11630), .s(n11543), .op(\CORTEXM0DS_INST/u_logic/Pkjvx4 ) );
  mux2_1 U13160 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [18]), .ip2(n11631), .s(n11612), .op(\CORTEXM0DS_INST/u_logic/Epjvx4 ) );
  mux2_1 U13161 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [19]), .ip2(n11632), .s(n11543), .op(\CORTEXM0DS_INST/u_logic/Ttjvx4 ) );
  mux2_1 U13162 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [20]), .ip2(n11633), .s(n11612), .op(\CORTEXM0DS_INST/u_logic/Iyjvx4 ) );
  mux2_1 U13163 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [21]), .ip2(n11634), .s(n11543), .op(\CORTEXM0DS_INST/u_logic/X2kvx4 ) );
  mux2_1 U13164 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [22]), .ip2(n11635), .s(n11543), .op(\CORTEXM0DS_INST/u_logic/M7kvx4 ) );
  mux2_1 U13165 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [3]), .ip2(n11636), .s(n11543), 
        .op(\CORTEXM0DS_INST/u_logic/Ickvx4 ) );
  mux2_1 U13166 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [4]), .ip2(n11637), .s(n11543), 
        .op(\CORTEXM0DS_INST/u_logic/Xgkvx4 ) );
  mux2_1 U13167 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [5]), .ip2(n11638), .s(n11543), 
        .op(\CORTEXM0DS_INST/u_logic/Mlkvx4 ) );
  mux2_1 U13168 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [6]), .ip2(n11639), .s(n11543), 
        .op(\CORTEXM0DS_INST/u_logic/Bqkvx4 ) );
  mux2_1 U13169 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [24]), .ip2(n11640), .s(n11543), .op(\CORTEXM0DS_INST/u_logic/Qukvx4 ) );
  mux2_1 U13170 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [25]), .ip2(n11641), .s(n11612), .op(\CORTEXM0DS_INST/u_logic/Yykvx4 ) );
  mux2_1 U13171 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [26]), .ip2(n11642), .s(n11543), .op(\CORTEXM0DS_INST/u_logic/N3lvx4 ) );
  mux2_1 U13172 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [27]), .ip2(n11644), .s(n11612), .op(\CORTEXM0DS_INST/u_logic/C8lvx4 ) );
  mux2_1 U13173 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [29]), .ip2(n11647), .s(n11543), .op(\CORTEXM0DS_INST/u_logic/Rclvx4 ) );
  mux2_1 U13174 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [30]), .ip2(n11648), .s(n11612), .op(\CORTEXM0DS_INST/u_logic/Nhlvx4 ) );
  mux2_1 U13175 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [0]), .ip2(n11649), .s(n11543), 
        .op(\CORTEXM0DS_INST/u_logic/Cmlvx4 ) );
  mux2_1 U13176 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [1]), .ip2(n11650), .s(n11612), 
        .op(\CORTEXM0DS_INST/u_logic/Jmlvx4 ) );
  mux2_1 U13177 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [7]), .ip2(n11651), .s(n11612), 
        .op(\CORTEXM0DS_INST/u_logic/Qmlvx4 ) );
  mux2_1 U13178 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [28]), .ip2(n11652), .s(n11612), .op(\CORTEXM0DS_INST/u_logic/Xmlvx4 ) );
  mux2_1 U13179 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [31]), .ip2(n11654), .s(n11612), .op(\CORTEXM0DS_INST/u_logic/Enlvx4 ) );
  nand2_1 U13180 ( .ip1(n11549), .ip2(n11547), .op(n11614) );
  nor2_1 U13181 ( .ip1(n11550), .ip2(n11614), .op(n11544) );
  mux2_1 U13182 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [9]), .ip2(n11622), .s(n11544), 
        .op(\CORTEXM0DS_INST/u_logic/Sjivx4 ) );
  buf_1 U13183 ( .ip(n11544), .op(n11613) );
  mux2_1 U13184 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [2]), .ip2(n11623), .s(n11613), 
        .op(\CORTEXM0DS_INST/u_logic/Hoivx4 ) );
  mux2_1 U13185 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [10]), .ip2(n11624), .s(n11544), .op(\CORTEXM0DS_INST/u_logic/Wsivx4 ) );
  mux2_1 U13186 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [11]), .ip2(n11625), .s(n11613), .op(\CORTEXM0DS_INST/u_logic/Lxivx4 ) );
  mux2_1 U13187 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [12]), .ip2(n11626), .s(n11544), .op(\CORTEXM0DS_INST/u_logic/A2jvx4 ) );
  mux2_1 U13188 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [13]), .ip2(n11627), .s(n11613), .op(\CORTEXM0DS_INST/u_logic/P6jvx4 ) );
  mux2_1 U13189 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [14]), .ip2(n11628), .s(n11544), .op(\CORTEXM0DS_INST/u_logic/Ebjvx4 ) );
  mux2_1 U13190 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [16]), .ip2(n11629), .s(n11613), .op(\CORTEXM0DS_INST/u_logic/Tfjvx4 ) );
  mux2_1 U13191 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [17]), .ip2(n11630), .s(n11544), .op(\CORTEXM0DS_INST/u_logic/Ikjvx4 ) );
  mux2_1 U13192 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [18]), .ip2(n11631), .s(n11613), .op(\CORTEXM0DS_INST/u_logic/Xojvx4 ) );
  mux2_1 U13193 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [19]), .ip2(n11632), .s(n11544), .op(\CORTEXM0DS_INST/u_logic/Mtjvx4 ) );
  mux2_1 U13194 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [20]), .ip2(n11633), .s(n11613), .op(\CORTEXM0DS_INST/u_logic/Byjvx4 ) );
  mux2_1 U13195 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [21]), .ip2(n11634), .s(n11544), .op(\CORTEXM0DS_INST/u_logic/Q2kvx4 ) );
  mux2_1 U13196 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [22]), .ip2(n11635), .s(n11544), .op(\CORTEXM0DS_INST/u_logic/F7kvx4 ) );
  mux2_1 U13197 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [3]), .ip2(n11636), .s(n11544), 
        .op(\CORTEXM0DS_INST/u_logic/Bckvx4 ) );
  mux2_1 U13198 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [4]), .ip2(n11637), .s(n11544), 
        .op(\CORTEXM0DS_INST/u_logic/Qgkvx4 ) );
  mux2_1 U13199 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [5]), .ip2(n11638), .s(n11544), 
        .op(\CORTEXM0DS_INST/u_logic/Flkvx4 ) );
  mux2_1 U13200 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [6]), .ip2(n11639), .s(n11544), 
        .op(\CORTEXM0DS_INST/u_logic/Upkvx4 ) );
  mux2_1 U13201 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [24]), .ip2(n11640), .s(n11544), .op(\CORTEXM0DS_INST/u_logic/Jukvx4 ) );
  mux2_1 U13202 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [25]), .ip2(n11641), .s(n11613), .op(\CORTEXM0DS_INST/u_logic/Rykvx4 ) );
  mux2_1 U13203 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [26]), .ip2(n11642), .s(n11544), .op(\CORTEXM0DS_INST/u_logic/G3lvx4 ) );
  mux2_1 U13204 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [27]), .ip2(n11644), .s(n11613), .op(\CORTEXM0DS_INST/u_logic/V7lvx4 ) );
  mux2_1 U13205 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [29]), .ip2(n11647), .s(n11544), .op(\CORTEXM0DS_INST/u_logic/Kclvx4 ) );
  mux2_1 U13206 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [30]), .ip2(n11648), .s(n11613), .op(\CORTEXM0DS_INST/u_logic/Ghlvx4 ) );
  mux2_1 U13207 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [0]), .ip2(n11649), .s(n11544), 
        .op(\CORTEXM0DS_INST/u_logic/Eulvx4 ) );
  mux2_1 U13208 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [1]), .ip2(n11650), .s(n11613), 
        .op(\CORTEXM0DS_INST/u_logic/Lulvx4 ) );
  mux2_1 U13209 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [7]), .ip2(n11651), .s(n11613), 
        .op(\CORTEXM0DS_INST/u_logic/Sulvx4 ) );
  mux2_1 U13210 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [28]), .ip2(n11652), .s(n11613), .op(\CORTEXM0DS_INST/u_logic/Zulvx4 ) );
  mux2_1 U13211 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [31]), .ip2(n11654), .s(n11613), .op(\CORTEXM0DS_INST/u_logic/Gvlvx4 ) );
  nor2_1 U13212 ( .ip1(n11552), .ip2(n11614), .op(n11545) );
  mux2_1 U13213 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [9]), .ip2(n11622), .s(n11545), 
        .op(\CORTEXM0DS_INST/u_logic/Ejivx4 ) );
  buf_1 U13214 ( .ip(n11545), .op(n11617) );
  mux2_1 U13215 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [2]), .ip2(n11623), .s(n11617), 
        .op(\CORTEXM0DS_INST/u_logic/Tnivx4 ) );
  mux2_1 U13216 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [10]), .ip2(n11624), .s(n11545), .op(\CORTEXM0DS_INST/u_logic/Isivx4 ) );
  mux2_1 U13217 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [11]), .ip2(n11625), .s(n11617), .op(\CORTEXM0DS_INST/u_logic/Xwivx4 ) );
  mux2_1 U13218 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [12]), .ip2(n11626), .s(n11545), .op(\CORTEXM0DS_INST/u_logic/M1jvx4 ) );
  mux2_1 U13219 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [13]), .ip2(n11627), .s(n11617), .op(\CORTEXM0DS_INST/u_logic/B6jvx4 ) );
  mux2_1 U13220 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [14]), .ip2(n11628), .s(n11545), .op(\CORTEXM0DS_INST/u_logic/Qajvx4 ) );
  mux2_1 U13221 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [16]), .ip2(n11629), .s(n11617), .op(\CORTEXM0DS_INST/u_logic/Ffjvx4 ) );
  mux2_1 U13222 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [17]), .ip2(n11630), .s(n11545), .op(\CORTEXM0DS_INST/u_logic/Ujjvx4 ) );
  mux2_1 U13223 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [18]), .ip2(n11631), .s(n11617), .op(\CORTEXM0DS_INST/u_logic/Jojvx4 ) );
  mux2_1 U13224 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [19]), .ip2(n11632), .s(n11545), .op(\CORTEXM0DS_INST/u_logic/Ysjvx4 ) );
  mux2_1 U13225 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [20]), .ip2(n11633), .s(n11617), .op(\CORTEXM0DS_INST/u_logic/Nxjvx4 ) );
  mux2_1 U13226 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [21]), .ip2(n11634), .s(n11545), .op(\CORTEXM0DS_INST/u_logic/C2kvx4 ) );
  mux2_1 U13227 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [22]), .ip2(n11635), .s(n11545), .op(\CORTEXM0DS_INST/u_logic/R6kvx4 ) );
  mux2_1 U13228 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [3]), .ip2(n11636), .s(n11545), 
        .op(\CORTEXM0DS_INST/u_logic/Nbkvx4 ) );
  mux2_1 U13229 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [4]), .ip2(n11637), .s(n11545), 
        .op(\CORTEXM0DS_INST/u_logic/Cgkvx4 ) );
  mux2_1 U13230 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [5]), .ip2(n11638), .s(n11545), 
        .op(\CORTEXM0DS_INST/u_logic/Rkkvx4 ) );
  mux2_1 U13231 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [6]), .ip2(n11639), .s(n11545), 
        .op(\CORTEXM0DS_INST/u_logic/Gpkvx4 ) );
  mux2_1 U13232 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [24]), .ip2(n11640), .s(n11545), .op(\CORTEXM0DS_INST/u_logic/Vtkvx4 ) );
  mux2_1 U13233 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [25]), .ip2(n11641), .s(n11617), .op(\CORTEXM0DS_INST/u_logic/Dykvx4 ) );
  mux2_1 U13234 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [26]), .ip2(n11642), .s(n11545), .op(\CORTEXM0DS_INST/u_logic/S2lvx4 ) );
  mux2_1 U13235 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [27]), .ip2(n11644), .s(n11617), .op(\CORTEXM0DS_INST/u_logic/H7lvx4 ) );
  mux2_1 U13236 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [29]), .ip2(n11647), .s(n11545), .op(\CORTEXM0DS_INST/u_logic/Wblvx4 ) );
  mux2_1 U13237 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [30]), .ip2(n11648), .s(n11617), .op(\CORTEXM0DS_INST/u_logic/Sglvx4 ) );
  mux2_1 U13238 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [0]), .ip2(n11649), .s(n11545), 
        .op(\CORTEXM0DS_INST/u_logic/Wwlvx4 ) );
  mux2_1 U13239 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [1]), .ip2(n11650), .s(n11617), 
        .op(\CORTEXM0DS_INST/u_logic/Dxlvx4 ) );
  mux2_1 U13240 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [7]), .ip2(n11651), .s(n11617), 
        .op(\CORTEXM0DS_INST/u_logic/Kxlvx4 ) );
  mux2_1 U13241 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [28]), .ip2(n11652), .s(n11617), .op(\CORTEXM0DS_INST/u_logic/Rxlvx4 ) );
  mux2_1 U13242 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [31]), .ip2(n11654), .s(n11617), .op(\CORTEXM0DS_INST/u_logic/Yxlvx4 ) );
  nor2_1 U13243 ( .ip1(n11554), .ip2(n11614), .op(n11546) );
  mux2_1 U13244 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [9]), .ip2(n11622), .s(n11546), 
        .op(\CORTEXM0DS_INST/u_logic/Xiivx4 ) );
  buf_1 U13245 ( .ip(n11546), .op(n11618) );
  mux2_1 U13246 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [2]), .ip2(n11623), .s(n11618), 
        .op(\CORTEXM0DS_INST/u_logic/Mnivx4 ) );
  mux2_1 U13247 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [10]), .ip2(n11624), .s(n11546), .op(\CORTEXM0DS_INST/u_logic/Bsivx4 ) );
  mux2_1 U13248 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [11]), .ip2(n11625), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/Qwivx4 ) );
  mux2_1 U13249 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [12]), .ip2(n11626), .s(n11546), .op(\CORTEXM0DS_INST/u_logic/F1jvx4 ) );
  mux2_1 U13250 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [13]), .ip2(n11627), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/U5jvx4 ) );
  mux2_1 U13251 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [14]), .ip2(n11628), .s(n11546), .op(\CORTEXM0DS_INST/u_logic/Jajvx4 ) );
  mux2_1 U13252 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [16]), .ip2(n11629), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/Yejvx4 ) );
  mux2_1 U13253 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [17]), .ip2(n11630), .s(n11546), .op(\CORTEXM0DS_INST/u_logic/Njjvx4 ) );
  mux2_1 U13254 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [18]), .ip2(n11631), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/Cojvx4 ) );
  mux2_1 U13255 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [19]), .ip2(n11632), .s(n11546), .op(\CORTEXM0DS_INST/u_logic/Rsjvx4 ) );
  mux2_1 U13256 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [20]), .ip2(n11633), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/Gxjvx4 ) );
  mux2_1 U13257 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [21]), .ip2(n11634), .s(n11546), .op(\CORTEXM0DS_INST/u_logic/V1kvx4 ) );
  mux2_1 U13258 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [22]), .ip2(n11635), .s(n11546), .op(\CORTEXM0DS_INST/u_logic/K6kvx4 ) );
  mux2_1 U13259 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [3]), .ip2(n11636), .s(n11546), 
        .op(\CORTEXM0DS_INST/u_logic/Gbkvx4 ) );
  mux2_1 U13260 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [4]), .ip2(n11637), .s(n11546), 
        .op(\CORTEXM0DS_INST/u_logic/Vfkvx4 ) );
  mux2_1 U13261 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [5]), .ip2(n11638), .s(n11546), 
        .op(\CORTEXM0DS_INST/u_logic/Kkkvx4 ) );
  mux2_1 U13262 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [6]), .ip2(n11639), .s(n11546), 
        .op(\CORTEXM0DS_INST/u_logic/Zokvx4 ) );
  mux2_1 U13263 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [24]), .ip2(n11640), .s(n11546), .op(\CORTEXM0DS_INST/u_logic/Otkvx4 ) );
  mux2_1 U13264 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [25]), .ip2(n11641), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/Wxkvx4 ) );
  mux2_1 U13265 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [26]), .ip2(n11642), .s(n11546), .op(\CORTEXM0DS_INST/u_logic/L2lvx4 ) );
  mux2_1 U13266 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [27]), .ip2(n11644), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/A7lvx4 ) );
  mux2_1 U13267 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [29]), .ip2(n11647), .s(n11546), .op(\CORTEXM0DS_INST/u_logic/Pblvx4 ) );
  mux2_1 U13268 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [30]), .ip2(n11648), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/Lglvx4 ) );
  mux2_1 U13269 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [0]), .ip2(n11649), .s(n11546), 
        .op(\CORTEXM0DS_INST/u_logic/Fylvx4 ) );
  mux2_1 U13270 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [1]), .ip2(n11650), .s(n11618), 
        .op(\CORTEXM0DS_INST/u_logic/Mylvx4 ) );
  mux2_1 U13271 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [7]), .ip2(n11651), .s(n11618), 
        .op(\CORTEXM0DS_INST/u_logic/Tylvx4 ) );
  mux2_1 U13272 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [28]), .ip2(n11652), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/Azlvx4 ) );
  mux2_1 U13273 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [31]), .ip2(n11654), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/Hzlvx4 ) );
  inv_1 U13274 ( .ip(n11547), .op(n11548) );
  nand2_1 U13275 ( .ip1(n11549), .ip2(n11548), .op(n11621) );
  nor2_1 U13276 ( .ip1(n11550), .ip2(n11621), .op(n11551) );
  mux2_1 U13277 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [9]), .ip2(n11622), .s(n11551), 
        .op(\CORTEXM0DS_INST/u_logic/Qiivx4 ) );
  buf_1 U13278 ( .ip(n11551), .op(n11619) );
  mux2_1 U13279 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [2]), .ip2(n11623), .s(n11619), 
        .op(\CORTEXM0DS_INST/u_logic/Fnivx4 ) );
  mux2_1 U13280 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [10]), .ip2(n11624), .s(n11551), .op(\CORTEXM0DS_INST/u_logic/Urivx4 ) );
  mux2_1 U13281 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [11]), .ip2(n11625), .s(n11619), .op(\CORTEXM0DS_INST/u_logic/Jwivx4 ) );
  mux2_1 U13282 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [12]), .ip2(n11626), .s(n11551), .op(\CORTEXM0DS_INST/u_logic/Y0jvx4 ) );
  mux2_1 U13283 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [13]), .ip2(n11627), .s(n11619), .op(\CORTEXM0DS_INST/u_logic/N5jvx4 ) );
  mux2_1 U13284 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [14]), .ip2(n11628), .s(n11551), .op(\CORTEXM0DS_INST/u_logic/Cajvx4 ) );
  mux2_1 U13285 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [16]), .ip2(n11629), .s(n11619), .op(\CORTEXM0DS_INST/u_logic/Rejvx4 ) );
  mux2_1 U13286 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [17]), .ip2(n11630), .s(n11551), .op(\CORTEXM0DS_INST/u_logic/Gjjvx4 ) );
  mux2_1 U13287 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [18]), .ip2(n11631), .s(n11619), .op(\CORTEXM0DS_INST/u_logic/Vnjvx4 ) );
  mux2_1 U13288 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [19]), .ip2(n11632), .s(n11551), .op(\CORTEXM0DS_INST/u_logic/Ksjvx4 ) );
  mux2_1 U13289 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [20]), .ip2(n11633), .s(n11619), .op(\CORTEXM0DS_INST/u_logic/Zwjvx4 ) );
  mux2_1 U13290 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [21]), .ip2(n11634), .s(n11551), .op(\CORTEXM0DS_INST/u_logic/O1kvx4 ) );
  mux2_1 U13291 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [22]), .ip2(n11635), .s(n11551), .op(\CORTEXM0DS_INST/u_logic/D6kvx4 ) );
  mux2_1 U13292 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [3]), .ip2(n11636), .s(n11551), 
        .op(\CORTEXM0DS_INST/u_logic/Zakvx4 ) );
  mux2_1 U13293 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [4]), .ip2(n11637), .s(n11551), 
        .op(\CORTEXM0DS_INST/u_logic/Ofkvx4 ) );
  mux2_1 U13294 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [5]), .ip2(n11638), .s(n11551), 
        .op(\CORTEXM0DS_INST/u_logic/Dkkvx4 ) );
  mux2_1 U13295 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [6]), .ip2(n11639), .s(n11551), 
        .op(\CORTEXM0DS_INST/u_logic/Sokvx4 ) );
  mux2_1 U13296 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [24]), .ip2(n11640), .s(n11551), .op(\CORTEXM0DS_INST/u_logic/Htkvx4 ) );
  mux2_1 U13297 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [25]), .ip2(n11641), .s(n11619), .op(\CORTEXM0DS_INST/u_logic/Pxkvx4 ) );
  mux2_1 U13298 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [26]), .ip2(n11642), .s(n11551), .op(\CORTEXM0DS_INST/u_logic/E2lvx4 ) );
  mux2_1 U13299 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [27]), .ip2(n11644), .s(n11619), .op(\CORTEXM0DS_INST/u_logic/T6lvx4 ) );
  mux2_1 U13300 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [29]), .ip2(n11647), .s(n11551), .op(\CORTEXM0DS_INST/u_logic/Iblvx4 ) );
  mux2_1 U13301 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [30]), .ip2(n11648), .s(n11619), .op(\CORTEXM0DS_INST/u_logic/Eglvx4 ) );
  mux2_1 U13302 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [0]), .ip2(n11649), .s(n11551), 
        .op(\CORTEXM0DS_INST/u_logic/Ozlvx4 ) );
  mux2_1 U13303 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [1]), .ip2(n11650), .s(n11619), 
        .op(\CORTEXM0DS_INST/u_logic/Vzlvx4 ) );
  mux2_1 U13304 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [7]), .ip2(n11651), .s(n11619), 
        .op(\CORTEXM0DS_INST/u_logic/C0mvx4 ) );
  mux2_1 U13305 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [28]), .ip2(n11652), .s(n11619), .op(\CORTEXM0DS_INST/u_logic/J0mvx4 ) );
  mux2_1 U13306 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [31]), .ip2(n11654), .s(n11619), .op(\CORTEXM0DS_INST/u_logic/Q0mvx4 ) );
  nor2_1 U13307 ( .ip1(n11552), .ip2(n11621), .op(n11553) );
  mux2_1 U13308 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [9]), .ip2(n11622), .s(n11553), 
        .op(\CORTEXM0DS_INST/u_logic/Ciivx4 ) );
  buf_1 U13309 ( .ip(n11553), .op(n11655) );
  mux2_1 U13310 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [2]), .ip2(n11623), .s(n11655), 
        .op(\CORTEXM0DS_INST/u_logic/Rmivx4 ) );
  mux2_1 U13311 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [10]), .ip2(n11624), .s(n11553), .op(\CORTEXM0DS_INST/u_logic/Grivx4 ) );
  mux2_1 U13312 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [11]), .ip2(n11625), .s(n11655), .op(\CORTEXM0DS_INST/u_logic/Vvivx4 ) );
  mux2_1 U13313 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [12]), .ip2(n11626), .s(n11553), .op(\CORTEXM0DS_INST/u_logic/K0jvx4 ) );
  mux2_1 U13314 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [13]), .ip2(n11627), .s(n11655), .op(\CORTEXM0DS_INST/u_logic/Z4jvx4 ) );
  mux2_1 U13315 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [14]), .ip2(n11628), .s(n11553), .op(\CORTEXM0DS_INST/u_logic/O9jvx4 ) );
  mux2_1 U13316 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [16]), .ip2(n11629), .s(n11655), .op(\CORTEXM0DS_INST/u_logic/Dejvx4 ) );
  mux2_1 U13317 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [17]), .ip2(n11630), .s(n11553), .op(\CORTEXM0DS_INST/u_logic/Sijvx4 ) );
  mux2_1 U13318 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [18]), .ip2(n11631), .s(n11655), .op(\CORTEXM0DS_INST/u_logic/Hnjvx4 ) );
  mux2_1 U13319 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [19]), .ip2(n11632), .s(n11553), .op(\CORTEXM0DS_INST/u_logic/Wrjvx4 ) );
  mux2_1 U13320 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [20]), .ip2(n11633), .s(n11655), .op(\CORTEXM0DS_INST/u_logic/Lwjvx4 ) );
  mux2_1 U13321 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [21]), .ip2(n11634), .s(n11553), .op(\CORTEXM0DS_INST/u_logic/A1kvx4 ) );
  mux2_1 U13322 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [22]), .ip2(n11635), .s(n11553), .op(\CORTEXM0DS_INST/u_logic/P5kvx4 ) );
  mux2_1 U13323 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [3]), .ip2(n11636), .s(n11553), 
        .op(\CORTEXM0DS_INST/u_logic/Lakvx4 ) );
  mux2_1 U13324 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [4]), .ip2(n11637), .s(n11553), 
        .op(\CORTEXM0DS_INST/u_logic/Afkvx4 ) );
  mux2_1 U13325 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [5]), .ip2(n11638), .s(n11553), 
        .op(\CORTEXM0DS_INST/u_logic/Pjkvx4 ) );
  mux2_1 U13326 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [6]), .ip2(n11639), .s(n11553), 
        .op(\CORTEXM0DS_INST/u_logic/Eokvx4 ) );
  mux2_1 U13327 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [24]), .ip2(n11640), .s(n11553), .op(\CORTEXM0DS_INST/u_logic/Tskvx4 ) );
  mux2_1 U13328 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [25]), .ip2(n11641), .s(n11655), .op(\CORTEXM0DS_INST/u_logic/Bxkvx4 ) );
  mux2_1 U13329 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [26]), .ip2(n11642), .s(n11553), .op(\CORTEXM0DS_INST/u_logic/Q1lvx4 ) );
  mux2_1 U13330 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [27]), .ip2(n11644), .s(n11655), .op(\CORTEXM0DS_INST/u_logic/F6lvx4 ) );
  mux2_1 U13331 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [29]), .ip2(n11647), .s(n11553), .op(\CORTEXM0DS_INST/u_logic/Ualvx4 ) );
  mux2_1 U13332 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [30]), .ip2(n11648), .s(n11655), .op(\CORTEXM0DS_INST/u_logic/Qflvx4 ) );
  mux2_1 U13333 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [0]), .ip2(n11649), .s(n11553), 
        .op(\CORTEXM0DS_INST/u_logic/Eenvx4 ) );
  mux2_1 U13334 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [1]), .ip2(n11650), .s(n11655), 
        .op(\CORTEXM0DS_INST/u_logic/Lenvx4 ) );
  mux2_1 U13335 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [7]), .ip2(n11651), .s(n11655), 
        .op(\CORTEXM0DS_INST/u_logic/Senvx4 ) );
  mux2_1 U13336 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [28]), .ip2(n11652), .s(n11655), .op(\CORTEXM0DS_INST/u_logic/Zenvx4 ) );
  mux2_1 U13337 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [31]), .ip2(n11654), .s(n11655), .op(\CORTEXM0DS_INST/u_logic/Gfnvx4 ) );
  nor2_1 U13338 ( .ip1(n11554), .ip2(n11621), .op(n11555) );
  mux2_1 U13339 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [9]), .ip2(n11622), .s(n11555), 
        .op(\CORTEXM0DS_INST/u_logic/Vhivx4 ) );
  buf_1 U13340 ( .ip(n11555), .op(n11658) );
  mux2_1 U13341 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [2]), .ip2(n11623), .s(n11658), 
        .op(\CORTEXM0DS_INST/u_logic/Kmivx4 ) );
  mux2_1 U13342 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [10]), .ip2(n11624), .s(n11555), .op(\CORTEXM0DS_INST/u_logic/Zqivx4 ) );
  mux2_1 U13343 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [11]), .ip2(n11625), .s(n11658), .op(\CORTEXM0DS_INST/u_logic/Ovivx4 ) );
  mux2_1 U13344 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [12]), .ip2(n11626), .s(n11555), .op(\CORTEXM0DS_INST/u_logic/D0jvx4 ) );
  mux2_1 U13345 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [13]), .ip2(n11627), .s(n11658), .op(\CORTEXM0DS_INST/u_logic/S4jvx4 ) );
  mux2_1 U13346 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [14]), .ip2(n11628), .s(n11555), .op(\CORTEXM0DS_INST/u_logic/H9jvx4 ) );
  mux2_1 U13347 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [16]), .ip2(n11629), .s(n11658), .op(\CORTEXM0DS_INST/u_logic/Wdjvx4 ) );
  mux2_1 U13348 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [17]), .ip2(n11630), .s(n11555), .op(\CORTEXM0DS_INST/u_logic/Lijvx4 ) );
  mux2_1 U13349 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [18]), .ip2(n11631), .s(n11658), .op(\CORTEXM0DS_INST/u_logic/Anjvx4 ) );
  mux2_1 U13350 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [19]), .ip2(n11632), .s(n11555), .op(\CORTEXM0DS_INST/u_logic/Prjvx4 ) );
  mux2_1 U13351 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [20]), .ip2(n11633), .s(n11658), .op(\CORTEXM0DS_INST/u_logic/Ewjvx4 ) );
  mux2_1 U13352 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [21]), .ip2(n11634), .s(n11555), .op(\CORTEXM0DS_INST/u_logic/T0kvx4 ) );
  mux2_1 U13353 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [22]), .ip2(n11635), .s(n11555), .op(\CORTEXM0DS_INST/u_logic/I5kvx4 ) );
  mux2_1 U13354 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [3]), .ip2(n11636), .s(n11555), 
        .op(\CORTEXM0DS_INST/u_logic/Eakvx4 ) );
  mux2_1 U13355 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [4]), .ip2(n11637), .s(n11555), 
        .op(\CORTEXM0DS_INST/u_logic/Tekvx4 ) );
  mux2_1 U13356 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [5]), .ip2(n11638), .s(n11555), 
        .op(\CORTEXM0DS_INST/u_logic/Ijkvx4 ) );
  mux2_1 U13357 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [6]), .ip2(n11639), .s(n11555), 
        .op(\CORTEXM0DS_INST/u_logic/Xnkvx4 ) );
  mux2_1 U13358 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [24]), .ip2(n11640), .s(n11555), .op(\CORTEXM0DS_INST/u_logic/Mskvx4 ) );
  mux2_1 U13359 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [25]), .ip2(n11641), .s(n11658), .op(\CORTEXM0DS_INST/u_logic/Uwkvx4 ) );
  mux2_1 U13360 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [26]), .ip2(n11642), .s(n11555), .op(\CORTEXM0DS_INST/u_logic/J1lvx4 ) );
  mux2_1 U13361 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [27]), .ip2(n11644), .s(n11658), .op(\CORTEXM0DS_INST/u_logic/Y5lvx4 ) );
  mux2_1 U13362 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [29]), .ip2(n11647), .s(n11555), .op(\CORTEXM0DS_INST/u_logic/Nalvx4 ) );
  mux2_1 U13363 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [30]), .ip2(n11648), .s(n11658), .op(\CORTEXM0DS_INST/u_logic/Jflvx4 ) );
  mux2_1 U13364 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [0]), .ip2(n11649), .s(n11555), 
        .op(\CORTEXM0DS_INST/u_logic/Bgnvx4 ) );
  mux2_1 U13365 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [7]), .ip2(n11651), .s(n11658), 
        .op(\CORTEXM0DS_INST/u_logic/Ignvx4 ) );
  mux2_1 U13366 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [31]), .ip2(n11654), .s(n11658), .op(\CORTEXM0DS_INST/u_logic/Wgnvx4 ) );
  mux2_1 U13367 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [28]), .ip2(n11652), .s(n11658), .op(\CORTEXM0DS_INST/u_logic/Dhnvx4 ) );
  mux2_1 U13368 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [1]), .ip2(n11650), .s(n11658), 
        .op(\CORTEXM0DS_INST/u_logic/Minvx4 ) );
  nand2_1 U13369 ( .ip1(n11556), .ip2(n11578), .op(n11569) );
  nor2_1 U13370 ( .ip1(n11588), .ip2(n11557), .op(n11563) );
  or2_1 U13371 ( .ip1(n11558), .ip2(n12158), .op(n11561) );
  or2_1 U13372 ( .ip1(n11559), .ip2(n12158), .op(n11560) );
  nand2_1 U13373 ( .ip1(n11561), .ip2(n11560), .op(n11562) );
  not_ab_or_c_or_d U13374 ( .ip1(n11565), .ip2(n11564), .ip3(n11563), .ip4(
        n11562), .op(n11566) );
  not_ab_or_c_or_d U13375 ( .ip1(n11594), .ip2(n12661), .ip3(n11593), .ip4(
        n11566), .op(n11568) );
  nand3_1 U13376 ( .ip1(n11569), .ip2(n11568), .ip3(n11567), .op(n11659) );
  nor2_1 U13377 ( .ip1(n11571), .ip2(n11570), .op(n11572) );
  mux2_1 U13378 ( .ip1(\CORTEXM0DS_INST/vis_psp [6]), .ip2(n11659), .s(n11572), 
        .op(\CORTEXM0DS_INST/u_logic/Hhivx4 ) );
  buf_1 U13379 ( .ip(n11572), .op(n11598) );
  mux2_1 U13380 ( .ip1(\CORTEXM0DS_INST/vis_psp [7]), .ip2(n11622), .s(n11598), 
        .op(\CORTEXM0DS_INST/u_logic/Wlivx4 ) );
  mux2_1 U13381 ( .ip1(\CORTEXM0DS_INST/vis_psp [0]), .ip2(n11623), .s(n11572), 
        .op(\CORTEXM0DS_INST/u_logic/Lqivx4 ) );
  mux2_1 U13382 ( .ip1(\CORTEXM0DS_INST/vis_psp [8]), .ip2(n11624), .s(n11598), 
        .op(\CORTEXM0DS_INST/u_logic/Avivx4 ) );
  mux2_1 U13383 ( .ip1(\CORTEXM0DS_INST/vis_psp [9]), .ip2(n11625), .s(n11572), 
        .op(\CORTEXM0DS_INST/u_logic/Pzivx4 ) );
  mux2_1 U13384 ( .ip1(\CORTEXM0DS_INST/vis_psp [10]), .ip2(n11626), .s(n11598), .op(\CORTEXM0DS_INST/u_logic/E4jvx4 ) );
  mux2_1 U13385 ( .ip1(\CORTEXM0DS_INST/vis_psp [11]), .ip2(n11627), .s(n11572), .op(\CORTEXM0DS_INST/u_logic/T8jvx4 ) );
  mux2_1 U13386 ( .ip1(\CORTEXM0DS_INST/vis_psp [12]), .ip2(n11628), .s(n11598), .op(\CORTEXM0DS_INST/u_logic/Idjvx4 ) );
  mux2_1 U13387 ( .ip1(\CORTEXM0DS_INST/vis_psp [14]), .ip2(n11629), .s(n11572), .op(\CORTEXM0DS_INST/u_logic/Xhjvx4 ) );
  mux2_1 U13388 ( .ip1(\CORTEXM0DS_INST/vis_psp [15]), .ip2(n11630), .s(n11598), .op(\CORTEXM0DS_INST/u_logic/Mmjvx4 ) );
  mux2_1 U13389 ( .ip1(\CORTEXM0DS_INST/vis_psp [16]), .ip2(n11631), .s(n11572), .op(\CORTEXM0DS_INST/u_logic/Brjvx4 ) );
  mux2_1 U13390 ( .ip1(\CORTEXM0DS_INST/vis_psp [17]), .ip2(n11632), .s(n11598), .op(\CORTEXM0DS_INST/u_logic/Qvjvx4 ) );
  mux2_1 U13391 ( .ip1(\CORTEXM0DS_INST/vis_psp [18]), .ip2(n11633), .s(n11572), .op(\CORTEXM0DS_INST/u_logic/F0kvx4 ) );
  mux2_1 U13392 ( .ip1(\CORTEXM0DS_INST/vis_psp [19]), .ip2(n11634), .s(n11572), .op(\CORTEXM0DS_INST/u_logic/U4kvx4 ) );
  mux2_1 U13393 ( .ip1(\CORTEXM0DS_INST/vis_psp [20]), .ip2(n11635), .s(n11572), .op(\CORTEXM0DS_INST/u_logic/J9kvx4 ) );
  mux2_1 U13394 ( .ip1(\CORTEXM0DS_INST/vis_psp [1]), .ip2(n11636), .s(n11572), 
        .op(\CORTEXM0DS_INST/u_logic/Fekvx4 ) );
  mux2_1 U13395 ( .ip1(\CORTEXM0DS_INST/vis_psp [2]), .ip2(n11637), .s(n11572), 
        .op(\CORTEXM0DS_INST/u_logic/Uikvx4 ) );
  mux2_1 U13396 ( .ip1(\CORTEXM0DS_INST/vis_psp [3]), .ip2(n11638), .s(n11598), 
        .op(\CORTEXM0DS_INST/u_logic/Jnkvx4 ) );
  mux2_1 U13397 ( .ip1(\CORTEXM0DS_INST/vis_psp [4]), .ip2(n11639), .s(n11572), 
        .op(\CORTEXM0DS_INST/u_logic/Yrkvx4 ) );
  mux2_1 U13398 ( .ip1(\CORTEXM0DS_INST/vis_psp [22]), .ip2(n11640), .s(n11598), .op(\CORTEXM0DS_INST/u_logic/Nwkvx4 ) );
  mux2_1 U13399 ( .ip1(\CORTEXM0DS_INST/vis_psp [23]), .ip2(n11641), .s(n11572), .op(\CORTEXM0DS_INST/u_logic/V0lvx4 ) );
  mux2_1 U13400 ( .ip1(\CORTEXM0DS_INST/vis_psp [24]), .ip2(n11642), .s(n11598), .op(\CORTEXM0DS_INST/u_logic/K5lvx4 ) );
  mux2_1 U13401 ( .ip1(\CORTEXM0DS_INST/vis_psp [25]), .ip2(n11644), .s(n11572), .op(\CORTEXM0DS_INST/u_logic/Z9lvx4 ) );
  mux2_1 U13402 ( .ip1(\CORTEXM0DS_INST/vis_psp [27]), .ip2(n11647), .s(n11598), .op(\CORTEXM0DS_INST/u_logic/Oelvx4 ) );
  mux2_1 U13403 ( .ip1(\CORTEXM0DS_INST/vis_psp [28]), .ip2(n11648), .s(n11572), .op(\CORTEXM0DS_INST/u_logic/Kjlvx4 ) );
  mux2_1 U13404 ( .ip1(\CORTEXM0DS_INST/vis_psp [29]), .ip2(n11654), .s(n11598), .op(\CORTEXM0DS_INST/u_logic/Mklvx4 ) );
  mux2_1 U13405 ( .ip1(\CORTEXM0DS_INST/vis_psp [26]), .ip2(n11652), .s(n11598), .op(\CORTEXM0DS_INST/u_logic/Tklvx4 ) );
  mux2_1 U13406 ( .ip1(\CORTEXM0DS_INST/vis_psp [5]), .ip2(n11651), .s(n11598), 
        .op(\CORTEXM0DS_INST/u_logic/Allvx4 ) );
  not_ab_or_c_or_d U13407 ( .ip1(n11594), .ip2(n12682), .ip3(n11574), .ip4(
        n11573), .op(n11576) );
  nand3_1 U13408 ( .ip1(n11577), .ip2(n11576), .ip3(n11575), .op(n11656) );
  mux2_1 U13409 ( .ip1(\CORTEXM0DS_INST/vis_psp [21]), .ip2(n11656), .s(n11598), .op(\CORTEXM0DS_INST/u_logic/D8ivx4 ) );
  nand2_1 U13410 ( .ip1(n11579), .ip2(n11578), .op(n11597) );
  or2_1 U13411 ( .ip1(n11581), .ip2(n11580), .op(n11582) );
  nand2_1 U13412 ( .ip1(n11589), .ip2(n11582), .op(n11584) );
  or2_1 U13413 ( .ip1(n11583), .ip2(n11584), .op(n11587) );
  or2_1 U13414 ( .ip1(n11585), .ip2(n11584), .op(n11586) );
  nand2_1 U13415 ( .ip1(n11587), .ip2(n11586), .op(n11591) );
  nor2_1 U13416 ( .ip1(n11589), .ip2(n11588), .op(n11590) );
  nor2_1 U13417 ( .ip1(n11591), .ip2(n11590), .op(n11592) );
  not_ab_or_c_or_d U13418 ( .ip1(n11594), .ip2(n12669), .ip3(n11593), .ip4(
        n11592), .op(n11596) );
  nand3_1 U13419 ( .ip1(n11597), .ip2(n11596), .ip3(n11595), .op(n11657) );
  mux2_1 U13420 ( .ip1(\CORTEXM0DS_INST/vis_psp [13]), .ip2(n11657), .s(n11598), .op(\CORTEXM0DS_INST/u_logic/Scivx4 ) );
  mux2_1 U13421 ( .ip1(\CORTEXM0DS_INST/vis_msp [21]), .ip2(n11656), .s(n11599), .op(\CORTEXM0DS_INST/u_logic/W7ivx4 ) );
  mux2_1 U13422 ( .ip1(\CORTEXM0DS_INST/vis_msp [13]), .ip2(n11657), .s(n11599), .op(\CORTEXM0DS_INST/u_logic/Lcivx4 ) );
  mux2_1 U13423 ( .ip1(\CORTEXM0DS_INST/vis_msp [6]), .ip2(n11659), .s(n11599), 
        .op(\CORTEXM0DS_INST/u_logic/Ahivx4 ) );
  nor2_1 U13424 ( .ip1(n11601), .ip2(n11600), .op(n11607) );
  nand2_1 U13425 ( .ip1(n11602), .ip2(n11607), .op(n11603) );
  mux2_1 U13426 ( .ip1(n11656), .ip2(\CORTEXM0DS_INST/cm0_r14 [23]), .s(n11603), .op(\CORTEXM0DS_INST/u_logic/P7ivx4 ) );
  buf_1 U13427 ( .ip(n11603), .op(n11604) );
  mux2_1 U13428 ( .ip1(n11657), .ip2(\CORTEXM0DS_INST/cm0_r14 [15]), .s(n11604), .op(\CORTEXM0DS_INST/u_logic/Ecivx4 ) );
  mux2_1 U13429 ( .ip1(n11659), .ip2(\CORTEXM0DS_INST/cm0_r14 [8]), .s(n11603), 
        .op(\CORTEXM0DS_INST/u_logic/Tgivx4 ) );
  mux2_1 U13430 ( .ip1(n11622), .ip2(\CORTEXM0DS_INST/cm0_r14 [9]), .s(n11604), 
        .op(\CORTEXM0DS_INST/u_logic/Ilivx4 ) );
  mux2_1 U13431 ( .ip1(n11623), .ip2(\CORTEXM0DS_INST/cm0_r14 [2]), .s(n11603), 
        .op(\CORTEXM0DS_INST/u_logic/Xpivx4 ) );
  mux2_1 U13432 ( .ip1(n11624), .ip2(\CORTEXM0DS_INST/cm0_r14 [10]), .s(n11604), .op(\CORTEXM0DS_INST/u_logic/Muivx4 ) );
  mux2_1 U13433 ( .ip1(n11625), .ip2(\CORTEXM0DS_INST/cm0_r14 [11]), .s(n11603), .op(\CORTEXM0DS_INST/u_logic/Bzivx4 ) );
  mux2_1 U13434 ( .ip1(n11626), .ip2(\CORTEXM0DS_INST/cm0_r14 [12]), .s(n11604), .op(\CORTEXM0DS_INST/u_logic/Q3jvx4 ) );
  mux2_1 U13435 ( .ip1(n11627), .ip2(\CORTEXM0DS_INST/cm0_r14 [13]), .s(n11603), .op(\CORTEXM0DS_INST/u_logic/F8jvx4 ) );
  mux2_1 U13436 ( .ip1(n11628), .ip2(\CORTEXM0DS_INST/cm0_r14 [14]), .s(n11604), .op(\CORTEXM0DS_INST/u_logic/Ucjvx4 ) );
  mux2_1 U13437 ( .ip1(n11629), .ip2(\CORTEXM0DS_INST/cm0_r14 [16]), .s(n11603), .op(\CORTEXM0DS_INST/u_logic/Jhjvx4 ) );
  mux2_1 U13438 ( .ip1(n11630), .ip2(\CORTEXM0DS_INST/cm0_r14 [17]), .s(n11604), .op(\CORTEXM0DS_INST/u_logic/Yljvx4 ) );
  mux2_1 U13439 ( .ip1(n11631), .ip2(\CORTEXM0DS_INST/cm0_r14 [18]), .s(n11603), .op(\CORTEXM0DS_INST/u_logic/Nqjvx4 ) );
  mux2_1 U13440 ( .ip1(n11632), .ip2(\CORTEXM0DS_INST/cm0_r14 [19]), .s(n11603), .op(\CORTEXM0DS_INST/u_logic/Cvjvx4 ) );
  mux2_1 U13441 ( .ip1(n11633), .ip2(\CORTEXM0DS_INST/cm0_r14 [20]), .s(n11603), .op(\CORTEXM0DS_INST/u_logic/Rzjvx4 ) );
  mux2_1 U13442 ( .ip1(n11634), .ip2(\CORTEXM0DS_INST/cm0_r14 [21]), .s(n11603), .op(\CORTEXM0DS_INST/u_logic/G4kvx4 ) );
  mux2_1 U13443 ( .ip1(n11635), .ip2(\CORTEXM0DS_INST/cm0_r14 [22]), .s(n11603), .op(\CORTEXM0DS_INST/u_logic/V8kvx4 ) );
  mux2_1 U13444 ( .ip1(n11636), .ip2(\CORTEXM0DS_INST/cm0_r14 [3]), .s(n11603), 
        .op(\CORTEXM0DS_INST/u_logic/Rdkvx4 ) );
  mux2_1 U13445 ( .ip1(n11637), .ip2(\CORTEXM0DS_INST/cm0_r14 [4]), .s(n11603), 
        .op(\CORTEXM0DS_INST/u_logic/Gikvx4 ) );
  mux2_1 U13446 ( .ip1(n11638), .ip2(\CORTEXM0DS_INST/cm0_r14 [5]), .s(n11604), 
        .op(\CORTEXM0DS_INST/u_logic/Vmkvx4 ) );
  mux2_1 U13447 ( .ip1(n11639), .ip2(\CORTEXM0DS_INST/cm0_r14 [6]), .s(n11603), 
        .op(\CORTEXM0DS_INST/u_logic/Krkvx4 ) );
  mux2_1 U13448 ( .ip1(n11640), .ip2(\CORTEXM0DS_INST/cm0_r14 [24]), .s(n11604), .op(\CORTEXM0DS_INST/u_logic/Zvkvx4 ) );
  mux2_1 U13449 ( .ip1(n11641), .ip2(\CORTEXM0DS_INST/cm0_r14 [25]), .s(n11603), .op(\CORTEXM0DS_INST/u_logic/H0lvx4 ) );
  mux2_1 U13450 ( .ip1(n11642), .ip2(\CORTEXM0DS_INST/cm0_r14 [26]), .s(n11604), .op(\CORTEXM0DS_INST/u_logic/W4lvx4 ) );
  mux2_1 U13451 ( .ip1(n11644), .ip2(\CORTEXM0DS_INST/cm0_r14 [27]), .s(n11603), .op(\CORTEXM0DS_INST/u_logic/L9lvx4 ) );
  mux2_1 U13452 ( .ip1(n11647), .ip2(\CORTEXM0DS_INST/cm0_r14 [29]), .s(n11604), .op(\CORTEXM0DS_INST/u_logic/Aelvx4 ) );
  mux2_1 U13453 ( .ip1(n11648), .ip2(\CORTEXM0DS_INST/cm0_r14 [30]), .s(n11604), .op(\CORTEXM0DS_INST/u_logic/Wilvx4 ) );
  mux2_1 U13454 ( .ip1(n11649), .ip2(\CORTEXM0DS_INST/cm0_r14 [0]), .s(n11604), 
        .op(\CORTEXM0DS_INST/u_logic/Vslvx4 ) );
  mux2_1 U13455 ( .ip1(n11650), .ip2(\CORTEXM0DS_INST/cm0_r14 [1]), .s(n11604), 
        .op(\CORTEXM0DS_INST/u_logic/Ctlvx4 ) );
  mux2_1 U13456 ( .ip1(n11651), .ip2(\CORTEXM0DS_INST/cm0_r14 [7]), .s(n11604), 
        .op(\CORTEXM0DS_INST/u_logic/Jtlvx4 ) );
  mux2_1 U13457 ( .ip1(n11652), .ip2(\CORTEXM0DS_INST/cm0_r14 [28]), .s(n11604), .op(\CORTEXM0DS_INST/u_logic/Qtlvx4 ) );
  mux2_1 U13458 ( .ip1(n11654), .ip2(\CORTEXM0DS_INST/cm0_r14 [31]), .s(n11604), .op(\CORTEXM0DS_INST/u_logic/Xtlvx4 ) );
  mux2_1 U13459 ( .ip1(n11656), .ip2(\CORTEXM0DS_INST/cm0_r12 [23]), .s(n11605), .op(\CORTEXM0DS_INST/u_logic/I7ivx4 ) );
  mux2_1 U13460 ( .ip1(n11657), .ip2(\CORTEXM0DS_INST/cm0_r12 [15]), .s(n11605), .op(\CORTEXM0DS_INST/u_logic/Xbivx4 ) );
  mux2_1 U13461 ( .ip1(n11659), .ip2(\CORTEXM0DS_INST/cm0_r12 [8]), .s(n11605), 
        .op(\CORTEXM0DS_INST/u_logic/Mgivx4 ) );
  mux2_1 U13462 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [23]), .ip2(n11656), .s(n11606), .op(\CORTEXM0DS_INST/u_logic/B7ivx4 ) );
  mux2_1 U13463 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [15]), .ip2(n11657), .s(n11606), .op(\CORTEXM0DS_INST/u_logic/Qbivx4 ) );
  mux2_1 U13464 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [8]), .ip2(n11659), .s(n11606), 
        .op(\CORTEXM0DS_INST/u_logic/Fgivx4 ) );
  inv_1 U13465 ( .ip(n11607), .op(n11620) );
  nor2_1 U13466 ( .ip1(n11608), .ip2(n11620), .op(n11609) );
  mux2_1 U13467 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [23]), .ip2(n11656), .s(n11609), .op(\CORTEXM0DS_INST/u_logic/U6ivx4 ) );
  buf_1 U13468 ( .ip(n11609), .op(n11610) );
  mux2_1 U13469 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [15]), .ip2(n11657), .s(n11610), .op(\CORTEXM0DS_INST/u_logic/Jbivx4 ) );
  mux2_1 U13470 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [8]), .ip2(n11659), .s(n11609), 
        .op(\CORTEXM0DS_INST/u_logic/Yfivx4 ) );
  mux2_1 U13471 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [9]), .ip2(n11622), .s(n11610), 
        .op(\CORTEXM0DS_INST/u_logic/Nkivx4 ) );
  mux2_1 U13472 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [2]), .ip2(n11623), .s(n11609), 
        .op(\CORTEXM0DS_INST/u_logic/Cpivx4 ) );
  mux2_1 U13473 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [10]), .ip2(n11624), .s(n11610), .op(\CORTEXM0DS_INST/u_logic/Rtivx4 ) );
  mux2_1 U13474 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [11]), .ip2(n11625), .s(n11609), .op(\CORTEXM0DS_INST/u_logic/Gyivx4 ) );
  mux2_1 U13475 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [12]), .ip2(n11626), .s(n11610), .op(\CORTEXM0DS_INST/u_logic/V2jvx4 ) );
  mux2_1 U13476 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [13]), .ip2(n11627), .s(n11609), .op(\CORTEXM0DS_INST/u_logic/K7jvx4 ) );
  mux2_1 U13477 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [14]), .ip2(n11628), .s(n11610), .op(\CORTEXM0DS_INST/u_logic/Zbjvx4 ) );
  mux2_1 U13478 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [16]), .ip2(n11629), .s(n11609), .op(\CORTEXM0DS_INST/u_logic/Ogjvx4 ) );
  mux2_1 U13479 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [17]), .ip2(n11630), .s(n11610), .op(\CORTEXM0DS_INST/u_logic/Dljvx4 ) );
  mux2_1 U13480 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [18]), .ip2(n11631), .s(n11609), .op(\CORTEXM0DS_INST/u_logic/Spjvx4 ) );
  mux2_1 U13481 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [19]), .ip2(n11632), .s(n11609), .op(\CORTEXM0DS_INST/u_logic/Hujvx4 ) );
  mux2_1 U13482 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [20]), .ip2(n11633), .s(n11609), .op(\CORTEXM0DS_INST/u_logic/Wyjvx4 ) );
  mux2_1 U13483 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [21]), .ip2(n11634), .s(n11609), .op(\CORTEXM0DS_INST/u_logic/L3kvx4 ) );
  mux2_1 U13484 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [22]), .ip2(n11635), .s(n11609), .op(\CORTEXM0DS_INST/u_logic/A8kvx4 ) );
  mux2_1 U13485 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [3]), .ip2(n11636), .s(n11609), 
        .op(\CORTEXM0DS_INST/u_logic/Wckvx4 ) );
  mux2_1 U13486 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [4]), .ip2(n11637), .s(n11609), 
        .op(\CORTEXM0DS_INST/u_logic/Lhkvx4 ) );
  mux2_1 U13487 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [5]), .ip2(n11638), .s(n11610), 
        .op(\CORTEXM0DS_INST/u_logic/Amkvx4 ) );
  mux2_1 U13488 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [6]), .ip2(n11639), .s(n11609), 
        .op(\CORTEXM0DS_INST/u_logic/Pqkvx4 ) );
  mux2_1 U13489 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [24]), .ip2(n11640), .s(n11610), .op(\CORTEXM0DS_INST/u_logic/Evkvx4 ) );
  mux2_1 U13490 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [25]), .ip2(n11641), .s(n11609), .op(\CORTEXM0DS_INST/u_logic/Mzkvx4 ) );
  mux2_1 U13491 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [26]), .ip2(n11642), .s(n11610), .op(\CORTEXM0DS_INST/u_logic/B4lvx4 ) );
  mux2_1 U13492 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [27]), .ip2(n11644), .s(n11609), .op(\CORTEXM0DS_INST/u_logic/Q8lvx4 ) );
  mux2_1 U13493 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [29]), .ip2(n11647), .s(n11610), .op(\CORTEXM0DS_INST/u_logic/Fdlvx4 ) );
  mux2_1 U13494 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [30]), .ip2(n11648), .s(n11610), .op(\CORTEXM0DS_INST/u_logic/Bilvx4 ) );
  mux2_1 U13495 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [0]), .ip2(n11649), .s(n11610), 
        .op(\CORTEXM0DS_INST/u_logic/Uolvx4 ) );
  mux2_1 U13496 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [1]), .ip2(n11650), .s(n11610), 
        .op(\CORTEXM0DS_INST/u_logic/Bplvx4 ) );
  mux2_1 U13497 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [7]), .ip2(n11651), .s(n11610), 
        .op(\CORTEXM0DS_INST/u_logic/Iplvx4 ) );
  mux2_1 U13498 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [28]), .ip2(n11652), .s(n11610), .op(\CORTEXM0DS_INST/u_logic/Pplvx4 ) );
  mux2_1 U13499 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [31]), .ip2(n11654), .s(n11610), .op(\CORTEXM0DS_INST/u_logic/Wplvx4 ) );
  mux2_1 U13500 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [23]), .ip2(n11656), .s(n11611), .op(\CORTEXM0DS_INST/u_logic/N6ivx4 ) );
  mux2_1 U13501 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [15]), .ip2(n11657), .s(n11611), .op(\CORTEXM0DS_INST/u_logic/Cbivx4 ) );
  mux2_1 U13502 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [8]), .ip2(n11659), .s(n11611), 
        .op(\CORTEXM0DS_INST/u_logic/Rfivx4 ) );
  mux2_1 U13503 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [23]), .ip2(n11656), .s(n11612), .op(\CORTEXM0DS_INST/u_logic/G6ivx4 ) );
  mux2_1 U13504 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [15]), .ip2(n11657), .s(n11612), .op(\CORTEXM0DS_INST/u_logic/Vaivx4 ) );
  mux2_1 U13505 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [8]), .ip2(n11659), .s(n11612), 
        .op(\CORTEXM0DS_INST/u_logic/Kfivx4 ) );
  mux2_1 U13506 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [23]), .ip2(n11656), .s(n11613), .op(\CORTEXM0DS_INST/u_logic/Z5ivx4 ) );
  mux2_1 U13507 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [15]), .ip2(n11657), .s(n11613), .op(\CORTEXM0DS_INST/u_logic/Oaivx4 ) );
  mux2_1 U13508 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [8]), .ip2(n11659), .s(n11613), 
        .op(\CORTEXM0DS_INST/u_logic/Dfivx4 ) );
  nor2_1 U13509 ( .ip1(n11614), .ip2(n11620), .op(n11615) );
  mux2_1 U13510 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [23]), .ip2(n11656), .s(n11615), .op(\CORTEXM0DS_INST/u_logic/S5ivx4 ) );
  buf_1 U13511 ( .ip(n11615), .op(n11616) );
  mux2_1 U13512 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [15]), .ip2(n11657), .s(n11616), .op(\CORTEXM0DS_INST/u_logic/Haivx4 ) );
  mux2_1 U13513 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [8]), .ip2(n11659), .s(n11615), 
        .op(\CORTEXM0DS_INST/u_logic/Weivx4 ) );
  mux2_1 U13514 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [9]), .ip2(n11622), .s(n11616), 
        .op(\CORTEXM0DS_INST/u_logic/Ljivx4 ) );
  mux2_1 U13515 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [2]), .ip2(n11623), .s(n11615), 
        .op(\CORTEXM0DS_INST/u_logic/Aoivx4 ) );
  mux2_1 U13516 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [10]), .ip2(n11624), .s(n11616), .op(\CORTEXM0DS_INST/u_logic/Psivx4 ) );
  mux2_1 U13517 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [11]), .ip2(n11625), .s(n11615), .op(\CORTEXM0DS_INST/u_logic/Exivx4 ) );
  mux2_1 U13518 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [12]), .ip2(n11626), .s(n11616), .op(\CORTEXM0DS_INST/u_logic/T1jvx4 ) );
  mux2_1 U13519 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [13]), .ip2(n11627), .s(n11615), .op(\CORTEXM0DS_INST/u_logic/I6jvx4 ) );
  mux2_1 U13520 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [14]), .ip2(n11628), .s(n11616), .op(\CORTEXM0DS_INST/u_logic/Xajvx4 ) );
  mux2_1 U13521 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [16]), .ip2(n11629), .s(n11615), .op(\CORTEXM0DS_INST/u_logic/Mfjvx4 ) );
  mux2_1 U13522 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [17]), .ip2(n11630), .s(n11616), .op(\CORTEXM0DS_INST/u_logic/Bkjvx4 ) );
  mux2_1 U13523 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [18]), .ip2(n11631), .s(n11615), .op(\CORTEXM0DS_INST/u_logic/Qojvx4 ) );
  mux2_1 U13524 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [19]), .ip2(n11632), .s(n11615), .op(\CORTEXM0DS_INST/u_logic/Ftjvx4 ) );
  mux2_1 U13525 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [20]), .ip2(n11633), .s(n11615), .op(\CORTEXM0DS_INST/u_logic/Uxjvx4 ) );
  mux2_1 U13526 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [21]), .ip2(n11634), .s(n11615), .op(\CORTEXM0DS_INST/u_logic/J2kvx4 ) );
  mux2_1 U13527 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [22]), .ip2(n11635), .s(n11615), .op(\CORTEXM0DS_INST/u_logic/Y6kvx4 ) );
  mux2_1 U13528 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [3]), .ip2(n11636), .s(n11615), 
        .op(\CORTEXM0DS_INST/u_logic/Ubkvx4 ) );
  mux2_1 U13529 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [4]), .ip2(n11637), .s(n11615), 
        .op(\CORTEXM0DS_INST/u_logic/Jgkvx4 ) );
  mux2_1 U13530 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [5]), .ip2(n11638), .s(n11616), 
        .op(\CORTEXM0DS_INST/u_logic/Ykkvx4 ) );
  mux2_1 U13531 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [6]), .ip2(n11639), .s(n11615), 
        .op(\CORTEXM0DS_INST/u_logic/Npkvx4 ) );
  mux2_1 U13532 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [24]), .ip2(n11640), .s(n11616), .op(\CORTEXM0DS_INST/u_logic/Cukvx4 ) );
  mux2_1 U13533 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [25]), .ip2(n11641), .s(n11615), .op(\CORTEXM0DS_INST/u_logic/Kykvx4 ) );
  mux2_1 U13534 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [26]), .ip2(n11642), .s(n11616), .op(\CORTEXM0DS_INST/u_logic/Z2lvx4 ) );
  mux2_1 U13535 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [27]), .ip2(n11644), .s(n11615), .op(\CORTEXM0DS_INST/u_logic/O7lvx4 ) );
  mux2_1 U13536 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [29]), .ip2(n11647), .s(n11616), .op(\CORTEXM0DS_INST/u_logic/Dclvx4 ) );
  mux2_1 U13537 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [30]), .ip2(n11648), .s(n11616), .op(\CORTEXM0DS_INST/u_logic/Zglvx4 ) );
  mux2_1 U13538 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [0]), .ip2(n11649), .s(n11616), 
        .op(\CORTEXM0DS_INST/u_logic/Nvlvx4 ) );
  mux2_1 U13539 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [1]), .ip2(n11650), .s(n11616), 
        .op(\CORTEXM0DS_INST/u_logic/Uvlvx4 ) );
  mux2_1 U13540 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [7]), .ip2(n11651), .s(n11616), 
        .op(\CORTEXM0DS_INST/u_logic/Bwlvx4 ) );
  mux2_1 U13541 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [28]), .ip2(n11652), .s(n11616), .op(\CORTEXM0DS_INST/u_logic/Iwlvx4 ) );
  mux2_1 U13542 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [31]), .ip2(n11654), .s(n11616), .op(\CORTEXM0DS_INST/u_logic/Pwlvx4 ) );
  mux2_1 U13543 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [23]), .ip2(n11656), .s(n11617), .op(\CORTEXM0DS_INST/u_logic/L5ivx4 ) );
  mux2_1 U13544 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [15]), .ip2(n11657), .s(n11617), .op(\CORTEXM0DS_INST/u_logic/Aaivx4 ) );
  mux2_1 U13545 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [8]), .ip2(n11659), .s(n11617), 
        .op(\CORTEXM0DS_INST/u_logic/Peivx4 ) );
  mux2_1 U13546 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [23]), .ip2(n11656), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/E5ivx4 ) );
  mux2_1 U13547 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [15]), .ip2(n11657), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/T9ivx4 ) );
  mux2_1 U13548 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [8]), .ip2(n11659), .s(n11618), 
        .op(\CORTEXM0DS_INST/u_logic/Ieivx4 ) );
  mux2_1 U13549 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [23]), .ip2(n11656), .s(n11619), .op(\CORTEXM0DS_INST/u_logic/X4ivx4 ) );
  mux2_1 U13550 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [15]), .ip2(n11657), .s(n11619), .op(\CORTEXM0DS_INST/u_logic/M9ivx4 ) );
  mux2_1 U13551 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [8]), .ip2(n11659), .s(n11619), 
        .op(\CORTEXM0DS_INST/u_logic/Beivx4 ) );
  nor2_1 U13552 ( .ip1(n11621), .ip2(n11620), .op(n11643) );
  mux2_1 U13553 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [23]), .ip2(n11656), .s(n11643), .op(\CORTEXM0DS_INST/u_logic/Q4ivx4 ) );
  buf_1 U13554 ( .ip(n11643), .op(n11653) );
  mux2_1 U13555 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [15]), .ip2(n11657), .s(n11653), .op(\CORTEXM0DS_INST/u_logic/F9ivx4 ) );
  mux2_1 U13556 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [8]), .ip2(n11659), .s(n11643), 
        .op(\CORTEXM0DS_INST/u_logic/Udivx4 ) );
  mux2_1 U13557 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [9]), .ip2(n11622), .s(n11653), 
        .op(\CORTEXM0DS_INST/u_logic/Jiivx4 ) );
  mux2_1 U13558 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [2]), .ip2(n11623), .s(n11643), 
        .op(\CORTEXM0DS_INST/u_logic/Ymivx4 ) );
  mux2_1 U13559 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [10]), .ip2(n11624), .s(n11653), .op(\CORTEXM0DS_INST/u_logic/Nrivx4 ) );
  mux2_1 U13560 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [11]), .ip2(n11625), .s(n11643), .op(\CORTEXM0DS_INST/u_logic/Cwivx4 ) );
  mux2_1 U13561 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [12]), .ip2(n11626), .s(n11653), .op(\CORTEXM0DS_INST/u_logic/R0jvx4 ) );
  mux2_1 U13562 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [13]), .ip2(n11627), .s(n11643), .op(\CORTEXM0DS_INST/u_logic/G5jvx4 ) );
  mux2_1 U13563 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [14]), .ip2(n11628), .s(n11653), .op(\CORTEXM0DS_INST/u_logic/V9jvx4 ) );
  mux2_1 U13564 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [16]), .ip2(n11629), .s(n11643), .op(\CORTEXM0DS_INST/u_logic/Kejvx4 ) );
  mux2_1 U13565 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [17]), .ip2(n11630), .s(n11653), .op(\CORTEXM0DS_INST/u_logic/Zijvx4 ) );
  mux2_1 U13566 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [18]), .ip2(n11631), .s(n11643), .op(\CORTEXM0DS_INST/u_logic/Onjvx4 ) );
  mux2_1 U13567 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [19]), .ip2(n11632), .s(n11643), .op(\CORTEXM0DS_INST/u_logic/Dsjvx4 ) );
  mux2_1 U13568 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [20]), .ip2(n11633), .s(n11643), .op(\CORTEXM0DS_INST/u_logic/Swjvx4 ) );
  mux2_1 U13569 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [21]), .ip2(n11634), .s(n11643), .op(\CORTEXM0DS_INST/u_logic/H1kvx4 ) );
  mux2_1 U13570 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [22]), .ip2(n11635), .s(n11643), .op(\CORTEXM0DS_INST/u_logic/W5kvx4 ) );
  mux2_1 U13571 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [3]), .ip2(n11636), .s(n11643), 
        .op(\CORTEXM0DS_INST/u_logic/Sakvx4 ) );
  mux2_1 U13572 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [4]), .ip2(n11637), .s(n11643), 
        .op(\CORTEXM0DS_INST/u_logic/Hfkvx4 ) );
  mux2_1 U13573 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [5]), .ip2(n11638), .s(n11653), 
        .op(\CORTEXM0DS_INST/u_logic/Wjkvx4 ) );
  mux2_1 U13574 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [6]), .ip2(n11639), .s(n11643), 
        .op(\CORTEXM0DS_INST/u_logic/Lokvx4 ) );
  mux2_1 U13575 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [24]), .ip2(n11640), .s(n11653), .op(\CORTEXM0DS_INST/u_logic/Atkvx4 ) );
  mux2_1 U13576 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [25]), .ip2(n11641), .s(n11643), .op(\CORTEXM0DS_INST/u_logic/Ixkvx4 ) );
  mux2_1 U13577 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [26]), .ip2(n11642), .s(n11653), .op(\CORTEXM0DS_INST/u_logic/X1lvx4 ) );
  mux2_1 U13578 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [27]), .ip2(n11644), .s(n11643), .op(\CORTEXM0DS_INST/u_logic/M6lvx4 ) );
  and2_1 U13579 ( .ip1(n11646), .ip2(n11645), .op(n4180) );
  mux2_1 U13580 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [29]), .ip2(n11647), .s(n11653), .op(\CORTEXM0DS_INST/u_logic/Bblvx4 ) );
  mux2_1 U13581 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [30]), .ip2(n11648), .s(n11653), .op(\CORTEXM0DS_INST/u_logic/Xflvx4 ) );
  mux2_1 U13582 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [0]), .ip2(n11649), .s(n11653), 
        .op(\CORTEXM0DS_INST/u_logic/X0mvx4 ) );
  mux2_1 U13583 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [1]), .ip2(n11650), .s(n11653), 
        .op(\CORTEXM0DS_INST/u_logic/E1mvx4 ) );
  mux2_1 U13584 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [7]), .ip2(n11651), .s(n11653), 
        .op(\CORTEXM0DS_INST/u_logic/L1mvx4 ) );
  mux2_1 U13585 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [28]), .ip2(n11652), .s(n11653), .op(\CORTEXM0DS_INST/u_logic/S1mvx4 ) );
  mux2_1 U13586 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [31]), .ip2(n11654), .s(n11653), .op(\CORTEXM0DS_INST/u_logic/Z1mvx4 ) );
  mux2_1 U13587 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [23]), .ip2(n11656), .s(n11655), .op(\CORTEXM0DS_INST/u_logic/J4ivx4 ) );
  mux2_1 U13588 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [15]), .ip2(n11657), .s(n11655), .op(\CORTEXM0DS_INST/u_logic/Y8ivx4 ) );
  mux2_1 U13589 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [8]), .ip2(n11659), .s(n11655), 
        .op(\CORTEXM0DS_INST/u_logic/Ndivx4 ) );
  mux2_1 U13590 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [23]), .ip2(n11656), .s(n11658), .op(\CORTEXM0DS_INST/u_logic/C4ivx4 ) );
  mux2_1 U13591 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [15]), .ip2(n11657), .s(n11658), .op(\CORTEXM0DS_INST/u_logic/R8ivx4 ) );
  mux2_1 U13592 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [8]), .ip2(n11659), .s(n11658), 
        .op(\CORTEXM0DS_INST/u_logic/Gdivx4 ) );
  nor2_1 U13593 ( .ip1(n11661), .ip2(n11660), .op(n3959) );
  nor2_1 U13594 ( .ip1(n11662), .ip2(n11820), .op(n11666) );
  nor2_1 U13595 ( .ip1(n11664), .ip2(n11663), .op(n11665) );
  ab_or_c_or_d U13596 ( .ip1(n11668), .ip2(n11667), .ip3(n11666), .ip4(n11665), 
        .op(n11670) );
  not_ab_or_c_or_d U13597 ( .ip1(n11669), .ip2(n11825), .ip3(1'b0), .ip4(n5932), .op(n11676) );
  mux2_1 U13598 ( .ip1(\CORTEXM0DS_INST/vis_apsr [3]), .ip2(n11670), .s(n11676), .op(\CORTEXM0DS_INST/u_logic/V3ivx4 ) );
  nor2_1 U13599 ( .ip1(n11671), .ip2(n11818), .op(n11674) );
  nor2_1 U13600 ( .ip1(n11672), .ip2(n11820), .op(n11673) );
  ab_or_c_or_d U13601 ( .ip1(n11825), .ip2(n11675), .ip3(n11674), .ip4(n11673), 
        .op(n11677) );
  mux2_1 U13602 ( .ip1(\CORTEXM0DS_INST/vis_apsr [2]), .ip2(n11677), .s(n11676), .op(\CORTEXM0DS_INST/u_logic/Cflvx4 ) );
  and3_1 U13603 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n11679), .ip3(
        n11678), .op(TXEV_top_out) );
  nor4_1 U13604 ( .ip1(n11683), .ip2(n11682), .ip3(n11681), .ip4(n11680), .op(
        n11704) );
  nor2_1 U13605 ( .ip1(n11684), .ip2(n11704), .op(n11685) );
  nor2_1 U13606 ( .ip1(n11703), .ip2(n11685), .op(n11889) );
  nand2_1 U13607 ( .ip1(n11889), .ip2(n11885), .op(n11749) );
  nor2_1 U13608 ( .ip1(n11687), .ip2(n11686), .op(n12409) );
  nand2_1 U13609 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Dmgvx4 ), .op(n12412) );
  not_ab_or_c_or_d U13610 ( .ip1(n12409), .ip2(n12652), .ip3(
        \CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip4(n12412), .op(n11702) );
  or2_1 U13611 ( .ip1(n11688), .ip2(\CORTEXM0DS_INST/u_logic/Rkgvx4 ), .op(
        n11700) );
  nor2_1 U13612 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n11689), .op(
        n11696) );
  nor3_1 U13613 ( .ip1(n12118), .ip2(n5639), .ip3(n12413), .op(n11695) );
  nor4_1 U13614 ( .ip1(n11693), .ip2(n11692), .ip3(n11691), .ip4(n11690), .op(
        n11694) );
  not_ab_or_c_or_d U13615 ( .ip1(n11697), .ip2(n11696), .ip3(n11695), .ip4(
        n11694), .op(n11698) );
  or2_1 U13616 ( .ip1(n11698), .ip2(\CORTEXM0DS_INST/u_logic/Rkgvx4 ), .op(
        n11699) );
  nand2_1 U13617 ( .ip1(n11700), .ip2(n11699), .op(n11701) );
  not_ab_or_c_or_d U13618 ( .ip1(n11704), .ip2(n11703), .ip3(n11702), .ip4(
        n11701), .op(n11883) );
  nor2_1 U13619 ( .ip1(\CORTEXM0DS_INST/u_logic/Krgvx4 ), .ip2(n11883), .op(
        n11736) );
  nor2_1 U13620 ( .ip1(n3233), .ip2(n11705), .op(n11725) );
  inv_1 U13621 ( .ip(\CORTEXM0DS_INST/u_logic/P0ivx4 ), .op(n11706) );
  nor2_1 U13622 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [8]), .ip2(n11706), 
        .op(n11715) );
  nand2_1 U13623 ( .ip1(\CORTEXM0DS_INST/u_logic/Nzhvx4 ), .ip2(n11707), .op(
        n11713) );
  nand2_1 U13624 ( .ip1(\CORTEXM0DS_INST/u_logic/Y1ivx4 ), .ip2(n11708), .op(
        n11712) );
  nand2_1 U13625 ( .ip1(\CORTEXM0DS_INST/u_logic/D1ivx4 ), .ip2(n11709), .op(
        n11711) );
  inv_1 U13626 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [15]), .op(n11831) );
  nand2_1 U13627 ( .ip1(\CORTEXM0DS_INST/u_logic/Syhvx4 ), .ip2(n11831), .op(
        n11710) );
  nand4_1 U13628 ( .ip1(n11713), .ip2(n11712), .ip3(n11711), .ip4(n11710), 
        .op(n11714) );
  not_ab_or_c_or_d U13629 ( .ip1(\CORTEXM0DS_INST/u_logic/T2ivx4 ), .ip2(
        n11716), .ip3(n11715), .ip4(n11714), .op(n11723) );
  inv_1 U13630 ( .ip(\CORTEXM0DS_INST/u_logic/Eqgvx4 ), .op(n11717) );
  nand2_1 U13631 ( .ip1(\CORTEXM0DS_INST/u_logic/Owgvx4 ), .ip2(n11717), .op(
        n11722) );
  nand2_1 U13632 ( .ip1(\CORTEXM0DS_INST/u_logic/Gzhvx4 ), .ip2(n11718), .op(
        n11721) );
  inv_1 U13633 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [10]), .op(n11719) );
  nand2_1 U13634 ( .ip1(\CORTEXM0DS_INST/u_logic/B0ivx4 ), .ip2(n11719), .op(
        n11720) );
  nand4_1 U13635 ( .ip1(n11723), .ip2(n11722), .ip3(n11721), .ip4(n11720), 
        .op(n11724) );
  not_ab_or_c_or_d U13636 ( .ip1(\CORTEXM0DS_INST/u_logic/Zyhvx4 ), .ip2(
        n11726), .ip3(n11725), .ip4(n11724), .op(n11734) );
  nand2_1 U13637 ( .ip1(\CORTEXM0DS_INST/u_logic/Uzhvx4 ), .ip2(n11727), .op(
        n11733) );
  inv_1 U13638 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [9]), .op(n11728) );
  nand2_1 U13639 ( .ip1(\CORTEXM0DS_INST/u_logic/I0ivx4 ), .ip2(n11728), .op(
        n11732) );
  nor2_1 U13640 ( .ip1(n2326), .ip2(n3224), .op(n11729) );
  nor2_1 U13641 ( .ip1(n12747), .ip2(n11729), .op(n12048) );
  nand2_1 U13642 ( .ip1(n12048), .ip2(n11730), .op(n11731) );
  nand4_1 U13643 ( .ip1(n11734), .ip2(n11733), .ip3(n11732), .ip4(n11731), 
        .op(n11735) );
  not_ab_or_c_or_d U13644 ( .ip1(\CORTEXM0DS_INST/u_logic/W0ivx4 ), .ip2(n3223), .ip3(n11736), .ip4(n11735), .op(n11748) );
  inv_1 U13645 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [1]), .op(n11746) );
  inv_1 U13646 ( .ip(n3224), .op(n11737) );
  nor3_1 U13647 ( .ip1(\CORTEXM0DS_INST/u_logic/Qsgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Sx3wx4 ), .ip3(n11737), .op(n11745) );
  inv_1 U13648 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [2]), .op(n11738) );
  nand2_1 U13649 ( .ip1(n11738), .ip2(\CORTEXM0DS_INST/u_logic/F2ivx4 ), .op(
        n11743) );
  nand2_1 U13650 ( .ip1(\CORTEXM0DS_INST/u_logic/K1ivx4 ), .ip2(n11739), .op(
        n11742) );
  nand2_1 U13651 ( .ip1(\CORTEXM0DS_INST/u_logic/R1ivx4 ), .ip2(n11740), .op(
        n11741) );
  nand3_1 U13652 ( .ip1(n11743), .ip2(n11742), .ip3(n11741), .op(n11744) );
  not_ab_or_c_or_d U13653 ( .ip1(\CORTEXM0DS_INST/u_logic/M2ivx4 ), .ip2(
        n11746), .ip3(n11745), .ip4(n11744), .op(n11747) );
  nand3_1 U13654 ( .ip1(n11749), .ip2(n11748), .ip3(n11747), .op(n11750) );
  nand2_1 U13655 ( .ip1(\CORTEXM0DS_INST/u_logic/Vogvx4 ), .ip2(n11750), .op(
        n11753) );
  not_ab_or_c_or_d U13656 ( .ip1(n11751), .ip2(n12623), .ip3(TXEV_top_out), 
        .ip4(n3276), .op(n11752) );
  nand2_1 U13657 ( .ip1(n11753), .ip2(n11752), .op(n11759) );
  or4_1 U13658 ( .ip1(n11757), .ip2(n11756), .ip3(n11755), .ip4(n11754), .op(
        n11758) );
  mux2_1 U13659 ( .ip1(n11759), .ip2(n11758), .s(
        \CORTEXM0DS_INST/u_logic/Ih8vx4 ), .op(
        \CORTEXM0DS_INST/u_logic/H3ivx4 ) );
  inv_1 U13660 ( .ip(n12409), .op(n3217) );
  inv_1 U13661 ( .ip(n11760), .op(n11762) );
  mux2_1 U13662 ( .ip1(n11762), .ip2(n11761), .s(n3217), .op(n11767) );
  not_ab_or_c_or_d U13663 ( .ip1(n11765), .ip2(n11764), .ip3(n5932), .ip4(
        n11763), .op(n11766) );
  mux2_1 U13664 ( .ip1(\CORTEXM0DS_INST/u_logic/Oy8vx4 ), .ip2(n11767), .s(
        n11766), .op(\CORTEXM0DS_INST/u_logic/Sqivx4 ) );
  nand3_1 U13665 ( .ip1(\CORTEXM0DS_INST/u_logic/B19vx4 ), .ip2(n11768), .ip3(
        n11796), .op(n11785) );
  or2_1 U13666 ( .ip1(n12138), .ip2(\CORTEXM0DS_INST/cm0_control[1] ), .op(
        n11770) );
  or2_1 U13667 ( .ip1(\CORTEXM0DS_INST/vis_pc [1]), .ip2(
        \CORTEXM0DS_INST/cm0_control[1] ), .op(n11769) );
  nand2_1 U13668 ( .ip1(n11770), .ip2(n11769), .op(n11781) );
  nor2_1 U13669 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n11789), .op(
        n11778) );
  or2_1 U13670 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n8424), .op(
        n11772) );
  or2_1 U13671 ( .ip1(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), .ip2(n8424), .op(
        n11771) );
  nand2_1 U13672 ( .ip1(n11772), .ip2(n11771), .op(n11777) );
  or2_1 U13673 ( .ip1(\CORTEXM0DS_INST/u_logic/P39vx4 ), .ip2(n11773), .op(
        n11775) );
  or2_1 U13674 ( .ip1(n11796), .ip2(n11773), .op(n11774) );
  nand2_1 U13675 ( .ip1(n11775), .ip2(n11774), .op(n11776) );
  nor4_1 U13676 ( .ip1(n11779), .ip2(n11778), .ip3(n11777), .ip4(n11776), .op(
        n11780) );
  or2_1 U13677 ( .ip1(n11781), .ip2(n11780), .op(n11784) );
  nand3_1 U13678 ( .ip1(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), .ip2(n11782), .ip3(
        n8424), .op(n11783) );
  nand3_1 U13679 ( .ip1(n11785), .ip2(n11784), .ip3(n11783), .op(n11806) );
  nand2_1 U13680 ( .ip1(n11787), .ip2(n11786), .op(n11800) );
  nor3_1 U13681 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n11789), .ip3(
        n11788), .op(n11790) );
  not_ab_or_c_or_d U13682 ( .ip1(n11792), .ip2(n12134), .ip3(n11791), .ip4(
        n11790), .op(n11799) );
  nor2_1 U13683 ( .ip1(n11793), .ip2(n12070), .op(n11795) );
  not_ab_or_c_or_d U13684 ( .ip1(n11797), .ip2(n11796), .ip3(n11795), .ip4(
        n11794), .op(n11798) );
  nand3_1 U13685 ( .ip1(n11800), .ip2(n11799), .ip3(n11798), .op(n11801) );
  not_ab_or_c_or_d U13686 ( .ip1(n11803), .ip2(
        \CORTEXM0DS_INST/u_logic/P39vx4 ), .ip3(n11802), .ip4(n11801), .op(
        n11804) );
  nor2_1 U13687 ( .ip1(n5932), .ip2(n11804), .op(n11805) );
  mux2_1 U13688 ( .ip1(\CORTEXM0DS_INST/u_logic/O7evx4 ), .ip2(n11806), .s(
        n11805), .op(\CORTEXM0DS_INST/u_logic/Hllvx4 ) );
  nand2_1 U13689 ( .ip1(\CORTEXM0DS_INST/vis_pc [1]), .ip2(
        \CORTEXM0DS_INST/u_logic/Hx8vx4 ), .op(n11809) );
  or2_1 U13690 ( .ip1(n11812), .ip2(n11807), .op(n11808) );
  nand2_1 U13691 ( .ip1(n11809), .ip2(n11808), .op(n11816) );
  nor3_1 U13692 ( .ip1(n11812), .ip2(n11811), .ip3(n11810), .op(n11813) );
  nor3_1 U13693 ( .ip1(n11813), .ip2(n12138), .ip3(n3276), .op(n11814) );
  nor2_1 U13694 ( .ip1(n5932), .ip2(n11814), .op(n11815) );
  mux2_1 U13695 ( .ip1(\CORTEXM0DS_INST/cm0_control[1] ), .ip2(n11816), .s(
        n11815), .op(\CORTEXM0DS_INST/u_logic/Ollvx4 ) );
  nor2_1 U13696 ( .ip1(n12687), .ip2(n11817), .op(n3129) );
  nor2_1 U13697 ( .ip1(n11819), .ip2(n11818), .op(n11823) );
  nor2_1 U13698 ( .ip1(n11821), .ip2(n11820), .op(n11822) );
  ab_or_c_or_d U13699 ( .ip1(n11825), .ip2(n11824), .ip3(n11823), .ip4(n11822), 
        .op(n11828) );
  not_ab_or_c_or_d U13700 ( .ip1(n11826), .ip2(n11825), .ip3(1'b0), .ip4(n5932), .op(n11827) );
  mux2_1 U13701 ( .ip1(\CORTEXM0DS_INST/vis_apsr [1]), .ip2(n11828), .s(n11827), .op(\CORTEXM0DS_INST/u_logic/Finvx4 ) );
  nor2_1 U13702 ( .ip1(n11875), .ip2(n11937), .op(n3082) );
  and2_1 U13703 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [5]), .ip2(n11829), 
        .op(n3083) );
  nor2_1 U13704 ( .ip1(n11831), .ip2(n11830), .op(n3030) );
  and2_1 U13705 ( .ip1(n11832), .ip2(n11853), .op(n3017) );
  inv_1 U13706 ( .ip(n11841), .op(n11859) );
  nor2_1 U13707 ( .ip1(n11859), .ip2(n11833), .op(n11838) );
  nand2_1 U13708 ( .ip1(n11864), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [13]), 
        .op(n11836) );
  nand2_1 U13709 ( .ip1(\CORTEXM0DS_INST/u_logic/Psh2z4 [1]), .ip2(n12643), 
        .op(n11835) );
  nand2_1 U13710 ( .ip1(n11842), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [29]), 
        .op(n11834) );
  nand3_1 U13711 ( .ip1(n11836), .ip2(n11835), .ip3(n11834), .op(n11837) );
  not_ab_or_c_or_d U13712 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [21]), .ip2(
        n11863), .ip3(n11838), .ip4(n11837), .op(n11839) );
  nor2_1 U13713 ( .ip1(n11839), .ip2(n11871), .op(n3018) );
  and2_1 U13714 ( .ip1(n11840), .ip2(n11853), .op(n3008) );
  and2_1 U13715 ( .ip1(n11841), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [7]), 
        .op(n11850) );
  nand2_1 U13716 ( .ip1(\CORTEXM0DS_INST/u_logic/Uth2z4 [1]), .ip2(n12642), 
        .op(n11846) );
  nand2_1 U13717 ( .ip1(n11864), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [15]), 
        .op(n11845) );
  nand2_1 U13718 ( .ip1(n11842), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [31]), 
        .op(n11844) );
  nand2_1 U13719 ( .ip1(\CORTEXM0DS_INST/u_logic/Txh2z4 [1]), .ip2(n12643), 
        .op(n11843) );
  nand4_1 U13720 ( .ip1(n11846), .ip2(n11845), .ip3(n11844), .ip4(n11843), 
        .op(n11847) );
  ab_or_c_or_d U13721 ( .ip1(n11863), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [23]), .ip3(n11848), .ip4(n11847), 
        .op(n11849) );
  not_ab_or_c_or_d U13722 ( .ip1(n11851), .ip2(
        \CORTEXM0DS_INST/u_logic/Eqgvx4 ), .ip3(n11850), .ip4(n11849), .op(
        n11852) );
  nor2_1 U13723 ( .ip1(n11852), .ip2(n11871), .op(n3009) );
  nand2_1 U13724 ( .ip1(n11854), .ip2(n11853), .op(n11874) );
  nor2_1 U13725 ( .ip1(n11856), .ip2(n11855), .op(n11869) );
  nand2_1 U13726 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [7]), .ip2(n11857), 
        .op(n11867) );
  nor2_1 U13727 ( .ip1(n11859), .ip2(n11858), .op(n11862) );
  nor2_1 U13728 ( .ip1(n3223), .ip2(n11860), .op(n11861) );
  not_ab_or_c_or_d U13729 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [17]), .ip2(
        n11863), .ip3(n11862), .ip4(n11861), .op(n11866) );
  nand2_1 U13730 ( .ip1(n11864), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [9]), 
        .op(n11865) );
  nand3_1 U13731 ( .ip1(n11867), .ip2(n11866), .ip3(n11865), .op(n11868) );
  not_ab_or_c_or_d U13732 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [7]), .ip2(
        n11870), .ip3(n11869), .ip4(n11868), .op(n11872) );
  or2_1 U13733 ( .ip1(n11872), .ip2(n11871), .op(n11873) );
  nand2_1 U13734 ( .ip1(n11874), .ip2(n11873), .op(n2994) );
  inv_1 U13735 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [7]), .op(n11949) );
  nor2_1 U13736 ( .ip1(n11875), .ip2(n11949), .op(n2995) );
  nor2_1 U13737 ( .ip1(n11876), .ip2(n11895), .op(n2791) );
  mux2_1 U13738 ( .ip1(n11898), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [0]), .s(
        n2786), .op(n6186) );
  mux2_1 U13739 ( .ip1(n11898), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [1]), .s(
        n2774), .op(n6183) );
  mux2_1 U13740 ( .ip1(n11898), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [14]), 
        .s(n2757), .op(n6177) );
  nor2_1 U13741 ( .ip1(n11877), .ip2(n11895), .op(n2714) );
  mux2_1 U13742 ( .ip1(n11898), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [6]), .s(
        n2711), .op(n6176) );
  mux2_1 U13743 ( .ip1(n11898), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [5]), .s(
        n2686), .op(n6174) );
  nor2_1 U13744 ( .ip1(n11878), .ip2(n11895), .op(n2648) );
  mux2_1 U13745 ( .ip1(n11898), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [12]), 
        .s(n2645), .op(n6171) );
  mux2_1 U13746 ( .ip1(n11898), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [4]), .s(
        n2644), .op(n6169) );
  nor3_1 U13747 ( .ip1(n11880), .ip2(n11879), .ip3(n11895), .op(n2627) );
  mux2_1 U13748 ( .ip1(n11898), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [3]), .s(
        n2624), .op(n6167) );
  mux2_1 U13749 ( .ip1(n11898), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [2]), .s(
        n2623), .op(n6165) );
  mux2_1 U13750 ( .ip1(n11898), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [7]), .s(
        n2577), .op(n6160) );
  nand3_1 U13751 ( .ip1(n12402), .ip2(n3276), .ip3(n12403), .op(n11881) );
  nand2_1 U13752 ( .ip1(\CORTEXM0DS_INST/u_logic/Krgvx4 ), .ip2(n11881), .op(
        n11882) );
  nand2_1 U13753 ( .ip1(n11883), .ip2(n11882), .op(n6158) );
  or2_1 U13754 ( .ip1(n11884), .ip2(n11885), .op(n11887) );
  or2_1 U13755 ( .ip1(n3276), .ip2(n11885), .op(n11886) );
  nand2_1 U13756 ( .ip1(n11887), .ip2(n11886), .op(n11888) );
  or2_1 U13757 ( .ip1(n11889), .ip2(n11888), .op(n6157) );
  and2_1 U13758 ( .ip1(n11890), .ip2(n3276), .op(n2544) );
  mux2_1 U13759 ( .ip1(n11898), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [10]), 
        .s(n2541), .op(n6156) );
  mux2_1 U13760 ( .ip1(n11898), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [11]), 
        .s(n2533), .op(n6153) );
  mux2_1 U13761 ( .ip1(n11898), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [9]), .s(
        n2514), .op(n6151) );
  mux2_1 U13762 ( .ip1(n11898), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [8]), .s(
        n2513), .op(n6150) );
  nor2_1 U13763 ( .ip1(n11891), .ip2(n11895), .op(n2512) );
  mux2_1 U13764 ( .ip1(n11898), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [13]), 
        .s(n2500), .op(n6147) );
  nand2_1 U13765 ( .ip1(n11892), .ip2(n3276), .op(n11893) );
  nand3_1 U13766 ( .ip1(n11893), .ip2(n2490), .ip3(
        \CORTEXM0DS_INST/u_logic/Qsgvx4 ), .op(n11894) );
  nand2_1 U13767 ( .ip1(n2492), .ip2(n11894), .op(n6143) );
  nor3_1 U13768 ( .ip1(n11897), .ip2(n11896), .ip3(n11895), .op(n2464) );
  mux2_1 U13769 ( .ip1(n11898), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [15]), 
        .s(n2460), .op(n6141) );
  nor2_1 U13770 ( .ip1(n11899), .ip2(n12687), .op(n2785) );
  nand2_1 U13771 ( .ip1(\CORTEXM0DS_INST/u_logic/Z7hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/B5hvx4 ), .op(n11900) );
  nor4_1 U13772 ( .ip1(n12689), .ip2(n11901), .ip3(n11900), .ip4(n12687), .op(
        n11913) );
  inv_1 U13773 ( .ip(n11913), .op(n11907) );
  nand3_1 U13774 ( .ip1(n11903), .ip2(n11902), .ip3(n12687), .op(n11904) );
  nand3_1 U13775 ( .ip1(n11907), .ip2(\CORTEXM0DS_INST/u_logic/Izgvx4 ), .ip3(
        n11904), .op(n11906) );
  nand3_1 U13776 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [0]), .ip2(
        \CORTEXM0DS_INST/u_logic/F2hvx4 ), .ip3(n11908), .op(n11905) );
  nand2_1 U13777 ( .ip1(n11906), .ip2(n11905), .op(n6139) );
  nand2_1 U13778 ( .ip1(n11907), .ip2(\CORTEXM0DS_INST/u_logic/F2hvx4 ), .op(
        n11909) );
  inv_1 U13779 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [0]), .op(n11914) );
  nand2_1 U13780 ( .ip1(n11908), .ip2(n11914), .op(n11910) );
  nor2_1 U13781 ( .ip1(n11909), .ip2(n11910), .op(n12041) );
  inv_1 U13782 ( .ip(n11909), .op(n11929) );
  nand2_1 U13783 ( .ip1(n11929), .ip2(n11910), .op(n11974) );
  nor2_1 U13784 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [0]), .ip2(n11974), 
        .op(n11912) );
  nor3_1 U13785 ( .ip1(\CORTEXM0DS_INST/u_logic/F2hvx4 ), .ip2(n11913), .ip3(
        n11914), .op(n11911) );
  ab_or_c_or_d U13786 ( .ip1(n12041), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [0]), .ip3(n11912), .ip4(n11911), .op(n6138) );
  or2_1 U13787 ( .ip1(\CORTEXM0DS_INST/u_logic/F2hvx4 ), .ip2(n11913), .op(
        n11916) );
  or2_1 U13788 ( .ip1(n11914), .ip2(n11913), .op(n11915) );
  nand2_1 U13789 ( .ip1(n11916), .ip2(n11915), .op(n11924) );
  nor3_1 U13790 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [0]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [1]), .ip3(n11974), .op(n11918) );
  and2_1 U13791 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [1]), .ip2(n12041), 
        .op(n11917) );
  ab_or_c_or_d U13792 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [1]), .ip2(n11924), .ip3(n11918), .ip4(n11917), .op(n6137) );
  nand2_1 U13793 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [2]), .ip2(n12041), 
        .op(n11923) );
  inv_1 U13794 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [2]), .op(n11920) );
  nand2_1 U13795 ( .ip1(n11918), .ip2(n11920), .op(n11932) );
  or2_1 U13796 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [1]), .ip2(n11924), .op(
        n11919) );
  inv_1 U13797 ( .ip(n11974), .op(n12042) );
  or2_1 U13798 ( .ip1(n12042), .ip2(n11924), .op(n12036) );
  nand2_1 U13799 ( .ip1(n11919), .ip2(n12036), .op(n11921) );
  or2_1 U13800 ( .ip1(n11921), .ip2(n11920), .op(n11922) );
  nand3_1 U13801 ( .ip1(n11923), .ip2(n11932), .ip3(n11922), .op(n6136) );
  or2_1 U13802 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [1]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [2]), .op(n11925) );
  or2_1 U13803 ( .ip1(n11925), .ip2(n11924), .op(n11926) );
  nand2_1 U13804 ( .ip1(n12036), .ip2(n11926), .op(n11931) );
  mux2_1 U13805 ( .ip1(n11932), .ip2(n11931), .s(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [3]), .op(n11928) );
  nand2_1 U13806 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [3]), .ip2(n12041), 
        .op(n11927) );
  nand2_1 U13807 ( .ip1(n11928), .ip2(n11927), .op(n6135) );
  nand2_1 U13808 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [3]), .ip2(n11929), 
        .op(n11930) );
  nand2_1 U13809 ( .ip1(n11931), .ip2(n11930), .op(n11935) );
  nor3_1 U13810 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [4]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [3]), .ip3(n11932), .op(n11934) );
  and2_1 U13811 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [4]), .ip2(n12041), 
        .op(n11933) );
  ab_or_c_or_d U13812 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [4]), .ip2(n11935), .ip3(n11934), .ip4(n11933), .op(n6134) );
  nand2_1 U13813 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [5]), .ip2(n12041), 
        .op(n11939) );
  nand2_1 U13814 ( .ip1(n11934), .ip2(n11937), .op(n11940) );
  or2_1 U13815 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [4]), .ip2(n11935), .op(
        n11936) );
  nand2_1 U13816 ( .ip1(n11936), .ip2(n12036), .op(n11948) );
  or2_1 U13817 ( .ip1(n11948), .ip2(n11937), .op(n11938) );
  nand3_1 U13818 ( .ip1(n11939), .ip2(n11940), .ip3(n11938), .op(n6133) );
  nor2_1 U13819 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [6]), .ip2(n11940), 
        .op(n11950) );
  or2_1 U13820 ( .ip1(n11948), .ip2(n11941), .op(n11944) );
  nand2_1 U13821 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [5]), .ip2(n12042), 
        .op(n11942) );
  or2_1 U13822 ( .ip1(n11942), .ip2(n11941), .op(n11943) );
  nand2_1 U13823 ( .ip1(n11944), .ip2(n11943), .op(n11945) );
  ab_or_c_or_d U13824 ( .ip1(n12041), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [6]), .ip3(n11950), .ip4(n11945), .op(n6132) );
  nand2_1 U13825 ( .ip1(n12042), .ip2(n11946), .op(n11947) );
  nand2_1 U13826 ( .ip1(n11948), .ip2(n11947), .op(n11954) );
  nand2_1 U13827 ( .ip1(n11954), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [7]), 
        .op(n11952) );
  nand2_1 U13828 ( .ip1(n12041), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [7]), 
        .op(n11951) );
  nand2_1 U13829 ( .ip1(n11950), .ip2(n11949), .op(n11953) );
  nand3_1 U13830 ( .ip1(n11952), .ip2(n11951), .ip3(n11953), .op(n6131) );
  nor2_1 U13831 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [8]), .ip2(n11953), 
        .op(n11957) );
  or2_1 U13832 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [7]), .ip2(n11954), .op(
        n11955) );
  nand2_1 U13833 ( .ip1(n11955), .ip2(n12036), .op(n11976) );
  inv_1 U13834 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [8]), .op(n11963) );
  nor2_1 U13835 ( .ip1(n11976), .ip2(n11963), .op(n11956) );
  ab_or_c_or_d U13836 ( .ip1(n12041), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [8]), .ip3(n11957), .ip4(n11956), .op(n6130) );
  nand2_1 U13837 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [9]), .ip2(n12041), 
        .op(n11961) );
  inv_1 U13838 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [9]), .op(n11964) );
  nand2_1 U13839 ( .ip1(n11957), .ip2(n11964), .op(n11962) );
  nand2_1 U13840 ( .ip1(n12042), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [8]), 
        .op(n11958) );
  nand2_1 U13841 ( .ip1(n11976), .ip2(n11958), .op(n11959) );
  nand2_1 U13842 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [9]), .ip2(n11959), 
        .op(n11960) );
  nand3_1 U13843 ( .ip1(n11961), .ip2(n11962), .ip3(n11960), .op(n6129) );
  nor2_1 U13844 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [10]), .ip2(n11962), 
        .op(n11972) );
  inv_1 U13845 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [10]), .op(n11966) );
  or2_1 U13846 ( .ip1(n11976), .ip2(n11966), .op(n11969) );
  nand2_1 U13847 ( .ip1(n11964), .ip2(n11963), .op(n11965) );
  nand2_1 U13848 ( .ip1(n12042), .ip2(n11965), .op(n11967) );
  or2_1 U13849 ( .ip1(n11967), .ip2(n11966), .op(n11968) );
  nand2_1 U13850 ( .ip1(n11969), .ip2(n11968), .op(n11970) );
  ab_or_c_or_d U13851 ( .ip1(n12041), .ip2(
        \CORTEXM0DS_INST/u_logic/Czh2z4 [10]), .ip3(n11972), .ip4(n11970), 
        .op(n6128) );
  nand2_1 U13852 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [11]), .ip2(n12041), 
        .op(n11978) );
  inv_1 U13853 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [11]), .op(n11971) );
  nand2_1 U13854 ( .ip1(n11972), .ip2(n11971), .op(n11979) );
  or2_1 U13855 ( .ip1(n11974), .ip2(n11973), .op(n11975) );
  nand2_1 U13856 ( .ip1(n11976), .ip2(n11975), .op(n11980) );
  nand2_1 U13857 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [11]), .ip2(n11980), 
        .op(n11977) );
  nand3_1 U13858 ( .ip1(n11978), .ip2(n11979), .ip3(n11977), .op(n6127) );
  nor2_1 U13859 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [12]), .ip2(n11979), 
        .op(n11984) );
  or2_1 U13860 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [11]), .ip2(n11980), 
        .op(n11981) );
  nand2_1 U13861 ( .ip1(n11981), .ip2(n12036), .op(n11986) );
  inv_1 U13862 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [12]), .op(n11982) );
  nor2_1 U13863 ( .ip1(n11986), .ip2(n11982), .op(n11983) );
  ab_or_c_or_d U13864 ( .ip1(n12041), .ip2(
        \CORTEXM0DS_INST/u_logic/Czh2z4 [12]), .ip3(n11984), .ip4(n11983), 
        .op(n6126) );
  nand2_1 U13865 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [13]), .ip2(n12041), 
        .op(n11988) );
  nand2_1 U13866 ( .ip1(n11984), .ip2(n11994), .op(n11989) );
  nand2_1 U13867 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [12]), .ip2(n12042), 
        .op(n11985) );
  nand2_1 U13868 ( .ip1(n11986), .ip2(n11985), .op(n11996) );
  nand2_1 U13869 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [13]), .ip2(n11996), 
        .op(n11987) );
  nand3_1 U13870 ( .ip1(n11988), .ip2(n11989), .ip3(n11987), .op(n6125) );
  nor2_1 U13871 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [14]), .ip2(n11989), 
        .op(n11993) );
  or2_1 U13872 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [13]), .ip2(n11996), 
        .op(n11990) );
  nand2_1 U13873 ( .ip1(n11990), .ip2(n12036), .op(n11991) );
  inv_1 U13874 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [14]), .op(n11995) );
  nor2_1 U13875 ( .ip1(n11991), .ip2(n11995), .op(n11992) );
  ab_or_c_or_d U13876 ( .ip1(n12041), .ip2(
        \CORTEXM0DS_INST/u_logic/Czh2z4 [14]), .ip3(n11993), .ip4(n11992), 
        .op(n6124) );
  inv_1 U13877 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [15]), .op(n11999) );
  nand2_1 U13878 ( .ip1(n11993), .ip2(n11999), .op(n12004) );
  nand2_1 U13879 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [15]), .ip2(n12041), 
        .op(n12001) );
  nand2_1 U13880 ( .ip1(n11995), .ip2(n11994), .op(n11997) );
  or2_1 U13881 ( .ip1(n11997), .ip2(n11996), .op(n11998) );
  nand2_1 U13882 ( .ip1(n12036), .ip2(n11998), .op(n12003) );
  or2_1 U13883 ( .ip1(n11999), .ip2(n12003), .op(n12000) );
  nand3_1 U13884 ( .ip1(n12004), .ip2(n12001), .ip3(n12000), .op(n6123) );
  nand2_1 U13885 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [15]), .ip2(n12042), 
        .op(n12002) );
  nand2_1 U13886 ( .ip1(n12003), .ip2(n12002), .op(n12013) );
  nor2_1 U13887 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [16]), .ip2(n12004), 
        .op(n12006) );
  and2_1 U13888 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [16]), .ip2(n12041), 
        .op(n12005) );
  ab_or_c_or_d U13889 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [16]), .ip2(
        n12013), .ip3(n12006), .ip4(n12005), .op(n6122) );
  nand2_1 U13890 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [17]), .ip2(n12041), 
        .op(n12011) );
  inv_1 U13891 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [17]), .op(n12008) );
  nand2_1 U13892 ( .ip1(n12006), .ip2(n12008), .op(n12012) );
  or2_1 U13893 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [16]), .ip2(n12013), 
        .op(n12007) );
  nand2_1 U13894 ( .ip1(n12007), .ip2(n12036), .op(n12009) );
  or2_1 U13895 ( .ip1(n12009), .ip2(n12008), .op(n12010) );
  nand3_1 U13896 ( .ip1(n12011), .ip2(n12012), .ip3(n12010), .op(n6121) );
  nor2_1 U13897 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [18]), .ip2(n12012), 
        .op(n12021) );
  or2_1 U13898 ( .ip1(n12014), .ip2(n12013), .op(n12015) );
  nand2_1 U13899 ( .ip1(n12036), .ip2(n12015), .op(n12019) );
  inv_1 U13900 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [18]), .op(n12016) );
  nor2_1 U13901 ( .ip1(n12019), .ip2(n12016), .op(n12017) );
  ab_or_c_or_d U13902 ( .ip1(n12041), .ip2(
        \CORTEXM0DS_INST/u_logic/Czh2z4 [18]), .ip3(n12021), .ip4(n12017), 
        .op(n6120) );
  nand2_1 U13903 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [18]), .ip2(n12042), 
        .op(n12018) );
  nand2_1 U13904 ( .ip1(n12019), .ip2(n12018), .op(n12025) );
  nand2_1 U13905 ( .ip1(n12025), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [19]), 
        .op(n12023) );
  nand2_1 U13906 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [19]), .ip2(n12041), 
        .op(n12022) );
  inv_1 U13907 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [19]), .op(n12020) );
  nand2_1 U13908 ( .ip1(n12021), .ip2(n12020), .op(n12024) );
  nand3_1 U13909 ( .ip1(n12023), .ip2(n12022), .ip3(n12024), .op(n6119) );
  nor2_1 U13910 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [20]), .ip2(n12024), 
        .op(n12032) );
  or2_1 U13911 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [19]), .ip2(n12025), 
        .op(n12026) );
  nand2_1 U13912 ( .ip1(n12026), .ip2(n12036), .op(n12030) );
  inv_1 U13913 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [20]), .op(n12027) );
  nor2_1 U13914 ( .ip1(n12030), .ip2(n12027), .op(n12028) );
  ab_or_c_or_d U13915 ( .ip1(n12041), .ip2(
        \CORTEXM0DS_INST/u_logic/Czh2z4 [20]), .ip3(n12032), .ip4(n12028), 
        .op(n6118) );
  nand2_1 U13916 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [20]), .ip2(n12042), 
        .op(n12029) );
  nand2_1 U13917 ( .ip1(n12030), .ip2(n12029), .op(n12035) );
  nand2_1 U13918 ( .ip1(n12035), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [21]), 
        .op(n12034) );
  nand2_1 U13919 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [21]), .ip2(n12041), 
        .op(n12033) );
  nand2_1 U13920 ( .ip1(n12032), .ip2(n12031), .op(n12038) );
  nand3_1 U13921 ( .ip1(n12034), .ip2(n12033), .ip3(n12038), .op(n6117) );
  or2_1 U13922 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [21]), .ip2(n12035), 
        .op(n12037) );
  nand2_1 U13923 ( .ip1(n12037), .ip2(n12036), .op(n12044) );
  mux2_1 U13924 ( .ip1(n12038), .ip2(n12044), .s(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [22]), .op(n12040) );
  nand2_1 U13925 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [22]), .ip2(n12041), 
        .op(n12039) );
  nand2_1 U13926 ( .ip1(n12040), .ip2(n12039), .op(n6116) );
  nand2_1 U13927 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [23]), .ip2(n12041), 
        .op(n12047) );
  nand2_1 U13928 ( .ip1(n12042), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [22]), 
        .op(n12043) );
  nand2_1 U13929 ( .ip1(n12044), .ip2(n12043), .op(n12045) );
  nand2_1 U13930 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [23]), .ip2(n12045), 
        .op(n12046) );
  nand2_1 U13931 ( .ip1(n12047), .ip2(n12046), .op(n6115) );
  inv_1 U13932 ( .ip(n12048), .op(n12052) );
  nand2_1 U13933 ( .ip1(n12049), .ip2(n3276), .op(n12050) );
  nand3_1 U13934 ( .ip1(n12050), .ip2(n2328), .ip3(
        \CORTEXM0DS_INST/u_logic/R3hvx4 ), .op(n12051) );
  nand2_1 U13935 ( .ip1(n12052), .ip2(n12051), .op(n6113) );
  nor3_1 U13936 ( .ip1(n3231), .ip2(n2269), .ip3(n2270), .op(n12053) );
  nand4_1 U13937 ( .ip1(\CORTEXM0DS_INST/u_logic/Sx3wx4 ), .ip2(n2266), .ip3(
        n12053), .ip4(\CORTEXM0DS_INST/u_logic/O24wx4 ), .op(n12054) );
  nor2_1 U13938 ( .ip1(n12055), .ip2(n12054), .op(n12056) );
  or2_1 U13939 ( .ip1(SYSRESETREQ_top_out), .ip2(n12056), .op(n6112) );
  nand3_1 U13940 ( .ip1(n2216), .ip2(n2215), .ip3(n2214), .op(n6111) );
  inv_1 U13941 ( .ip(n2212), .op(n2213) );
  or2_1 U13942 ( .ip1(\CORTEXM0DS_INST/u_logic/V2qvx4 ), .ip2(n2208), .op(
        n12059) );
  inv_1 U13943 ( .ip(n2207), .op(n12057) );
  or2_1 U13944 ( .ip1(n12057), .ip2(n2208), .op(n12058) );
  nand2_1 U13945 ( .ip1(n12059), .ip2(n12058), .op(n12060) );
  or2_1 U13946 ( .ip1(n2211), .ip2(n12060), .op(n6110) );
  inv_1 U13947 ( .ip(n12064), .op(n12477) );
  nor2_1 U13948 ( .ip1(n12477), .ip2(n2204), .op(n12061) );
  nor2_1 U13949 ( .ip1(n12062), .ip2(n12061), .op(n6109) );
  and2_1 U13950 ( .ip1(n12063), .ip2(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .op(
        n12067) );
  not_ab_or_c_or_d U13951 ( .ip1(n3217), .ip2(n12065), .ip3(n5932), .ip4(
        n12064), .op(n12066) );
  or2_1 U13952 ( .ip1(n12067), .ip2(n12066), .op(n6108) );
  nand3_1 U13953 ( .ip1(n12648), .ip2(n2196), .ip3(n2211), .op(n12069) );
  nand2_1 U13954 ( .ip1(\CORTEXM0DS_INST/u_logic/H0gvx4 ), .ip2(n2197), .op(
        n12068) );
  nand2_1 U13955 ( .ip1(n12069), .ip2(n12068), .op(n6107) );
  nand2_1 U13956 ( .ip1(n2211), .ip2(n2196), .op(
        \CORTEXM0DS_INST/u_logic/Xmywx4 ) );
  inv_1 U13957 ( .ip(n5772), .op(n12073) );
  nand3_1 U13958 ( .ip1(n12072), .ip2(n12071), .ip3(n12070), .op(n12095) );
  nand4_1 U13959 ( .ip1(\CORTEXM0DS_INST/u_logic/Fuevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip3(n12073), .ip4(n12095), .op(
        n12082) );
  nor2_1 U13960 ( .ip1(n12588), .ip2(n12074), .op(n12076) );
  and2_1 U13961 ( .ip1(n12094), .ip2(\CORTEXM0DS_INST/u_logic/W49vx4 ), .op(
        n12075) );
  not_ab_or_c_or_d U13962 ( .ip1(\CORTEXM0DS_INST/u_logic/D69vx4 ), .ip2(
        n12101), .ip3(n12076), .ip4(n12075), .op(n12078) );
  inv_1 U13963 ( .ip(\CORTEXM0DS_INST/u_logic/Cq9vx4 ), .op(n12077) );
  mux2_1 U13964 ( .ip1(n12078), .ip2(n12077), .s(n5772), .op(n12081) );
  or2_1 U13965 ( .ip1(n12079), .ip2(n12106), .op(n12080) );
  nand3_1 U13966 ( .ip1(n12082), .ip2(n12081), .ip3(n12080), .op(n6106) );
  nor2_1 U13967 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n12104), .op(
        n12083) );
  nor2_1 U13968 ( .ip1(n12084), .ip2(n12083), .op(n12085) );
  nor4_1 U13969 ( .ip1(n12088), .ip2(n12087), .ip3(n12086), .ip4(n12085), .op(
        n12092) );
  not_ab_or_c_or_d U13970 ( .ip1(n12090), .ip2(n12089), .ip3(
        \CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip4(n12588), .op(n12091) );
  not_ab_or_c_or_d U13971 ( .ip1(n12093), .ip2(
        \CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip3(n12092), .ip4(n12091), .op(
        n12098) );
  nand2_1 U13972 ( .ip1(\CORTEXM0DS_INST/u_logic/P39vx4 ), .ip2(n12094), .op(
        n12097) );
  nand3_1 U13973 ( .ip1(\CORTEXM0DS_INST/u_logic/Vsevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip3(n12095), .op(n12096) );
  nand4_1 U13974 ( .ip1(n12099), .ip2(n12098), .ip3(n12097), .ip4(n12096), 
        .op(n12100) );
  or2_1 U13975 ( .ip1(\CORTEXM0DS_INST/u_logic/W49vx4 ), .ip2(n12100), .op(
        n12103) );
  or2_1 U13976 ( .ip1(n12101), .ip2(n12100), .op(n12102) );
  nand2_1 U13977 ( .ip1(n12103), .ip2(n12102), .op(n12105) );
  mux2_1 U13978 ( .ip1(n12105), .ip2(n12104), .s(n5772), .op(n12110) );
  inv_1 U13979 ( .ip(n12106), .op(n12107) );
  nand2_1 U13980 ( .ip1(n12108), .ip2(n12107), .op(n12109) );
  nand2_1 U13981 ( .ip1(n12110), .ip2(n12109), .op(n6105) );
  nand3_1 U13982 ( .ip1(n12648), .ip2(n12112), .ip3(n12111), .op(n12115) );
  nand2_1 U13983 ( .ip1(\CORTEXM0DS_INST/u_logic/I4gvx4 ), .ip2(n12113), .op(
        n12114) );
  nand2_1 U13984 ( .ip1(n12115), .ip2(n12114), .op(n6104) );
  not_ab_or_c_or_d U13985 ( .ip1(n12117), .ip2(n5639), .ip3(n5932), .ip4(
        n12116), .op(n12119) );
  or2_1 U13986 ( .ip1(n12119), .ip2(n12118), .op(n12120) );
  nand2_1 U13987 ( .ip1(n2135), .ip2(n12120), .op(n6103) );
  nand2_1 U13988 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n12121), .op(
        n12141) );
  not_ab_or_c_or_d U13989 ( .ip1(n12124), .ip2(n12123), .ip3(n10492), .ip4(
        n12122), .op(n12130) );
  or2_1 U13990 ( .ip1(n12126), .ip2(n12125), .op(n12127) );
  nand2_1 U13991 ( .ip1(n12128), .ip2(n12127), .op(n12129) );
  not_ab_or_c_or_d U13992 ( .ip1(n12132), .ip2(n12131), .ip3(n12130), .ip4(
        n12129), .op(n12140) );
  nand3_1 U13993 ( .ip1(n12133), .ip2(n12609), .ip3(n9807), .op(n12136) );
  nand2_1 U13994 ( .ip1(n12134), .ip2(n12655), .op(n12135) );
  nand2_1 U13995 ( .ip1(n12136), .ip2(n12135), .op(n12137) );
  nand2_1 U13996 ( .ip1(n12138), .ip2(n12137), .op(n12139) );
  nand3_1 U13997 ( .ip1(n12141), .ip2(n12140), .ip3(n12139), .op(n2134) );
  nor2_1 U13998 ( .ip1(n12142), .ip2(n12347), .op(n12147) );
  inv_1 U13999 ( .ip(n12270), .op(n12145) );
  inv_1 U14000 ( .ip(n12346), .op(n12143) );
  not_ab_or_c_or_d U14001 ( .ip1(n12145), .ip2(n12144), .ip3(n12143), .ip4(
        n12343), .op(n12146) );
  not_ab_or_c_or_d U14002 ( .ip1(n12352), .ip2(n12148), .ip3(n12147), .ip4(
        n12146), .op(\CORTEXM0DS_INST/u_logic/Y92wx4 ) );
  nor2_1 U14003 ( .ip1(\CORTEXM0DS_INST/u_logic/Y92wx4 ), .ip2(n12355), .op(
        n12151) );
  nor2_1 U14004 ( .ip1(n12149), .ip2(n12353), .op(n12150) );
  ab_or_c_or_d U14005 ( .ip1(n12359), .ip2(\CORTEXM0DS_INST/vis_pc [22]), 
        .ip3(n12151), .ip4(n12150), .op(n6101) );
  nand2_1 U14006 ( .ip1(\CORTEXM0DS_INST/u_logic/Jjdvx4 ), .ip2(n2119), .op(
        n12153) );
  nand2_1 U14007 ( .ip1(\CORTEXM0DS_INST/vis_pc [14]), .ip2(n12359), .op(
        n12152) );
  nand3_1 U14008 ( .ip1(n12153), .ip2(n2094), .ip3(n12152), .op(n6100) );
  not_ab_or_c_or_d U14009 ( .ip1(n12333), .ip2(n12154), .ip3(n12162), .ip4(
        n12343), .op(n12157) );
  nor2_1 U14010 ( .ip1(n12155), .ip2(n12311), .op(n12156) );
  not_ab_or_c_or_d U14011 ( .ip1(n12316), .ip2(n12158), .ip3(n12157), .ip4(
        n12156), .op(\CORTEXM0DS_INST/u_logic/Z6ovx4 ) );
  nor2_1 U14012 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6ovx4 ), .ip2(n12355), .op(
        n12161) );
  nor2_1 U14013 ( .ip1(n12159), .ip2(n12353), .op(n12160) );
  ab_or_c_or_d U14014 ( .ip1(n12359), .ip2(\CORTEXM0DS_INST/vis_pc [7]), .ip3(
        n12161), .ip4(n12160), .op(n6099) );
  inv_1 U14015 ( .ip(n12162), .op(n12165) );
  inv_1 U14016 ( .ip(\CORTEXM0DS_INST/vis_pc [8]), .op(n12164) );
  nand2_1 U14017 ( .ip1(n12162), .ip2(\CORTEXM0DS_INST/vis_pc [8]), .op(n12175) );
  inv_1 U14018 ( .ip(n12175), .op(n12163) );
  not_ab_or_c_or_d U14019 ( .ip1(n12165), .ip2(n12164), .ip3(n12163), .ip4(
        n12343), .op(n12168) );
  nor2_1 U14020 ( .ip1(n12166), .ip2(n12347), .op(n12167) );
  not_ab_or_c_or_d U14021 ( .ip1(n12352), .ip2(n12169), .ip3(n12168), .ip4(
        n12167), .op(\CORTEXM0DS_INST/u_logic/Xxovx4 ) );
  nor2_1 U14022 ( .ip1(n12170), .ip2(n12353), .op(n12172) );
  nor2_1 U14023 ( .ip1(\CORTEXM0DS_INST/u_logic/Xxovx4 ), .ip2(n12355), .op(
        n12171) );
  not_ab_or_c_or_d U14024 ( .ip1(n12358), .ip2(
        \CORTEXM0DS_INST/u_logic/Oy8vx4 ), .ip3(n12172), .ip4(n12171), .op(
        n12174) );
  nand2_1 U14025 ( .ip1(\CORTEXM0DS_INST/vis_pc [8]), .ip2(n12359), .op(n12173) );
  nand2_1 U14026 ( .ip1(n12174), .ip2(n12173), .op(n6098) );
  inv_1 U14027 ( .ip(n12186), .op(n12184) );
  not_ab_or_c_or_d U14028 ( .ip1(n12176), .ip2(n12175), .ip3(n12184), .ip4(
        n12343), .op(n12179) );
  nor2_1 U14029 ( .ip1(n12177), .ip2(n12347), .op(n12178) );
  not_ab_or_c_or_d U14030 ( .ip1(n12352), .ip2(n12180), .ip3(n12179), .ip4(
        n12178), .op(\CORTEXM0DS_INST/u_logic/Jxovx4 ) );
  inv_1 U14031 ( .ip(\CORTEXM0DS_INST/u_logic/Jxovx4 ), .op(n2068) );
  nand2_1 U14032 ( .ip1(\CORTEXM0DS_INST/u_logic/Gcdvx4 ), .ip2(n2119), .op(
        n12183) );
  nand2_1 U14033 ( .ip1(n2118), .ip2(n2068), .op(n12182) );
  nand2_1 U14034 ( .ip1(\CORTEXM0DS_INST/vis_pc [9]), .ip2(n12359), .op(n12181) );
  nand3_1 U14035 ( .ip1(n12183), .ip2(n12182), .ip3(n12181), .op(n6097) );
  inv_1 U14036 ( .ip(\CORTEXM0DS_INST/vis_pc [10]), .op(n12187) );
  nand2_1 U14037 ( .ip1(\CORTEXM0DS_INST/vis_pc [10]), .ip2(n12184), .op(
        n12196) );
  inv_1 U14038 ( .ip(n12196), .op(n12185) );
  not_ab_or_c_or_d U14039 ( .ip1(n12187), .ip2(n12186), .ip3(n12185), .ip4(
        n12343), .op(n12190) );
  nor2_1 U14040 ( .ip1(n12188), .ip2(n12311), .op(n12189) );
  not_ab_or_c_or_d U14041 ( .ip1(n12316), .ip2(n12191), .ip3(n12190), .ip4(
        n12189), .op(\CORTEXM0DS_INST/u_logic/Owovx4 ) );
  inv_1 U14042 ( .ip(\CORTEXM0DS_INST/u_logic/Owovx4 ), .op(n2064) );
  nand2_1 U14043 ( .ip1(\CORTEXM0DS_INST/u_logic/Rddvx4 ), .ip2(n2119), .op(
        n12194) );
  nand2_1 U14044 ( .ip1(n2118), .ip2(n2064), .op(n12193) );
  nand2_1 U14045 ( .ip1(\CORTEXM0DS_INST/vis_pc [10]), .ip2(n12359), .op(
        n12192) );
  nand3_1 U14046 ( .ip1(n12194), .ip2(n12193), .ip3(n12192), .op(n6096) );
  not_ab_or_c_or_d U14047 ( .ip1(n12197), .ip2(n12196), .ip3(n12195), .ip4(
        n12343), .op(n12200) );
  nor2_1 U14048 ( .ip1(n12198), .ip2(n12311), .op(n12199) );
  not_ab_or_c_or_d U14049 ( .ip1(n12316), .ip2(n12201), .ip3(n12200), .ip4(
        n12199), .op(\CORTEXM0DS_INST/u_logic/Cqovx4 ) );
  nor2_1 U14050 ( .ip1(\CORTEXM0DS_INST/u_logic/Cqovx4 ), .ip2(n12355), .op(
        n12204) );
  nor2_1 U14051 ( .ip1(n12202), .ip2(n12353), .op(n12203) );
  ab_or_c_or_d U14052 ( .ip1(n12359), .ip2(\CORTEXM0DS_INST/vis_pc [11]), 
        .ip3(n12204), .ip4(n12203), .op(n6095) );
  nand2_1 U14053 ( .ip1(\CORTEXM0DS_INST/u_logic/Ngdvx4 ), .ip2(n2119), .op(
        n12206) );
  nand2_1 U14054 ( .ip1(\CORTEXM0DS_INST/vis_pc [12]), .ip2(n12359), .op(
        n12205) );
  nand3_1 U14055 ( .ip1(n12206), .ip2(n2059), .ip3(n12205), .op(n6094) );
  nand2_1 U14056 ( .ip1(\CORTEXM0DS_INST/u_logic/Yhdvx4 ), .ip2(n2119), .op(
        n12208) );
  nand2_1 U14057 ( .ip1(\CORTEXM0DS_INST/vis_pc [13]), .ip2(n12359), .op(
        n12207) );
  nand3_1 U14058 ( .ip1(n12208), .ip2(n2056), .ip3(n12207), .op(n6093) );
  inv_1 U14059 ( .ip(n12209), .op(n12212) );
  inv_1 U14060 ( .ip(n12221), .op(n12210) );
  not_ab_or_c_or_d U14061 ( .ip1(n12212), .ip2(n12211), .ip3(n12210), .ip4(
        n12343), .op(n12215) );
  nor2_1 U14062 ( .ip1(n12213), .ip2(n12311), .op(n12214) );
  not_ab_or_c_or_d U14063 ( .ip1(n12316), .ip2(n12216), .ip3(n12215), .ip4(
        n12214), .op(\CORTEXM0DS_INST/u_logic/Vpovx4 ) );
  nor2_1 U14064 ( .ip1(\CORTEXM0DS_INST/u_logic/Vpovx4 ), .ip2(n12355), .op(
        n12219) );
  nor2_1 U14065 ( .ip1(n12217), .ip2(n12353), .op(n12218) );
  ab_or_c_or_d U14066 ( .ip1(n12359), .ip2(\CORTEXM0DS_INST/vis_pc [15]), 
        .ip3(n12219), .ip4(n12218), .op(n6092) );
  not_ab_or_c_or_d U14067 ( .ip1(n12221), .ip2(n12220), .ip3(n12240), .ip4(
        n12343), .op(n12224) );
  nor2_1 U14068 ( .ip1(n12222), .ip2(n12311), .op(n12223) );
  not_ab_or_c_or_d U14069 ( .ip1(n12316), .ip2(n12225), .ip3(n12224), .ip4(
        n12223), .op(\CORTEXM0DS_INST/u_logic/Bv0wx4 ) );
  nor2_1 U14070 ( .ip1(\CORTEXM0DS_INST/u_logic/Bv0wx4 ), .ip2(n12355), .op(
        n12228) );
  nor2_1 U14071 ( .ip1(n12226), .ip2(n12353), .op(n12227) );
  ab_or_c_or_d U14072 ( .ip1(n12359), .ip2(\CORTEXM0DS_INST/vis_pc [16]), 
        .ip3(n12228), .ip4(n12227), .op(n6091) );
  inv_1 U14073 ( .ip(n12240), .op(n12230) );
  nand2_1 U14074 ( .ip1(\CORTEXM0DS_INST/vis_pc [17]), .ip2(n12240), .op(
        n12242) );
  inv_1 U14075 ( .ip(n12242), .op(n12229) );
  not_ab_or_c_or_d U14076 ( .ip1(n12231), .ip2(n12230), .ip3(n12229), .ip4(
        n12343), .op(n12234) );
  nor2_1 U14077 ( .ip1(n12232), .ip2(n12311), .op(n12233) );
  not_ab_or_c_or_d U14078 ( .ip1(n12316), .ip2(n12235), .ip3(n12234), .ip4(
        n12233), .op(\CORTEXM0DS_INST/u_logic/Fq0wx4 ) );
  nor2_1 U14079 ( .ip1(\CORTEXM0DS_INST/u_logic/Fq0wx4 ), .ip2(n12355), .op(
        n12238) );
  nor2_1 U14080 ( .ip1(n12236), .ip2(n12353), .op(n12237) );
  ab_or_c_or_d U14081 ( .ip1(n12359), .ip2(\CORTEXM0DS_INST/vis_pc [17]), 
        .ip3(n12238), .ip4(n12237), .op(n6090) );
  nor2_1 U14082 ( .ip1(n12239), .ip2(n12347), .op(n12245) );
  nand3_1 U14083 ( .ip1(\CORTEXM0DS_INST/vis_pc [17]), .ip2(
        \CORTEXM0DS_INST/vis_pc [18]), .ip3(n12240), .op(n12250) );
  inv_1 U14084 ( .ip(n12250), .op(n12241) );
  not_ab_or_c_or_d U14085 ( .ip1(n12243), .ip2(n12242), .ip3(n12241), .ip4(
        n12343), .op(n12244) );
  not_ab_or_c_or_d U14086 ( .ip1(n12352), .ip2(n12246), .ip3(n12245), .ip4(
        n12244), .op(\CORTEXM0DS_INST/u_logic/Ql0wx4 ) );
  nor2_1 U14087 ( .ip1(\CORTEXM0DS_INST/u_logic/Ql0wx4 ), .ip2(n12355), .op(
        n12249) );
  nor2_1 U14088 ( .ip1(n12247), .ip2(n12353), .op(n12248) );
  ab_or_c_or_d U14089 ( .ip1(n12359), .ip2(\CORTEXM0DS_INST/vis_pc [18]), 
        .ip3(n12249), .ip4(n12248), .op(n6089) );
  inv_1 U14090 ( .ip(n12261), .op(n12259) );
  not_ab_or_c_or_d U14091 ( .ip1(n12251), .ip2(n12250), .ip3(n12259), .ip4(
        n12343), .op(n12254) );
  nor2_1 U14092 ( .ip1(n12252), .ip2(n12311), .op(n12253) );
  not_ab_or_c_or_d U14093 ( .ip1(n12316), .ip2(n12255), .ip3(n12254), .ip4(
        n12253), .op(\CORTEXM0DS_INST/u_logic/Ug0wx4 ) );
  nor2_1 U14094 ( .ip1(\CORTEXM0DS_INST/u_logic/Ug0wx4 ), .ip2(n12355), .op(
        n12258) );
  nor2_1 U14095 ( .ip1(n12256), .ip2(n12353), .op(n12257) );
  ab_or_c_or_d U14096 ( .ip1(n12359), .ip2(\CORTEXM0DS_INST/vis_pc [19]), 
        .ip3(n12258), .ip4(n12257), .op(n6088) );
  inv_1 U14097 ( .ip(\CORTEXM0DS_INST/vis_pc [20]), .op(n12262) );
  nand2_1 U14098 ( .ip1(\CORTEXM0DS_INST/vis_pc [20]), .ip2(n12259), .op(
        n12271) );
  inv_1 U14099 ( .ip(n12271), .op(n12260) );
  not_ab_or_c_or_d U14100 ( .ip1(n12262), .ip2(n12261), .ip3(n12260), .ip4(
        n12343), .op(n12265) );
  nor2_1 U14101 ( .ip1(n12263), .ip2(n12311), .op(n12264) );
  not_ab_or_c_or_d U14102 ( .ip1(n12316), .ip2(n12266), .ip3(n12265), .ip4(
        n12264), .op(\CORTEXM0DS_INST/u_logic/Fc0wx4 ) );
  nor2_1 U14103 ( .ip1(\CORTEXM0DS_INST/u_logic/Fc0wx4 ), .ip2(n12355), .op(
        n12269) );
  nor2_1 U14104 ( .ip1(n12267), .ip2(n12353), .op(n12268) );
  ab_or_c_or_d U14105 ( .ip1(n12359), .ip2(\CORTEXM0DS_INST/vis_pc [20]), 
        .ip3(n12269), .ip4(n12268), .op(n6087) );
  not_ab_or_c_or_d U14106 ( .ip1(n12272), .ip2(n12271), .ip3(n12270), .ip4(
        n12343), .op(n12275) );
  nor2_1 U14107 ( .ip1(n12273), .ip2(n12347), .op(n12274) );
  not_ab_or_c_or_d U14108 ( .ip1(n12352), .ip2(n12276), .ip3(n12275), .ip4(
        n12274), .op(\CORTEXM0DS_INST/u_logic/C70wx4 ) );
  nor2_1 U14109 ( .ip1(\CORTEXM0DS_INST/u_logic/C70wx4 ), .ip2(n12355), .op(
        n12279) );
  nor2_1 U14110 ( .ip1(n12277), .ip2(n12353), .op(n12278) );
  ab_or_c_or_d U14111 ( .ip1(n12359), .ip2(\CORTEXM0DS_INST/vis_pc [21]), 
        .ip3(n12279), .ip4(n12278), .op(n6086) );
  not_ab_or_c_or_d U14112 ( .ip1(n12281), .ip2(n12280), .ip3(n12332), .ip4(
        n12343), .op(n12284) );
  nor2_1 U14113 ( .ip1(n12282), .ip2(n12311), .op(n12283) );
  not_ab_or_c_or_d U14114 ( .ip1(n12316), .ip2(n12285), .ip3(n12284), .ip4(
        n12283), .op(\CORTEXM0DS_INST/u_logic/Hszvx4 ) );
  nor2_1 U14115 ( .ip1(\CORTEXM0DS_INST/u_logic/Hszvx4 ), .ip2(n12355), .op(
        n12287) );
  and2_1 U14116 ( .ip1(\CORTEXM0DS_INST/vis_pc [5]), .ip2(n12359), .op(n12286)
         );
  ab_or_c_or_d U14117 ( .ip1(n2119), .ip2(\CORTEXM0DS_INST/u_logic/S6dvx4 ), 
        .ip3(n12287), .ip4(n12286), .op(n6082) );
  inv_1 U14118 ( .ip(n12288), .op(n12294) );
  inv_1 U14119 ( .ip(n12344), .op(n12290) );
  nor2_1 U14120 ( .ip1(n12290), .ip2(n12289), .op(n12298) );
  not_ab_or_c_or_d U14121 ( .ip1(n12290), .ip2(n12289), .ip3(n12298), .ip4(
        n12343), .op(n12293) );
  nor2_1 U14122 ( .ip1(n12291), .ip2(n12311), .op(n12292) );
  not_ab_or_c_or_d U14123 ( .ip1(n12316), .ip2(n12294), .ip3(n12293), .ip4(
        n12292), .op(\CORTEXM0DS_INST/u_logic/Rnovx4 ) );
  nor2_1 U14124 ( .ip1(\CORTEXM0DS_INST/u_logic/Rnovx4 ), .ip2(n12355), .op(
        n12297) );
  nor2_1 U14125 ( .ip1(n12295), .ip2(n12353), .op(n12296) );
  ab_or_c_or_d U14126 ( .ip1(n12359), .ip2(\CORTEXM0DS_INST/vis_pc [24]), 
        .ip3(n12297), .ip4(n12296), .op(n6081) );
  nor2_1 U14127 ( .ip1(\CORTEXM0DS_INST/vis_pc [25]), .ip2(n12298), .op(n12300) );
  inv_1 U14128 ( .ip(n12310), .op(n12299) );
  nor3_1 U14129 ( .ip1(n12300), .ip2(n12299), .ip3(n12343), .op(n12303) );
  nor2_1 U14130 ( .ip1(n12301), .ip2(n12311), .op(n12302) );
  not_ab_or_c_or_d U14131 ( .ip1(n12316), .ip2(n12304), .ip3(n12303), .ip4(
        n12302), .op(\CORTEXM0DS_INST/u_logic/Nhzvx4 ) );
  nor2_1 U14132 ( .ip1(\CORTEXM0DS_INST/u_logic/Nhzvx4 ), .ip2(n12355), .op(
        n12307) );
  nor2_1 U14133 ( .ip1(n12305), .ip2(n12353), .op(n12306) );
  ab_or_c_or_d U14134 ( .ip1(n12359), .ip2(\CORTEXM0DS_INST/vis_pc [25]), 
        .ip3(n12307), .ip4(n12306), .op(n6080) );
  not_ab_or_c_or_d U14135 ( .ip1(n12310), .ip2(n12309), .ip3(n12308), .ip4(
        n12343), .op(n12314) );
  nor2_1 U14136 ( .ip1(n12312), .ip2(n12311), .op(n12313) );
  not_ab_or_c_or_d U14137 ( .ip1(n12316), .ip2(n12315), .ip3(n12314), .ip4(
        n12313), .op(\CORTEXM0DS_INST/u_logic/Vezvx4 ) );
  nor2_1 U14138 ( .ip1(\CORTEXM0DS_INST/u_logic/Vezvx4 ), .ip2(n12355), .op(
        n12319) );
  nor2_1 U14139 ( .ip1(n12317), .ip2(n12353), .op(n12318) );
  ab_or_c_or_d U14140 ( .ip1(n12359), .ip2(\CORTEXM0DS_INST/vis_pc [26]), 
        .ip3(n12319), .ip4(n12318), .op(n6079) );
  or2_1 U14141 ( .ip1(\CORTEXM0DS_INST/cm0_xpsr[24] ), .ip2(n12323), .op(
        n12326) );
  nand3_1 U14142 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(n12320), .ip3(
        \CORTEXM0DS_INST/u_logic/Y99vx4 ), .op(n12322) );
  nand2_1 U14143 ( .ip1(n12322), .ip2(n12321), .op(n12324) );
  or2_1 U14144 ( .ip1(n12324), .ip2(n12323), .op(n12325) );
  nand2_1 U14145 ( .ip1(n12326), .ip2(n12325), .op(n12327) );
  nor2_1 U14146 ( .ip1(n12327), .ip2(n12355), .op(n12330) );
  nor2_1 U14147 ( .ip1(n12328), .ip2(n12353), .op(n12329) );
  ab_or_c_or_d U14148 ( .ip1(n12358), .ip2(\CORTEXM0DS_INST/vis_ipsr [0]), 
        .ip3(n12330), .ip4(n12329), .op(n6076) );
  nor2_1 U14149 ( .ip1(n12331), .ip2(n12347), .op(n12338) );
  inv_1 U14150 ( .ip(n12332), .op(n12336) );
  inv_1 U14151 ( .ip(n12333), .op(n12334) );
  not_ab_or_c_or_d U14152 ( .ip1(n12336), .ip2(n12335), .ip3(n12334), .ip4(
        n12343), .op(n12337) );
  not_ab_or_c_or_d U14153 ( .ip1(n12352), .ip2(n12339), .ip3(n12338), .ip4(
        n12337), .op(\CORTEXM0DS_INST/u_logic/S4qvx4 ) );
  nor2_1 U14154 ( .ip1(\CORTEXM0DS_INST/u_logic/S4qvx4 ), .ip2(n12355), .op(
        n12342) );
  nor2_1 U14155 ( .ip1(n12340), .ip2(n12353), .op(n12341) );
  ab_or_c_or_d U14156 ( .ip1(n12359), .ip2(\CORTEXM0DS_INST/vis_pc [6]), .ip3(
        n12342), .ip4(n12341), .op(n6074) );
  not_ab_or_c_or_d U14157 ( .ip1(n12346), .ip2(n12345), .ip3(n12344), .ip4(
        n12343), .op(n12350) );
  nor2_1 U14158 ( .ip1(n12348), .ip2(n12347), .op(n12349) );
  not_ab_or_c_or_d U14159 ( .ip1(n12352), .ip2(n12351), .ip3(n12350), .ip4(
        n12349), .op(\CORTEXM0DS_INST/u_logic/Y1pvx4 ) );
  nor2_1 U14160 ( .ip1(n12354), .ip2(n12353), .op(n12357) );
  nor2_1 U14161 ( .ip1(\CORTEXM0DS_INST/u_logic/Y1pvx4 ), .ip2(n12355), .op(
        n12356) );
  not_ab_or_c_or_d U14162 ( .ip1(\CORTEXM0DS_INST/cm0_xpsr[24] ), .ip2(n12358), 
        .ip3(n12357), .ip4(n12356), .op(n12361) );
  nand2_1 U14163 ( .ip1(\CORTEXM0DS_INST/vis_pc [23]), .ip2(n12359), .op(
        n12360) );
  nand2_1 U14164 ( .ip1(n12361), .ip2(n12360), .op(n6071) );
  nand2_1 U14165 ( .ip1(n12362), .ip2(n1769), .op(n12367) );
  nand2_1 U14166 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n12374), .op(
        n12365) );
  nand2_1 U14167 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(n12389), .op(
        n12364) );
  nand2_1 U14168 ( .ip1(\CORTEXM0DS_INST/u_logic/I29vx4 ), .ip2(n12375), .op(
        n12363) );
  nand4_1 U14169 ( .ip1(n12392), .ip2(n12365), .ip3(n12364), .ip4(n12363), 
        .op(n12366) );
  nand2_1 U14170 ( .ip1(n12367), .ip2(n12366), .op(n12372) );
  nor2_1 U14171 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n9807), .op(
        n12368) );
  nor2_1 U14172 ( .ip1(n12369), .ip2(n12368), .op(n12396) );
  nand2_1 U14173 ( .ip1(n12370), .ip2(n12396), .op(n12371) );
  nand2_1 U14174 ( .ip1(n12372), .ip2(n12371), .op(n6070) );
  nand2_1 U14175 ( .ip1(n12373), .ip2(n1769), .op(n12380) );
  nand2_1 U14176 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(n12374), .op(
        n12377) );
  nand2_1 U14177 ( .ip1(\CORTEXM0DS_INST/u_logic/B19vx4 ), .ip2(n12375), .op(
        n12376) );
  nand4_1 U14178 ( .ip1(n12392), .ip2(n12378), .ip3(n12377), .ip4(n12376), 
        .op(n12379) );
  nand2_1 U14179 ( .ip1(n12380), .ip2(n12379), .op(n12383) );
  nand2_1 U14180 ( .ip1(n12381), .ip2(n12396), .op(n12382) );
  nand2_1 U14181 ( .ip1(n12383), .ip2(n12382), .op(n6069) );
  nand2_1 U14182 ( .ip1(n12384), .ip2(n1769), .op(n12395) );
  nor2_1 U14183 ( .ip1(n12599), .ip2(n12385), .op(n12388) );
  nor2_1 U14184 ( .ip1(n12386), .ip2(n12592), .op(n12387) );
  not_ab_or_c_or_d U14185 ( .ip1(n12389), .ip2(
        \CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip3(n12388), .ip4(n12387), .op(
        n12393) );
  or2_1 U14186 ( .ip1(n12558), .ip2(n12390), .op(n12391) );
  nand3_1 U14187 ( .ip1(n12393), .ip2(n12392), .ip3(n12391), .op(n12394) );
  nand2_1 U14188 ( .ip1(n12395), .ip2(n12394), .op(n12399) );
  nand2_1 U14189 ( .ip1(n12397), .ip2(n12396), .op(n12398) );
  nand2_1 U14190 ( .ip1(n12399), .ip2(n12398), .op(n6068) );
  nand3_1 U14191 ( .ip1(n12401), .ip2(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip3(
        n12400), .op(n12405) );
  nand4_1 U14192 ( .ip1(n12403), .ip2(n12402), .ip3(n12409), .ip4(n12651), 
        .op(n12404) );
  nand2_1 U14193 ( .ip1(n12405), .ip2(n12404), .op(n12406) );
  nand3_1 U14194 ( .ip1(n12413), .ip2(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip3(
        n12406), .op(n12408) );
  nand2_1 U14195 ( .ip1(\CORTEXM0DS_INST/u_logic/Mk8vx4 ), .ip2(n1708), .op(
        n12407) );
  nand2_1 U14196 ( .ip1(n12408), .ip2(n12407), .op(n6066) );
  nand2_1 U14197 ( .ip1(n1708), .ip2(\CORTEXM0DS_INST/u_logic/Ul8vx4 ), .op(
        n12417) );
  nand2_1 U14198 ( .ip1(n12410), .ip2(n12409), .op(n12414) );
  nor2_1 U14199 ( .ip1(\CORTEXM0DS_INST/u_logic/Rkgvx4 ), .ip2(n12413), .op(
        n12411) );
  not_ab_or_c_or_d U14200 ( .ip1(n12414), .ip2(n12413), .ip3(n12412), .ip4(
        n12411), .op(n12415) );
  nand2_1 U14201 ( .ip1(n12415), .ip2(n12648), .op(n12416) );
  nand2_1 U14202 ( .ip1(n12417), .ip2(n12416), .op(n6065) );
  nand2_1 U14203 ( .ip1(n5932), .ip2(\CORTEXM0DS_INST/u_logic/N6hvx4 ), .op(
        n12426) );
  or2_1 U14204 ( .ip1(n1670), .ip2(n1671), .op(n12420) );
  nand3_1 U14205 ( .ip1(n1666), .ip2(n1667), .ip3(
        \CORTEXM0DS_INST/u_logic/Yuovx4 ), .op(n12418) );
  nand2_1 U14206 ( .ip1(n1669), .ip2(n12418), .op(n12419) );
  nand4_1 U14207 ( .ip1(n1674), .ip2(\CORTEXM0DS_INST/u_logic/Ekovx4 ), .ip3(
        n12420), .ip4(n12419), .op(n12422) );
  nand3_1 U14208 ( .ip1(n1671), .ip2(n1663), .ip3(n1662), .op(n12421) );
  not_ab_or_c_or_d U14209 ( .ip1(n12422), .ip2(n12421), .ip3(n1677), .ip4(
        n1676), .op(n12423) );
  and3_1 U14210 ( .ip1(\CORTEXM0DS_INST/u_logic/Rnovx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Vpovx4 ), .ip3(n12423), .op(n12427) );
  nand2_1 U14211 ( .ip1(n12427), .ip2(n1943), .op(n12424) );
  nand2_1 U14212 ( .ip1(n3128), .ip2(n12424), .op(n12425) );
  nand2_1 U14213 ( .ip1(n12426), .ip2(n12425), .op(n6064) );
  inv_1 U14214 ( .ip(n3128), .op(n12431) );
  nor2_1 U14215 ( .ip1(n12427), .ip2(n12431), .op(n12435) );
  nor2_1 U14216 ( .ip1(\CORTEXM0DS_INST/u_logic/Ekovx4 ), .ip2(n1690), .op(
        n12428) );
  not_ab_or_c_or_d U14217 ( .ip1(\CORTEXM0DS_INST/u_logic/Ekovx4 ), .ip2(n1690), .ip3(n12428), .ip4(n12431), .op(n12429) );
  ab_or_c_or_d U14218 ( .ip1(\CORTEXM0DS_INST/u_logic/Z7hvx4 ), .ip2(n5932), 
        .ip3(n12435), .ip4(n12429), .op(n6063) );
  nor2_1 U14219 ( .ip1(n1686), .ip2(n12431), .op(n12430) );
  ab_or_c_or_d U14220 ( .ip1(\CORTEXM0DS_INST/u_logic/L9hvx4 ), .ip2(n5932), 
        .ip3(n12435), .ip4(n12430), .op(n6062) );
  nor2_1 U14221 ( .ip1(n1684), .ip2(n12431), .op(n12432) );
  ab_or_c_or_d U14222 ( .ip1(\CORTEXM0DS_INST/u_logic/Xahvx4 ), .ip2(n5932), 
        .ip3(n12435), .ip4(n12432), .op(n6061) );
  nor2_1 U14223 ( .ip1(n12648), .ip2(n12433), .op(n12434) );
  ab_or_c_or_d U14224 ( .ip1(n3128), .ip2(\CORTEXM0DS_INST/u_logic/Z6ovx4 ), 
        .ip3(n12435), .ip4(n12434), .op(n6060) );
  mux2_1 U14225 ( .ip1(n2211), .ip2(\CORTEXM0DS_INST/u_logic/Xyfvx4 ), .s(
        n5932), .op(n6059) );
  nor2_1 U14226 ( .ip1(n5932), .ip2(n12436), .op(n12437) );
  nor2_1 U14227 ( .ip1(\CORTEXM0DS_INST/cm0_primask[0] ), .ip2(n12437), .op(
        n12438) );
  not_ab_or_c_or_d U14228 ( .ip1(n12439), .ip2(n12648), .ip3(1'b0), .ip4(
        n12438), .op(n6058) );
  nand2_1 U14229 ( .ip1(n12462), .ip2(n12477), .op(n12441) );
  nor2_1 U14230 ( .ip1(n12477), .ip2(n12519), .op(n12450) );
  nand2_1 U14231 ( .ip1(\CORTEXM0DS_INST/u_logic/Hnevx4 ), .ip2(n12450), .op(
        n12440) );
  nand3_1 U14232 ( .ip1(n12441), .ip2(n1514), .ip3(n12440), .op(n6057) );
  nand2_1 U14233 ( .ip1(n12477), .ip2(n12458), .op(n12443) );
  nand2_1 U14234 ( .ip1(n12450), .ip2(\CORTEXM0DS_INST/u_logic/Roevx4 ), .op(
        n12442) );
  nand3_1 U14235 ( .ip1(n12443), .ip2(n1509), .ip3(n12442), .op(n6056) );
  nand2_1 U14236 ( .ip1(n12470), .ip2(n12477), .op(n12445) );
  nand2_1 U14237 ( .ip1(n12450), .ip2(\CORTEXM0DS_INST/u_logic/Bqevx4 ), .op(
        n12444) );
  nand3_1 U14238 ( .ip1(n12445), .ip2(n1505), .ip3(n12444), .op(n6055) );
  nand2_1 U14239 ( .ip1(n12471), .ip2(n12477), .op(n12447) );
  nand2_1 U14240 ( .ip1(n12450), .ip2(\CORTEXM0DS_INST/u_logic/Lrevx4 ), .op(
        n12446) );
  nand3_1 U14241 ( .ip1(n12447), .ip2(n1504), .ip3(n12446), .op(n6054) );
  nand2_1 U14242 ( .ip1(n12457), .ip2(n12477), .op(n12449) );
  nand2_1 U14243 ( .ip1(n12450), .ip2(\CORTEXM0DS_INST/u_logic/Vsevx4 ), .op(
        n12448) );
  nand3_1 U14244 ( .ip1(n12449), .ip2(n1500), .ip3(n12448), .op(n6053) );
  nand2_1 U14245 ( .ip1(n12450), .ip2(\CORTEXM0DS_INST/u_logic/Fuevx4 ), .op(
        n12451) );
  nand2_1 U14246 ( .ip1(n1496), .ip2(n12451), .op(n6052) );
  inv_1 U14247 ( .ip(n4806), .op(n12517) );
  nand2_1 U14248 ( .ip1(\CORTEXM0DS_INST/u_logic/Pvevx4 ), .ip2(n12517), .op(
        n12479) );
  nor2_1 U14249 ( .ip1(\CORTEXM0DS_INST/u_logic/Pvevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Zwevx4 ), .op(n12480) );
  inv_1 U14250 ( .ip(n12480), .op(n12485) );
  inv_1 U14251 ( .ip(\CORTEXM0DS_INST/u_logic/O2fvx4 ), .op(n12594) );
  inv_1 U14252 ( .ip(\CORTEXM0DS_INST/u_logic/D1fvx4 ), .op(n12587) );
  inv_1 U14253 ( .ip(\CORTEXM0DS_INST/u_logic/Tzevx4 ), .op(n12582) );
  inv_1 U14254 ( .ip(\CORTEXM0DS_INST/u_logic/Jyevx4 ), .op(n12576) );
  nand4_1 U14255 ( .ip1(n12594), .ip2(n12587), .ip3(n12582), .ip4(n12576), 
        .op(n12452) );
  nor4_1 U14256 ( .ip1(\CORTEXM0DS_INST/u_logic/Z3fvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/K5fvx4 ), .ip3(n12485), .ip4(n12452), .op(
        n12454) );
  nor2_1 U14257 ( .ip1(n12454), .ip2(n12453), .op(n12650) );
  inv_1 U14258 ( .ip(\CORTEXM0DS_INST/u_logic/Pvevx4 ), .op(n12566) );
  nor2_1 U14259 ( .ip1(n12457), .ip2(n12456), .op(n12455) );
  not_ab_or_c_or_d U14260 ( .ip1(n12457), .ip2(n12456), .ip3(
        \CORTEXM0DS_INST/u_logic/Fuevx4 ), .ip4(n12455), .op(n12475) );
  inv_1 U14261 ( .ip(n12458), .op(n12469) );
  nor2_1 U14262 ( .ip1(n12462), .ip2(n12459), .op(n12468) );
  or2_1 U14263 ( .ip1(n12462), .ip2(n12458), .op(n12461) );
  or2_1 U14264 ( .ip1(n12459), .ip2(n12458), .op(n12460) );
  nand2_1 U14265 ( .ip1(n12461), .ip2(n12460), .op(n12466) );
  or2_1 U14266 ( .ip1(n12462), .ip2(n12547), .op(n12464) );
  inv_1 U14267 ( .ip(\CORTEXM0DS_INST/u_logic/Hnevx4 ), .op(n12543) );
  or2_1 U14268 ( .ip1(n12543), .ip2(n12547), .op(n12463) );
  nand2_1 U14269 ( .ip1(n12464), .ip2(n12463), .op(n12465) );
  nor2_1 U14270 ( .ip1(n12466), .ip2(n12465), .op(n12467) );
  not_ab_or_c_or_d U14271 ( .ip1(\CORTEXM0DS_INST/u_logic/Roevx4 ), .ip2(
        n12469), .ip3(n12468), .ip4(n12467), .op(n12474) );
  mux2_1 U14272 ( .ip1(n12553), .ip2(\CORTEXM0DS_INST/u_logic/Bqevx4 ), .s(
        n12470), .op(n12473) );
  inv_1 U14273 ( .ip(\CORTEXM0DS_INST/u_logic/Lrevx4 ), .op(n12557) );
  mux2_1 U14274 ( .ip1(n12557), .ip2(\CORTEXM0DS_INST/u_logic/Lrevx4 ), .s(
        n12471), .op(n12472) );
  nand4_1 U14275 ( .ip1(n12475), .ip2(n12474), .ip3(n12473), .ip4(n12472), 
        .op(n12476) );
  nand2_1 U14276 ( .ip1(n12477), .ip2(n12476), .op(n12514) );
  nand3_1 U14277 ( .ip1(n12650), .ip2(n12566), .ip3(n12514), .op(n12478) );
  nand3_1 U14278 ( .ip1(n12479), .ip2(n1494), .ip3(n12478), .op(n6051) );
  nand2_1 U14279 ( .ip1(n12517), .ip2(\CORTEXM0DS_INST/u_logic/Zwevx4 ), .op(
        n12484) );
  nand3_1 U14280 ( .ip1(\CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Zwevx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Pvevx4 ), .op(n12481) );
  nand2_1 U14281 ( .ip1(n12480), .ip2(n12650), .op(n12486) );
  nand2_1 U14282 ( .ip1(n12481), .ip2(n12486), .op(n12482) );
  nand2_1 U14283 ( .ip1(n12514), .ip2(n12482), .op(n12483) );
  nand3_1 U14284 ( .ip1(n12484), .ip2(n1490), .ip3(n12483), .op(n6050) );
  nand2_1 U14285 ( .ip1(n12517), .ip2(\CORTEXM0DS_INST/u_logic/Jyevx4 ), .op(
        n12490) );
  nand3_1 U14286 ( .ip1(n12485), .ip2(\CORTEXM0DS_INST/u_logic/Jyevx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Xlevx4 ), .op(n12487) );
  nor2_1 U14287 ( .ip1(\CORTEXM0DS_INST/u_logic/Jyevx4 ), .ip2(n12486), .op(
        n12504) );
  inv_1 U14288 ( .ip(n12504), .op(n12491) );
  nand2_1 U14289 ( .ip1(n12487), .ip2(n12491), .op(n12488) );
  nand2_1 U14290 ( .ip1(n12514), .ip2(n12488), .op(n12489) );
  nand3_1 U14291 ( .ip1(n12490), .ip2(n1487), .ip3(n12489), .op(n6049) );
  nand2_1 U14292 ( .ip1(n12517), .ip2(\CORTEXM0DS_INST/u_logic/Tzevx4 ), .op(
        n12494) );
  nand2_1 U14293 ( .ip1(\CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Tzevx4 ), .op(n12502) );
  xor2_1 U14294 ( .ip1(n12491), .ip2(n12502), .op(n12492) );
  nand2_1 U14295 ( .ip1(n12514), .ip2(n12492), .op(n12493) );
  nand3_1 U14296 ( .ip1(n12494), .ip2(n1484), .ip3(n12493), .op(n6048) );
  nand2_1 U14297 ( .ip1(n12517), .ip2(\CORTEXM0DS_INST/u_logic/D1fvx4 ), .op(
        n12498) );
  nand2_1 U14298 ( .ip1(n12504), .ip2(n12502), .op(n12495) );
  nand2_1 U14299 ( .ip1(\CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/D1fvx4 ), .op(n12503) );
  xor2_1 U14300 ( .ip1(n12495), .ip2(n12503), .op(n12496) );
  nand2_1 U14301 ( .ip1(n12514), .ip2(n12496), .op(n12497) );
  nand3_1 U14302 ( .ip1(n12498), .ip2(n1481), .ip3(n12497), .op(n6047) );
  nand2_1 U14303 ( .ip1(n12517), .ip2(\CORTEXM0DS_INST/u_logic/O2fvx4 ), .op(
        n12501) );
  nand3_1 U14304 ( .ip1(n12504), .ip2(n12502), .ip3(n12503), .op(n12509) );
  nand2_1 U14305 ( .ip1(\CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/O2fvx4 ), .op(n12511) );
  xor2_1 U14306 ( .ip1(n12509), .ip2(n12511), .op(n12499) );
  nand2_1 U14307 ( .ip1(n12514), .ip2(n12499), .op(n12500) );
  nand3_1 U14308 ( .ip1(n12501), .ip2(n1478), .ip3(n12500), .op(n6046) );
  nand2_1 U14309 ( .ip1(n12517), .ip2(\CORTEXM0DS_INST/u_logic/Z3fvx4 ), .op(
        n12508) );
  nand4_1 U14310 ( .ip1(n12504), .ip2(n12503), .ip3(n12502), .ip4(n12511), 
        .op(n12505) );
  nand2_1 U14311 ( .ip1(\CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Z3fvx4 ), .op(n12510) );
  xor2_1 U14312 ( .ip1(n12505), .ip2(n12510), .op(n12506) );
  nand2_1 U14313 ( .ip1(n12514), .ip2(n12506), .op(n12507) );
  nand3_1 U14314 ( .ip1(n12508), .ip2(n1475), .ip3(n12507), .op(n6045) );
  nand2_1 U14315 ( .ip1(n12517), .ip2(\CORTEXM0DS_INST/u_logic/K5fvx4 ), .op(
        n12516) );
  inv_1 U14316 ( .ip(n12509), .op(n12512) );
  nand3_1 U14317 ( .ip1(n12512), .ip2(n12511), .ip3(n12510), .op(n12513) );
  nand4_1 U14318 ( .ip1(\CORTEXM0DS_INST/u_logic/K5fvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip3(n12514), .ip4(n12513), .op(
        n12515) );
  nand3_1 U14319 ( .ip1(n12516), .ip2(n1472), .ip3(n12515), .op(n6044) );
  nand2_1 U14320 ( .ip1(n12517), .ip2(\CORTEXM0DS_INST/u_logic/V6fvx4 ), .op(
        n12518) );
  nand2_1 U14321 ( .ip1(n1402), .ip2(n12518), .op(n6043) );
  and2_1 U14322 ( .ip1(n12519), .ip2(n4807), .op(n1513) );
  nand2_1 U14323 ( .ip1(n1185), .ip2(\CORTEXM0DS_INST/u_logic/Cbfvx4 ), .op(
        n12520) );
  nand2_1 U14324 ( .ip1(n1187), .ip2(n12520), .op(n6041) );
  nand2_1 U14325 ( .ip1(n1185), .ip2(\CORTEXM0DS_INST/u_logic/Mcfvx4 ), .op(
        n12521) );
  nand2_1 U14326 ( .ip1(n1183), .ip2(n12521), .op(n6040) );
  nand2_1 U14327 ( .ip1(n1185), .ip2(\CORTEXM0DS_INST/u_logic/Wdfvx4 ), .op(
        n12522) );
  nand2_1 U14328 ( .ip1(n1181), .ip2(n12522), .op(n6039) );
  nand2_1 U14329 ( .ip1(n1185), .ip2(\CORTEXM0DS_INST/u_logic/Gffvx4 ), .op(
        n12523) );
  nand2_1 U14330 ( .ip1(n1179), .ip2(n12523), .op(n6038) );
  nand2_1 U14331 ( .ip1(n1185), .ip2(\CORTEXM0DS_INST/u_logic/Qgfvx4 ), .op(
        n12524) );
  nand2_1 U14332 ( .ip1(n1177), .ip2(n12524), .op(n6037) );
  nand2_1 U14333 ( .ip1(n1185), .ip2(\CORTEXM0DS_INST/u_logic/Aifvx4 ), .op(
        n12525) );
  nand2_1 U14334 ( .ip1(n1175), .ip2(n12525), .op(n6036) );
  nand2_1 U14335 ( .ip1(n1185), .ip2(\CORTEXM0DS_INST/u_logic/Kjfvx4 ), .op(
        n12526) );
  nand2_1 U14336 ( .ip1(n1173), .ip2(n12526), .op(n6035) );
  nand2_1 U14337 ( .ip1(n1185), .ip2(\CORTEXM0DS_INST/u_logic/Ukfvx4 ), .op(
        n12527) );
  nand2_1 U14338 ( .ip1(n1171), .ip2(n12527), .op(n6034) );
  nor2_1 U14339 ( .ip1(n1168), .ip2(n12535), .op(n12528) );
  mux2_1 U14340 ( .ip1(\CORTEXM0DS_INST/u_logic/Emfvx4 ), .ip2(n12528), .s(
        n12536), .op(n6033) );
  nand2_1 U14341 ( .ip1(n1185), .ip2(\CORTEXM0DS_INST/u_logic/Onfvx4 ), .op(
        n12529) );
  nand2_1 U14342 ( .ip1(n1167), .ip2(n12529), .op(n6032) );
  nand2_1 U14343 ( .ip1(n1185), .ip2(\CORTEXM0DS_INST/u_logic/Yofvx4 ), .op(
        n12530) );
  nand2_1 U14344 ( .ip1(n1165), .ip2(n12530), .op(n6031) );
  nand2_1 U14345 ( .ip1(n1185), .ip2(\CORTEXM0DS_INST/u_logic/Jqfvx4 ), .op(
        n12531) );
  nand2_1 U14346 ( .ip1(n1163), .ip2(n12531), .op(n6030) );
  nand2_1 U14347 ( .ip1(n1185), .ip2(\CORTEXM0DS_INST/u_logic/Urfvx4 ), .op(
        n12532) );
  nand2_1 U14348 ( .ip1(n1161), .ip2(n12532), .op(n6029) );
  nand2_1 U14349 ( .ip1(n1185), .ip2(\CORTEXM0DS_INST/u_logic/Ftfvx4 ), .op(
        n12533) );
  nand2_1 U14350 ( .ip1(n1159), .ip2(n12533), .op(n6028) );
  nor2_1 U14351 ( .ip1(n1185), .ip2(n12535), .op(n1184) );
  nor2_1 U14352 ( .ip1(n1156), .ip2(n12535), .op(n12534) );
  mux2_1 U14353 ( .ip1(\CORTEXM0DS_INST/u_logic/Qufvx4 ), .ip2(n12534), .s(
        n12536), .op(n6027) );
  nor2_1 U14354 ( .ip1(n1154), .ip2(n12535), .op(n12537) );
  mux2_1 U14355 ( .ip1(\CORTEXM0DS_INST/u_logic/Bwfvx4 ), .ip2(n12537), .s(
        n12536), .op(n6026) );
  and2_1 U14356 ( .ip1(\CORTEXM0DS_INST/u_logic/K5fvx4 ), .ip2(n12598), .op(
        n12540) );
  nor2_1 U14357 ( .ip1(n12600), .ip2(n12538), .op(n12539) );
  not_ab_or_c_or_d U14358 ( .ip1(n12603), .ip2(
        \CORTEXM0DS_INST/u_logic/Ftfvx4 ), .ip3(n12540), .ip4(n12539), .op(
        n12541) );
  nand3_1 U14359 ( .ip1(n1146), .ip2(n1144), .ip3(n12541), .op(n6024) );
  nor2_1 U14360 ( .ip1(n12600), .ip2(n12542), .op(n12545) );
  nor2_1 U14361 ( .ip1(n12543), .ip2(n12593), .op(n12544) );
  not_ab_or_c_or_d U14362 ( .ip1(n12603), .ip2(
        \CORTEXM0DS_INST/u_logic/Cbfvx4 ), .ip3(n12545), .ip4(n12544), .op(
        n12546) );
  nand3_1 U14363 ( .ip1(n1140), .ip2(n1138), .ip3(n12546), .op(n6023) );
  nor2_1 U14364 ( .ip1(n12547), .ip2(n12593), .op(n12550) );
  nor2_1 U14365 ( .ip1(n12600), .ip2(n12548), .op(n12549) );
  not_ab_or_c_or_d U14366 ( .ip1(n12603), .ip2(
        \CORTEXM0DS_INST/u_logic/Mcfvx4 ), .ip3(n12550), .ip4(n12549), .op(
        n12551) );
  nand3_1 U14367 ( .ip1(n1135), .ip2(n1133), .ip3(n12551), .op(n6022) );
  nor2_1 U14368 ( .ip1(n12600), .ip2(n12552), .op(n12555) );
  nor2_1 U14369 ( .ip1(n12553), .ip2(n12593), .op(n12554) );
  not_ab_or_c_or_d U14370 ( .ip1(n12603), .ip2(
        \CORTEXM0DS_INST/u_logic/Wdfvx4 ), .ip3(n12555), .ip4(n12554), .op(
        n12556) );
  nand3_1 U14371 ( .ip1(n1130), .ip2(n1128), .ip3(n12556), .op(n6021) );
  nor2_1 U14372 ( .ip1(n12557), .ip2(n12593), .op(n12560) );
  nor2_1 U14373 ( .ip1(n12600), .ip2(n12558), .op(n12559) );
  not_ab_or_c_or_d U14374 ( .ip1(n12603), .ip2(
        \CORTEXM0DS_INST/u_logic/Gffvx4 ), .ip3(n12560), .ip4(n12559), .op(
        n12561) );
  nand3_1 U14375 ( .ip1(n1125), .ip2(n1123), .ip3(n12561), .op(n6020) );
  and2_1 U14376 ( .ip1(\CORTEXM0DS_INST/u_logic/Fuevx4 ), .ip2(n12598), .op(
        n12564) );
  nor2_1 U14377 ( .ip1(n12600), .ip2(n12562), .op(n12563) );
  not_ab_or_c_or_d U14378 ( .ip1(n12603), .ip2(
        \CORTEXM0DS_INST/u_logic/Aifvx4 ), .ip3(n12564), .ip4(n12563), .op(
        n12565) );
  nand3_1 U14379 ( .ip1(n1115), .ip2(n1113), .ip3(n12565), .op(n6018) );
  nor2_1 U14380 ( .ip1(n12566), .ip2(n12593), .op(n12569) );
  nor2_1 U14381 ( .ip1(n12600), .ip2(n12567), .op(n12568) );
  not_ab_or_c_or_d U14382 ( .ip1(n12603), .ip2(
        \CORTEXM0DS_INST/u_logic/Kjfvx4 ), .ip3(n12569), .ip4(n12568), .op(
        n12570) );
  nand3_1 U14383 ( .ip1(n1110), .ip2(n1108), .ip3(n12570), .op(n6017) );
  nor2_1 U14384 ( .ip1(n12600), .ip2(n12571), .op(n12573) );
  and2_1 U14385 ( .ip1(\CORTEXM0DS_INST/u_logic/Zwevx4 ), .ip2(n12598), .op(
        n12572) );
  not_ab_or_c_or_d U14386 ( .ip1(n12603), .ip2(
        \CORTEXM0DS_INST/u_logic/Ukfvx4 ), .ip3(n12573), .ip4(n12572), .op(
        n12574) );
  nand3_1 U14387 ( .ip1(n1105), .ip2(n1103), .ip3(n12574), .op(n6016) );
  nand2_1 U14388 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n12575), .op(
        n12581) );
  nor2_1 U14389 ( .ip1(n12576), .ip2(n12593), .op(n12579) );
  nor2_1 U14390 ( .ip1(n1168), .ip2(n12577), .op(n12578) );
  not_ab_or_c_or_d U14391 ( .ip1(\CORTEXM0DS_INST/u_logic/Emfvx4 ), .ip2(
        n12603), .ip3(n12579), .ip4(n12578), .op(n12580) );
  nand3_1 U14392 ( .ip1(n12581), .ip2(n12580), .ip3(n1100), .op(n6015) );
  nor2_1 U14393 ( .ip1(n12582), .ip2(n12593), .op(n12585) );
  nor2_1 U14394 ( .ip1(n12600), .ip2(n12583), .op(n12584) );
  not_ab_or_c_or_d U14395 ( .ip1(n12603), .ip2(
        \CORTEXM0DS_INST/u_logic/Onfvx4 ), .ip3(n12585), .ip4(n12584), .op(
        n12586) );
  nand3_1 U14396 ( .ip1(n1095), .ip2(n1093), .ip3(n12586), .op(n6014) );
  nor2_1 U14397 ( .ip1(n12587), .ip2(n12593), .op(n12590) );
  nor2_1 U14398 ( .ip1(n12600), .ip2(n12588), .op(n12589) );
  not_ab_or_c_or_d U14399 ( .ip1(n12603), .ip2(
        \CORTEXM0DS_INST/u_logic/Yofvx4 ), .ip3(n12590), .ip4(n12589), .op(
        n12591) );
  nand3_1 U14400 ( .ip1(n1090), .ip2(n1088), .ip3(n12591), .op(n6013) );
  nor2_1 U14401 ( .ip1(n12600), .ip2(n12592), .op(n12596) );
  nor2_1 U14402 ( .ip1(n12594), .ip2(n12593), .op(n12595) );
  not_ab_or_c_or_d U14403 ( .ip1(n12603), .ip2(
        \CORTEXM0DS_INST/u_logic/Jqfvx4 ), .ip3(n12596), .ip4(n12595), .op(
        n12597) );
  nand3_1 U14404 ( .ip1(n1085), .ip2(n1083), .ip3(n12597), .op(n6012) );
  and2_1 U14405 ( .ip1(\CORTEXM0DS_INST/u_logic/Z3fvx4 ), .ip2(n12598), .op(
        n12602) );
  nor2_1 U14406 ( .ip1(n12600), .ip2(n12599), .op(n12601) );
  not_ab_or_c_or_d U14407 ( .ip1(n12603), .ip2(
        \CORTEXM0DS_INST/u_logic/Urfvx4 ), .ip3(n12602), .ip4(n12601), .op(
        n12604) );
  nand3_1 U14408 ( .ip1(n1080), .ip2(n1078), .ip3(n12604), .op(n6011) );
  or3_1 U14409 ( .ip1(n4578), .ip2(n12606), .ip3(n12605), .op(n12607) );
  nand2_1 U14410 ( .ip1(n1061), .ip2(n12607), .op(n6009) );
  nor2_1 U14411 ( .ip1(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip2(n12608), .op(
        n1059) );
  nand2_1 U14412 ( .ip1(n12618), .ip2(n12609), .op(n12616) );
  nand3_1 U14413 ( .ip1(n12610), .ip2(n12612), .ip3(n8424), .op(n12614) );
  nand2_1 U14414 ( .ip1(n12612), .ip2(n12611), .op(n12613) );
  nand4_1 U14415 ( .ip1(n12616), .ip2(n12615), .ip3(n12614), .ip4(n12613), 
        .op(n12640) );
  or2_1 U14416 ( .ip1(n12618), .ip2(n12617), .op(n12620) );
  nand2_1 U14417 ( .ip1(n12620), .ip2(n12619), .op(n12621) );
  nor2_1 U14418 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n12621), .op(
        n12639) );
  inv_1 U14419 ( .ip(n12622), .op(n12636) );
  nand2_1 U14420 ( .ip1(n12624), .ip2(n12623), .op(n12626) );
  nand2_1 U14421 ( .ip1(n12625), .ip2(n12626), .op(n12631) );
  nand2_1 U14422 ( .ip1(n12627), .ip2(n12626), .op(n12630) );
  inv_1 U14423 ( .ip(n12628), .op(n12629) );
  nand3_1 U14424 ( .ip1(n12631), .ip2(n12630), .ip3(n12629), .op(n12635) );
  nand2_1 U14425 ( .ip1(n12633), .ip2(n12632), .op(n12634) );
  nand4_1 U14426 ( .ip1(n12637), .ip2(n12636), .ip3(n12635), .ip4(n12634), 
        .op(n12638) );
  not_ab_or_c_or_d U14427 ( .ip1(n12641), .ip2(n12640), .ip3(n12639), .ip4(
        n12638), .op(n1060) );
  and2_1 U14428 ( .ip1(n12642), .ip2(\CORTEXM0DS_INST/u_logic/Mf8vx4 ), .op(
        n488) );
  mux2_1 U14429 ( .ip1(\CORTEXM0DS_INST/u_logic/Uth2z4 [1]), .ip2(n12644), .s(
        n488), .op(n6008) );
  nand2_1 U14430 ( .ip1(n12643), .ip2(\CORTEXM0DS_INST/u_logic/Mf8vx4 ), .op(
        n487) );
  mux2_1 U14431 ( .ip1(n12644), .ip2(\CORTEXM0DS_INST/u_logic/Txh2z4 [1]), .s(
        n487), .op(n6007) );
  mux2_1 U14432 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [23]), .ip2(n4704), .s(
        n12691), .op(n6006) );
  mux2_1 U14433 ( .ip1(n4704), .ip2(\CORTEXM0DS_INST/u_logic/Psh2z4 [1]), .s(
        n487), .op(n6005) );
  nor2_1 U14434 ( .ip1(\CORTEXM0DS_INST/u_logic/I4gvx4 ), .ip2(n12645), .op(
        n12646) );
  nor2_1 U14435 ( .ip1(n12647), .ip2(n12646), .op(n12649) );
  mux2_1 U14436 ( .ip1(\CORTEXM0DS_INST/u_logic/A3gvx4 ), .ip2(n12649), .s(
        n12648), .op(n6004) );
  mux2_1 U14437 ( .ip1(\CORTEXM0DS_INST/u_logic/Q5gvx4 ), .ip2(n12650), .s(
        n12651), .op(n6003) );
  mux2_1 U14438 ( .ip1(\CORTEXM0DS_INST/u_logic/Rkgvx4 ), .ip2(n12652), .s(
        n12651), .op(n6002) );
  nand3_1 U14439 ( .ip1(n12655), .ip2(n12654), .ip3(n12653), .op(n12658) );
  nand4_1 U14440 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip4(n12656), .op(n12657) );
  nand2_1 U14441 ( .ip1(n12658), .ip2(n12657), .op(n12659) );
  mux2_1 U14442 ( .ip1(n12659), .ip2(\CORTEXM0DS_INST/u_logic/Hx8vx4 ), .s(
        n5932), .op(n6001) );
  mux2_1 U14443 ( .ip1(n12660), .ip2(\CORTEXM0DS_INST/u_logic/Mxfvx4 ), .s(
        n1185), .op(n5999) );
  nand2_1 U14444 ( .ip1(n12661), .ip2(n12668), .op(n5997) );
  nand2_1 U14445 ( .ip1(n12662), .ip2(n12668), .op(n5995) );
  nand2_1 U14446 ( .ip1(n12663), .ip2(n12668), .op(n5993) );
  or2_1 U14447 ( .ip1(n12665), .ip2(n12664), .op(n5991) );
  nand2_1 U14448 ( .ip1(n12666), .ip2(n12668), .op(n5989) );
  nand2_1 U14449 ( .ip1(n12667), .ip2(n12668), .op(n5987) );
  nand2_1 U14450 ( .ip1(n12669), .ip2(n12668), .op(n5985) );
  or2_1 U14451 ( .ip1(n12684), .ip2(n12670), .op(n5983) );
  nand2_1 U14452 ( .ip1(n12671), .ip2(n12684), .op(n5984) );
  or2_1 U14453 ( .ip1(n12684), .ip2(n12672), .op(n5981) );
  nand2_1 U14454 ( .ip1(n12673), .ip2(n12684), .op(n5982) );
  or2_1 U14455 ( .ip1(n12684), .ip2(n12674), .op(n5979) );
  nand2_1 U14456 ( .ip1(n12675), .ip2(n12684), .op(n5980) );
  nand2_1 U14457 ( .ip1(n12683), .ip2(n12676), .op(n5977) );
  nand2_1 U14458 ( .ip1(n12677), .ip2(n12684), .op(n5978) );
  nand2_1 U14459 ( .ip1(n12683), .ip2(n12678), .op(n5975) );
  nand2_1 U14460 ( .ip1(n12679), .ip2(n12684), .op(n5976) );
  nand2_1 U14461 ( .ip1(n12683), .ip2(n12680), .op(n5973) );
  nand2_1 U14462 ( .ip1(n12681), .ip2(n12684), .op(n5974) );
  nand2_1 U14463 ( .ip1(n12683), .ip2(n12682), .op(n5971) );
  nand2_1 U14464 ( .ip1(n12685), .ip2(n12684), .op(n5972) );
  nor3_1 U14465 ( .ip1(n12689), .ip2(n12686), .ip3(n12687), .op(n2) );
  nor3_1 U14466 ( .ip1(n12689), .ip2(n12688), .ip3(n12687), .op(n1) );
  nor4_1 U14468 ( .ip1(PID_haddr_top[28]), .ip2(n2207), .ip3(n4578), .ip4(
        n2208), .op(n3128) );
  nor4_1 U14469 ( .ip1(PID_haddr_top[15]), .ip2(PID_haddr_top[16]), .ip3(n6111), .ip4(n5907), .op(n5925) );
  nand4_1 U14470 ( .ip1(HREADY_top), .ip2(n5014), .ip3(n5092), .ip4(n5013), 
        .op(n5420) );
  nand4_1 U14471 ( .ip1(HREADY_top), .ip2(PID_haddr_top[13]), .ip3(n5925), 
        .ip4(PID_haddr_top[12]), .op(n5924) );
  nor4_1 U14472 ( .ip1(PID_haddr_top[20]), .ip2(PID_haddr_top[19]), .ip3(
        PID_haddr_top[21]), .ip4(PID_haddr_top[18]), .op(n2216) );
  nor4_1 U14473 ( .ip1(PID_hwdata_top[26]), .ip2(PID_hwdata_top[22]), .ip3(
        PID_hwdata_top[18]), .ip4(PID_hwdata_top[19]), .op(n3229) );
  nor4_1 U14474 ( .ip1(PID_hwdata_top[16]), .ip2(PID_hwdata_top[28]), .ip3(
        PID_hwdata_top[24]), .ip4(PID_hwdata_top[17]), .op(n3228) );
  nor4_1 U14475 ( .ip1(PID_haddr_top[5]), .ip2(PID_haddr_top[10]), .ip3(
        PID_haddr_top[6]), .ip4(PID_haddr_top[11]), .op(n1667) );
  nand4_1 U14476 ( .ip1(\CORTEXM0DS_INST/u_logic/Cqovx4 ), .ip2(n2216), .ip3(
        PID_haddr_top[15]), .ip4(PID_hsize_top[1]), .op(n1676) );
  nor4_1 U14477 ( .ip1(PID_haddr_top[29]), .ip2(PID_haddr_top[30]), .ip3(
        PID_haddr_top[24]), .ip4(PID_haddr_top[22]), .op(n2215) );
  nand4_1 U14478 ( .ip1(PID_haddr_top[13]), .ip2(n2212), .ip3(
        PID_haddr_top[14]), .ip4(n1675), .op(n1677) );
  nor4_1 U14479 ( .ip1(PID_haddr_top[31]), .ip2(PID_haddr_top[28]), .ip3(
        PID_haddr_top[25]), .ip4(n2213), .op(n2214) );
  nor4_1 U14480 ( .ip1(PID_hwdata_top[20]), .ip2(PID_hwdata_top[21]), .ip3(
        n3231), .ip4(n3230), .op(n3233) );
  nand4_1 U14481 ( .ip1(PID_hwdata_top[2]), .ip2(PID_hwdata_top[21]), .ip3(
        PID_hwdata_top[20]), .ip4(n3227), .op(n2269) );
  nor2_1 U14482 ( .ip1(PID_hwdata_top[11]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [11]), .op(n12737) );
  nor2_1 U14483 ( .ip1(PID_hwdata_top[9]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [9]), .op(n12738) );
  nor2_1 U14484 ( .ip1(PID_hwdata_top[10]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [10]), .op(n12739) );
  nor2_1 U14485 ( .ip1(PID_hwdata_top[13]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [13]), .op(n12740) );
  nor2_1 U14486 ( .ip1(PID_hwdata_top[15]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [15]), .op(n12741) );
  nor2_1 U14487 ( .ip1(PID_hwdata_top[8]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [8]), .op(n12742) );
  nor2_1 U14488 ( .ip1(PID_hwdata_top[12]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [12]), .op(n12743) );
  nor2_1 U14489 ( .ip1(PID_hwdata_top[0]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [0]), .op(n12744) );
  nor2_1 U14490 ( .ip1(PID_hwdata_top[3]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [3]), .op(n12745) );
  nor2_1 U14491 ( .ip1(PID_hwdata_top[6]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [6]), .op(n12746) );
  nor2_1 U14492 ( .ip1(PID_hwdata_top[26]), .ip2(n2326), .op(n12747) );
  nor2_1 U14493 ( .ip1(PID_hwdata_top[7]), .ip2(n3223), .op(n12748) );
endmodule

