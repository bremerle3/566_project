
module i_i2c_DW_apb_i2c_regfile ( pclk, presetn, wr_en, rd_en, byte_en, 
        reg_addr, ipwdata, iprdata, ic_clr_intr_en, ic_clr_rx_under_en, 
        ic_clr_rx_over_en, ic_clr_tx_over_en, ic_clr_rd_req_en, 
        ic_clr_tx_abrt_en, ic_clr_rx_done_en, ic_clr_activity_en, 
        ic_clr_stop_det_en, ic_clr_start_det_en, ic_clr_gen_call_en, 
        mst_activity, slv_activity, activity, ic_tx_abrt_source, ic_en, 
        slv_rx_aborted_sync, slv_fifo_filled_and_flushed_sync, ic_tar, ic_sar, 
        ic_hs_maddr, ic_fs_hcnt, ic_fs_lcnt, ic_intr_mask, ic_rx_tl_int, 
        ic_enable, ic_hcnt, ic_lcnt, ic_fs_spklen, ic_hs_spklen, ic_intr_stat, 
        ic_raw_intr_stat, ic_hs, ic_fs, ic_ss, ic_master, ic_10bit_mst, 
        ic_10bit_slv, ic_slave_en, p_det_ifaddr, tx_empty_ctrl, rx_pop_data, 
        tx_push_data, fifo_rst_n, tx_fifo_rst_n, tx_pop_sync, rx_push_sync, 
        rx_pop, tx_push, tx_empty, rx_full, tx_full, rx_empty, tx_abrt_flg_edg, 
        abrt_in_rcve_trns, slv_clr_leftover_flg_edg, ic_rstrt_en, ic_sda_setup, 
        ic_sda_hold, ic_ack_general_call, ic_tx_tl_7_, ic_tx_tl_6_, 
        ic_tx_tl_5_, ic_tx_tl_4_, ic_tx_tl_3__BAR, ic_tx_tl_2_, ic_tx_tl_1_, 
        ic_tx_tl_0_ );
  input [3:0] byte_en;
  input [5:0] reg_addr;
  input [31:0] ipwdata;
  output [31:0] iprdata;
  input [16:0] ic_tx_abrt_source;
  output [11:0] ic_tar;
  output [9:0] ic_sar;
  output [2:0] ic_hs_maddr;
  output [15:0] ic_fs_hcnt;
  output [15:0] ic_fs_lcnt;
  output [13:0] ic_intr_mask;
  output [2:0] ic_rx_tl_int;
  output [1:0] ic_enable;
  output [15:0] ic_hcnt;
  output [15:0] ic_lcnt;
  output [7:0] ic_fs_spklen;
  output [7:0] ic_hs_spklen;
  input [13:0] ic_intr_stat;
  input [13:0] ic_raw_intr_stat;
  input [7:0] rx_pop_data;
  output [8:0] tx_push_data;
  output [7:0] ic_sda_setup;
  output [23:0] ic_sda_hold;
  input pclk, presetn, wr_en, rd_en, mst_activity, slv_activity, activity,
         ic_en, slv_rx_aborted_sync, slv_fifo_filled_and_flushed_sync,
         tx_pop_sync, rx_push_sync, tx_empty, rx_full, tx_full, rx_empty,
         tx_abrt_flg_edg, abrt_in_rcve_trns, slv_clr_leftover_flg_edg;
  output ic_clr_intr_en, ic_clr_rx_under_en, ic_clr_rx_over_en,
         ic_clr_tx_over_en, ic_clr_rd_req_en, ic_clr_tx_abrt_en,
         ic_clr_rx_done_en, ic_clr_activity_en, ic_clr_stop_det_en,
         ic_clr_start_det_en, ic_clr_gen_call_en, ic_hs, ic_fs, ic_ss,
         ic_master, ic_10bit_mst, ic_10bit_slv, ic_slave_en, p_det_ifaddr,
         tx_empty_ctrl, fifo_rst_n, tx_fifo_rst_n, rx_pop, tx_push,
         ic_rstrt_en, ic_ack_general_call, ic_tx_tl_7_, ic_tx_tl_6_,
         ic_tx_tl_5_, ic_tx_tl_4_, ic_tx_tl_3__BAR, ic_tx_tl_2_, ic_tx_tl_1_,
         ic_tx_tl_0_;
  wire   activity_r, mst_activity_r, slv_activity_r, ic_con_pre_6_,
         ic_con_pre_2_, ic_con_pre_1_, fifo_rst_n_int, fix_c, n1105, n1107,
         n1109, n1111, n1113, n1115, n1117, n1119, n1121, n1123, n1125, n1127,
         n1129, n1131, n1133, n1135, n1137, n1149, n1151, n1153, n1165, n1167,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n760;
  wire   [3:0] ic_txflr;
  wire   [3:0] ic_txflr_flushed;
  wire   [3:0] ic_rxflr;
  wire   [15:0] hcr_ic_ss_hcnt;
  wire   [15:0] hcr_ic_ss_lcnt;
  wire   [15:0] hcr_ic_hs_hcnt;
  wire   [15:0] hcr_ic_hs_lcnt;

  drp_1 mst_activity_r_reg ( .ip(mst_activity), .ck(pclk), .rb(presetn), .q(
        mst_activity_r) );
  drp_1 slv_activity_r_reg ( .ip(slv_activity), .ck(pclk), .rb(presetn), .q(
        slv_activity_r) );
  drp_1 activity_r_reg ( .ip(activity), .ck(pclk), .rb(presetn), .q(activity_r) );
  drp_1 ic_enable_reg_reg_0_ ( .ip(n1549), .ck(pclk), .rb(presetn), .q(
        ic_enable[0]) );
  drp_1 ic_enable_reg_reg_1_ ( .ip(n1548), .ck(pclk), .rb(presetn), .q(
        ic_enable[1]) );
  drp_1 ic_rxflr_reg_0_ ( .ip(n1546), .ck(pclk), .rb(presetn), .q(ic_rxflr[0])
         );
  drp_1 ic_rxflr_reg_2_ ( .ip(n1544), .ck(pclk), .rb(presetn), .q(ic_rxflr[2])
         );
  drp_1 ic_rxflr_reg_3_ ( .ip(n1547), .ck(pclk), .rb(presetn), .q(ic_rxflr[3])
         );
  drp_1 ic_rxflr_reg_1_ ( .ip(n1545), .ck(pclk), .rb(presetn), .q(ic_rxflr[1])
         );
  drp_1 ic_con_pre_reg_8_ ( .ip(n1543), .ck(pclk), .rb(presetn), .q(
        tx_empty_ctrl) );
  drp_1 ic_con_pre_reg_7_ ( .ip(n1542), .ck(pclk), .rb(presetn), .q(
        p_det_ifaddr) );
  drp_1 ic_tar_reg_reg_11_ ( .ip(n1529), .ck(pclk), .rb(presetn), .q(
        ic_tar[11]) );
  drp_1 ic_tar_reg_reg_10_ ( .ip(n1530), .ck(pclk), .rb(presetn), .q(
        ic_tar[10]) );
  drp_1 ic_tar_reg_reg_9_ ( .ip(n1531), .ck(pclk), .rb(presetn), .q(ic_tar[9])
         );
  drp_1 ic_tar_reg_reg_8_ ( .ip(n1532), .ck(pclk), .rb(presetn), .q(ic_tar[8])
         );
  drp_1 ic_tar_reg_reg_7_ ( .ip(n1513), .ck(pclk), .rb(presetn), .q(ic_tar[7])
         );
  drp_1 ic_tar_reg_reg_5_ ( .ip(n1515), .ck(pclk), .rb(presetn), .q(ic_tar[5])
         );
  drp_1 ic_tar_reg_reg_3_ ( .ip(n1517), .ck(pclk), .rb(presetn), .q(ic_tar[3])
         );
  drp_1 ic_tar_reg_reg_1_ ( .ip(n1519), .ck(pclk), .rb(presetn), .q(ic_tar[1])
         );
  drp_1 ic_sar_reg_9_ ( .ip(n1533), .ck(pclk), .rb(presetn), .q(ic_sar[9]) );
  drp_1 ic_sar_reg_8_ ( .ip(n1534), .ck(pclk), .rb(presetn), .q(ic_sar[8]) );
  drp_1 ic_sar_reg_7_ ( .ip(n1521), .ck(pclk), .rb(presetn), .q(ic_sar[7]) );
  drp_1 ic_sar_reg_5_ ( .ip(n1523), .ck(pclk), .rb(presetn), .q(ic_sar[5]) );
  drp_1 ic_sar_reg_3_ ( .ip(n1525), .ck(pclk), .rb(presetn), .q(ic_sar[3]) );
  drp_1 ic_sar_reg_1_ ( .ip(n1527), .ck(pclk), .rb(presetn), .q(ic_sar[1]) );
  drp_1 r_ic_ss_hcnt_reg_15_ ( .ip(n1504), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[15]) );
  drp_1 r_ic_ss_hcnt_reg_14_ ( .ip(n1497), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[14]) );
  drp_1 r_ic_ss_hcnt_reg_13_ ( .ip(n1498), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[13]) );
  drp_1 r_ic_ss_hcnt_reg_12_ ( .ip(n1499), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[12]) );
  drp_1 r_ic_ss_hcnt_reg_11_ ( .ip(n1500), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[11]) );
  drp_1 r_ic_ss_hcnt_reg_10_ ( .ip(n1501), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[10]) );
  drp_1 r_ic_ss_hcnt_reg_9_ ( .ip(n1502), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[9]) );
  drp_1 r_ic_ss_hcnt_reg_6_ ( .ip(n1506), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[6]) );
  drp_1 r_ic_ss_hcnt_reg_5_ ( .ip(n1507), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[5]) );
  drp_1 r_ic_ss_hcnt_reg_3_ ( .ip(n1509), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[3]) );
  drp_1 r_ic_ss_hcnt_reg_2_ ( .ip(n1510), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[2]) );
  drp_1 r_ic_ss_hcnt_reg_1_ ( .ip(n1511), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[1]) );
  drp_1 r_ic_ss_hcnt_reg_0_ ( .ip(n1512), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[0]) );
  drp_1 r_ic_ss_lcnt_reg_3_ ( .ip(n1493), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[3]) );
  drp_1 r_ic_ss_lcnt_reg_5_ ( .ip(n1491), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[5]) );
  drp_1 r_ic_ss_lcnt_reg_15_ ( .ip(n1488), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[15]) );
  drp_1 r_ic_ss_lcnt_reg_9_ ( .ip(n1486), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[9]) );
  drp_1 r_ic_ss_lcnt_reg_10_ ( .ip(n1485), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[10]) );
  drp_1 r_ic_ss_lcnt_reg_11_ ( .ip(n1484), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[11]) );
  drp_1 r_ic_ss_lcnt_reg_12_ ( .ip(n1483), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[12]) );
  drp_1 r_ic_ss_lcnt_reg_13_ ( .ip(n1482), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[13]) );
  drp_1 r_ic_ss_lcnt_reg_14_ ( .ip(n1481), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[14]) );
  drp_1 r_ic_ss_lcnt_reg_0_ ( .ip(n1496), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[0]) );
  drp_1 r_ic_fs_hcnt_reg_15_ ( .ip(n1472), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[15]) );
  drp_1 r_ic_fs_hcnt_reg_14_ ( .ip(n1465), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[14]) );
  drp_1 r_ic_fs_hcnt_reg_13_ ( .ip(n1466), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[13]) );
  drp_1 r_ic_fs_hcnt_reg_12_ ( .ip(n1467), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[12]) );
  drp_1 r_ic_fs_hcnt_reg_11_ ( .ip(n1468), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[11]) );
  drp_1 r_ic_fs_hcnt_reg_10_ ( .ip(n1469), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[10]) );
  drp_1 r_ic_fs_hcnt_reg_9_ ( .ip(n1470), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[9]) );
  drp_1 r_ic_fs_hcnt_reg_8_ ( .ip(n1471), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[8]) );
  drp_1 r_ic_fs_hcnt_reg_7_ ( .ip(n1473), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[7]) );
  drp_1 r_ic_fs_hcnt_reg_6_ ( .ip(n1474), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[6]) );
  drp_1 r_ic_fs_hcnt_reg_1_ ( .ip(n1479), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[1]) );
  drp_1 r_ic_fs_hcnt_reg_0_ ( .ip(n1480), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[0]) );
  drp_1 r_ic_fs_lcnt_reg_3_ ( .ip(n1461), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[3]) );
  drp_1 r_ic_fs_lcnt_reg_4_ ( .ip(n1460), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[4]) );
  drp_1 r_ic_fs_lcnt_reg_5_ ( .ip(n1459), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[5]) );
  drp_1 r_ic_fs_lcnt_reg_6_ ( .ip(n1458), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[6]) );
  drp_1 r_ic_fs_lcnt_reg_15_ ( .ip(n1456), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[15]) );
  drp_1 r_ic_fs_lcnt_reg_8_ ( .ip(n1455), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[8]) );
  drp_1 r_ic_fs_lcnt_reg_9_ ( .ip(n1454), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[9]) );
  drp_1 r_ic_fs_lcnt_reg_10_ ( .ip(n1453), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[10]) );
  drp_1 r_ic_fs_lcnt_reg_11_ ( .ip(n1452), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[11]) );
  drp_1 r_ic_fs_lcnt_reg_12_ ( .ip(n1451), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[12]) );
  drp_1 r_ic_fs_lcnt_reg_13_ ( .ip(n1450), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[13]) );
  drp_1 r_ic_fs_lcnt_reg_14_ ( .ip(n1449), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[14]) );
  drp_1 r_ic_fs_lcnt_reg_2_ ( .ip(n1462), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[2]) );
  drp_1 r_ic_fs_lcnt_reg_0_ ( .ip(n1464), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[0]) );
  drp_1 r_ic_hs_hcnt_reg_15_ ( .ip(n1440), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[15]) );
  drp_1 r_ic_hs_hcnt_reg_14_ ( .ip(n1433), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[14]) );
  drp_1 r_ic_hs_hcnt_reg_13_ ( .ip(n1434), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[13]) );
  drp_1 r_ic_hs_hcnt_reg_12_ ( .ip(n1435), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[12]) );
  drp_1 r_ic_hs_hcnt_reg_11_ ( .ip(n1436), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[11]) );
  drp_1 r_ic_hs_hcnt_reg_10_ ( .ip(n1437), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[10]) );
  drp_1 r_ic_hs_hcnt_reg_9_ ( .ip(n1438), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[9]) );
  drp_1 r_ic_hs_hcnt_reg_8_ ( .ip(n1439), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[8]) );
  drp_1 r_ic_hs_hcnt_reg_7_ ( .ip(n1441), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[7]) );
  drp_1 r_ic_hs_hcnt_reg_6_ ( .ip(n1442), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[6]) );
  drp_1 r_ic_hs_hcnt_reg_5_ ( .ip(n1443), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[5]) );
  drp_1 r_ic_hs_hcnt_reg_4_ ( .ip(n1444), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[4]) );
  drp_1 r_ic_hs_hcnt_reg_3_ ( .ip(n1445), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[3]) );
  drp_1 r_ic_hs_hcnt_reg_0_ ( .ip(n1448), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[0]) );
  drp_1 r_ic_hs_lcnt_reg_3_ ( .ip(n1429), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[3]) );
  drp_1 r_ic_hs_lcnt_reg_5_ ( .ip(n1427), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[5]) );
  drp_1 r_ic_hs_lcnt_reg_6_ ( .ip(n1426), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[6]) );
  drp_1 r_ic_hs_lcnt_reg_7_ ( .ip(n1425), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[7]) );
  drp_1 r_ic_hs_lcnt_reg_15_ ( .ip(n1424), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[15]) );
  drp_1 r_ic_hs_lcnt_reg_8_ ( .ip(n1423), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[8]) );
  drp_1 r_ic_hs_lcnt_reg_9_ ( .ip(n1422), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[9]) );
  drp_1 r_ic_hs_lcnt_reg_10_ ( .ip(n1421), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[10]) );
  drp_1 r_ic_hs_lcnt_reg_11_ ( .ip(n1420), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[11]) );
  drp_1 r_ic_hs_lcnt_reg_12_ ( .ip(n1419), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[12]) );
  drp_1 r_ic_hs_lcnt_reg_13_ ( .ip(n1418), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[13]) );
  drp_1 r_ic_hs_lcnt_reg_14_ ( .ip(n1417), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[14]) );
  drp_1 r_ic_hs_lcnt_reg_2_ ( .ip(n1430), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[2]) );
  drp_1 r_ic_hs_lcnt_reg_1_ ( .ip(n1431), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[1]) );
  drp_1 r_ic_hs_lcnt_reg_0_ ( .ip(n1432), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[0]) );
  drp_1 r_ic_fs_spklen_reg_7_ ( .ip(n1416), .ck(pclk), .rb(presetn), .q(
        ic_fs_spklen[7]) );
  drp_1 r_ic_fs_spklen_reg_6_ ( .ip(n1415), .ck(pclk), .rb(presetn), .q(
        ic_fs_spklen[6]) );
  drp_1 r_ic_fs_spklen_reg_5_ ( .ip(n1414), .ck(pclk), .rb(presetn), .q(
        ic_fs_spklen[5]) );
  drp_1 r_ic_fs_spklen_reg_4_ ( .ip(n1413), .ck(pclk), .rb(presetn), .q(
        ic_fs_spklen[4]) );
  drp_1 r_ic_fs_spklen_reg_3_ ( .ip(n1412), .ck(pclk), .rb(presetn), .q(
        ic_fs_spklen[3]) );
  drp_1 r_ic_fs_spklen_reg_1_ ( .ip(n1410), .ck(pclk), .rb(presetn), .q(
        ic_fs_spklen[1]) );
  drp_1 r_ic_hs_spklen_reg_7_ ( .ip(n1408), .ck(pclk), .rb(presetn), .q(
        ic_hs_spklen[7]) );
  drp_1 r_ic_hs_spklen_reg_6_ ( .ip(n1407), .ck(pclk), .rb(presetn), .q(
        ic_hs_spklen[6]) );
  drp_1 r_ic_hs_spklen_reg_5_ ( .ip(n1406), .ck(pclk), .rb(presetn), .q(
        ic_hs_spklen[5]) );
  drp_1 r_ic_hs_spklen_reg_4_ ( .ip(n1405), .ck(pclk), .rb(presetn), .q(
        ic_hs_spklen[4]) );
  drp_1 r_ic_hs_spklen_reg_3_ ( .ip(n1404), .ck(pclk), .rb(presetn), .q(
        ic_hs_spklen[3]) );
  drp_1 r_ic_hs_spklen_reg_2_ ( .ip(n1403), .ck(pclk), .rb(presetn), .q(
        ic_hs_spklen[2]) );
  drp_1 r_ic_hs_spklen_reg_1_ ( .ip(n1402), .ck(pclk), .rb(presetn), .q(
        ic_hs_spklen[1]) );
  drp_1 ic_intr_mask_reg_10_ ( .ip(n1398), .ck(pclk), .rb(presetn), .q(
        ic_intr_mask[10]) );
  drp_1 ic_intr_mask_reg_9_ ( .ip(n1399), .ck(pclk), .rb(presetn), .q(
        ic_intr_mask[9]) );
  drp_1 ic_intr_mask_reg_8_ ( .ip(n1400), .ck(pclk), .rb(presetn), .q(
        ic_intr_mask[8]) );
  drp_1 ic_sda_hold_reg_23_ ( .ip(n1388), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[23]) );
  drp_1 ic_sda_hold_reg_22_ ( .ip(n1387), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[22]) );
  drp_1 ic_sda_hold_reg_21_ ( .ip(n1386), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[21]) );
  drp_1 ic_sda_hold_reg_20_ ( .ip(n1385), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[20]) );
  drp_1 ic_sda_hold_reg_19_ ( .ip(n1384), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[19]) );
  drp_1 ic_sda_hold_reg_18_ ( .ip(n1383), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[18]) );
  drp_1 ic_sda_hold_reg_17_ ( .ip(n1382), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[17]) );
  drp_1 ic_sda_hold_reg_16_ ( .ip(n1381), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[16]) );
  drp_1 ic_sda_hold_reg_15_ ( .ip(n1380), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[15]) );
  drp_1 ic_sda_hold_reg_14_ ( .ip(n1379), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[14]) );
  drp_1 ic_sda_hold_reg_13_ ( .ip(n1378), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[13]) );
  drp_1 ic_sda_hold_reg_12_ ( .ip(n1377), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[12]) );
  drp_1 ic_sda_hold_reg_11_ ( .ip(n1376), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[11]) );
  drp_1 ic_sda_hold_reg_10_ ( .ip(n1375), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[10]) );
  drp_1 ic_sda_hold_reg_9_ ( .ip(n1374), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[9]) );
  drp_1 ic_sda_hold_reg_8_ ( .ip(n1373), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[8]) );
  drp_1 ic_sda_hold_reg_7_ ( .ip(n1372), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[7]) );
  drp_1 ic_sda_hold_reg_6_ ( .ip(n1371), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[6]) );
  drp_1 ic_sda_hold_reg_5_ ( .ip(n1370), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[5]) );
  drp_1 ic_sda_hold_reg_4_ ( .ip(n1369), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[4]) );
  drp_1 ic_sda_hold_reg_3_ ( .ip(n1368), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[3]) );
  drp_1 ic_sda_hold_reg_2_ ( .ip(n1367), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[2]) );
  drp_1 ic_sda_hold_reg_1_ ( .ip(n1366), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[1]) );
  drp_1 fifo_rst_n_int_reg ( .ip(fix_c), .ck(pclk), .rb(presetn), .q(
        fifo_rst_n_int) );
  drp_1 ic_txflr_reg_2_ ( .ip(n1361), .ck(pclk), .rb(presetn), .q(ic_txflr[2])
         );
  drp_1 ic_txflr_reg_3_ ( .ip(n1364), .ck(pclk), .rb(presetn), .q(ic_txflr[3])
         );
  drp_1 ic_txflr_reg_0_ ( .ip(n1363), .ck(pclk), .rb(presetn), .q(ic_txflr[0])
         );
  drp_1 ic_txflr_reg_1_ ( .ip(n1362), .ck(pclk), .rb(presetn), .q(ic_txflr[1])
         );
  drp_1 ic_hs_maddr_reg_2_ ( .ip(n1167), .ck(pclk), .rb(presetn), .q(
        ic_hs_maddr[2]) );
  drp_1 ic_hs_maddr_reg_1_ ( .ip(n1165), .ck(pclk), .rb(presetn), .q(
        ic_hs_maddr[1]) );
  drp_1 ic_rx_tl_reg_2_ ( .ip(n1153), .ck(pclk), .rb(presetn), .q(
        ic_rx_tl_int[2]) );
  drp_1 ic_rx_tl_reg_1_ ( .ip(n1151), .ck(pclk), .rb(presetn), .q(
        ic_rx_tl_int[1]) );
  drp_1 ic_rx_tl_reg_0_ ( .ip(n1149), .ck(pclk), .rb(presetn), .q(
        ic_rx_tl_int[0]) );
  drp_1 ic_tx_tl_reg_2_ ( .ip(n1137), .ck(pclk), .rb(presetn), .q(ic_tx_tl_2_)
         );
  drp_1 ic_tx_tl_reg_1_ ( .ip(n1135), .ck(pclk), .rb(presetn), .q(ic_tx_tl_1_)
         );
  drp_1 ic_tx_tl_reg_0_ ( .ip(n1133), .ck(pclk), .rb(presetn), .q(ic_tx_tl_0_)
         );
  drp_1 ic_sda_setup_reg_7_ ( .ip(n1131), .ck(pclk), .rb(presetn), .q(
        ic_sda_setup[7]) );
  drp_1 ic_sda_setup_reg_4_ ( .ip(n1129), .ck(pclk), .rb(presetn), .q(
        ic_sda_setup[4]) );
  drp_1 ic_sda_setup_reg_3_ ( .ip(n1127), .ck(pclk), .rb(presetn), .q(
        ic_sda_setup[3]) );
  drp_1 ic_sda_setup_reg_1_ ( .ip(n1125), .ck(pclk), .rb(presetn), .q(
        ic_sda_setup[1]) );
  drp_1 ic_sda_setup_reg_0_ ( .ip(n1123), .ck(pclk), .rb(presetn), .q(
        ic_sda_setup[0]) );
  drp_1 ic_txflr_flushed_reg_0_ ( .ip(n1121), .ck(pclk), .rb(presetn), .q(
        ic_txflr_flushed[0]) );
  drp_1 ic_txflr_flushed_reg_1_ ( .ip(n1119), .ck(pclk), .rb(presetn), .q(
        ic_txflr_flushed[1]) );
  drp_1 ic_txflr_flushed_reg_3_ ( .ip(n1117), .ck(pclk), .rb(presetn), .q(
        ic_txflr_flushed[3]) );
  drp_1 ic_txflr_flushed_reg_2_ ( .ip(n1115), .ck(pclk), .rb(presetn), .q(
        ic_txflr_flushed[2]) );
  drsp_1 ic_ack_general_call_reg ( .ip(n1105), .ck(pclk), .rb(1'b1), .s(n760), 
        .q(ic_ack_general_call) );
  drsp_1 ic_intr_mask_reg_11_ ( .ip(n1397), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_intr_mask[11]) );
  drsp_1 ic_intr_mask_reg_6_ ( .ip(n1390), .ck(pclk), .rb(1'b1), .s(n1), .q(
        ic_intr_mask[6]) );
  drsp_1 ic_intr_mask_reg_3_ ( .ip(n1393), .ck(pclk), .rb(1'b1), .s(n485), .q(
        ic_intr_mask[3]) );
  drsp_1 ic_intr_mask_reg_7_ ( .ip(n1389), .ck(pclk), .rb(1'b1), .s(n760), .q(
        ic_intr_mask[7]) );
  drsp_1 ic_intr_mask_reg_4_ ( .ip(n1392), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_intr_mask[4]) );
  drsp_1 ic_intr_mask_reg_1_ ( .ip(n1395), .ck(pclk), .rb(1'b1), .s(n1), .q(
        ic_intr_mask[1]) );
  drsp_1 ic_intr_mask_reg_5_ ( .ip(n1391), .ck(pclk), .rb(1'b1), .s(n485), .q(
        ic_intr_mask[5]) );
  drsp_1 ic_intr_mask_reg_2_ ( .ip(n1394), .ck(pclk), .rb(1'b1), .s(n760), .q(
        ic_intr_mask[2]) );
  drsp_1 ic_intr_mask_reg_0_ ( .ip(n1396), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_intr_mask[0]) );
  drsp_1 ic_hs_maddr_reg_0_ ( .ip(n1113), .ck(pclk), .rb(1'b1), .s(n1), .q(
        ic_hs_maddr[0]) );
  drsp_1 r_ic_hs_spklen_reg_0_ ( .ip(n1401), .ck(pclk), .rb(1'b1), .s(n485), 
        .q(ic_hs_spklen[0]) );
  drsp_1 r_ic_fs_spklen_reg_0_ ( .ip(n1409), .ck(pclk), .rb(1'b1), .s(n760), 
        .q(ic_fs_spklen[0]) );
  drsp_1 r_ic_fs_spklen_reg_2_ ( .ip(n1411), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_fs_spklen[2]) );
  drsp_1 ic_sda_setup_reg_6_ ( .ip(n1111), .ck(pclk), .rb(1'b1), .s(n1), .q(
        ic_sda_setup[6]) );
  drsp_1 ic_sda_setup_reg_5_ ( .ip(n1109), .ck(pclk), .rb(1'b1), .s(n485), .q(
        ic_sda_setup[5]) );
  drsp_1 ic_sda_setup_reg_2_ ( .ip(n1107), .ck(pclk), .rb(1'b1), .s(n760), .q(
        ic_sda_setup[2]) );
  drsp_1 ic_sar_reg_6_ ( .ip(n1522), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_sar[6]) );
  drsp_1 ic_sar_reg_4_ ( .ip(n1524), .ck(pclk), .rb(1'b1), .s(n1), .q(
        ic_sar[4]) );
  drsp_1 ic_sar_reg_2_ ( .ip(n1526), .ck(pclk), .rb(1'b1), .s(n485), .q(
        ic_sar[2]) );
  drsp_1 ic_sar_reg_0_ ( .ip(n1528), .ck(pclk), .rb(1'b1), .s(n760), .q(
        ic_sar[0]) );
  drsp_1 ic_con_pre_reg_2_ ( .ip(n1537), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_con_pre_2_) );
  drsp_1 ic_con_pre_reg_1_ ( .ip(n1536), .ck(pclk), .rb(1'b1), .s(n1), .q(
        ic_con_pre_1_) );
  drsp_1 ic_con_pre_reg_6_ ( .ip(n1541), .ck(pclk), .rb(1'b1), .s(n485), .q(
        ic_con_pre_6_) );
  drsp_1 ic_con_pre_reg_3_ ( .ip(n1538), .ck(pclk), .rb(1'b1), .s(n760), .q(
        ic_10bit_slv) );
  drsp_1 ic_con_pre_reg_4_ ( .ip(n1539), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_10bit_mst) );
  drsp_1 ic_con_pre_reg_5_ ( .ip(n1540), .ck(pclk), .rb(1'b1), .s(n1), .q(
        ic_rstrt_en) );
  drsp_1 ic_con_pre_reg_0_ ( .ip(n1535), .ck(pclk), .rb(1'b1), .s(n485), .q(
        ic_master) );
  drsp_1 ic_tar_reg_reg_6_ ( .ip(n1514), .ck(pclk), .rb(1'b1), .s(n760), .q(
        ic_tar[6]) );
  drsp_1 ic_tar_reg_reg_4_ ( .ip(n1516), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_tar[4]) );
  drsp_1 ic_tar_reg_reg_2_ ( .ip(n1518), .ck(pclk), .rb(1'b1), .s(n1), .q(
        ic_tar[2]) );
  drsp_1 ic_tar_reg_reg_0_ ( .ip(n1520), .ck(pclk), .rb(1'b1), .s(n485), .q(
        ic_tar[0]) );
  drsp_1 ic_sda_hold_reg_0_ ( .ip(n1365), .ck(pclk), .rb(1'b1), .s(n760), .q(
        ic_sda_hold[0]) );
  drsp_1 r_ic_hs_hcnt_reg_2_ ( .ip(n1446), .ck(pclk), .rb(1'b1), .s(n2), .q(
        hcr_ic_hs_hcnt[2]) );
  drsp_1 r_ic_hs_hcnt_reg_1_ ( .ip(n1447), .ck(pclk), .rb(1'b1), .s(n1), .q(
        hcr_ic_hs_hcnt[1]) );
  drsp_1 r_ic_fs_hcnt_reg_2_ ( .ip(n1478), .ck(pclk), .rb(1'b1), .s(n485), .q(
        ic_fs_hcnt[2]) );
  drsp_1 r_ic_fs_hcnt_reg_5_ ( .ip(n1475), .ck(pclk), .rb(1'b1), .s(n760), .q(
        ic_fs_hcnt[5]) );
  drsp_1 r_ic_fs_lcnt_reg_7_ ( .ip(n1457), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_fs_lcnt[7]) );
  drsp_1 r_ic_ss_lcnt_reg_2_ ( .ip(n1494), .ck(pclk), .rb(1'b1), .s(n1), .q(
        hcr_ic_ss_lcnt[2]) );
  drsp_1 r_ic_ss_lcnt_reg_1_ ( .ip(n1495), .ck(pclk), .rb(1'b1), .s(n485), .q(
        hcr_ic_ss_lcnt[1]) );
  drsp_1 r_ic_ss_lcnt_reg_8_ ( .ip(n1487), .ck(pclk), .rb(1'b1), .s(n760), .q(
        hcr_ic_ss_lcnt[8]) );
  drsp_1 r_ic_ss_lcnt_reg_6_ ( .ip(n1490), .ck(pclk), .rb(1'b1), .s(n2), .q(
        hcr_ic_ss_lcnt[6]) );
  drsp_1 r_ic_ss_lcnt_reg_7_ ( .ip(n1489), .ck(pclk), .rb(1'b1), .s(n1), .q(
        hcr_ic_ss_lcnt[7]) );
  drsp_1 r_ic_ss_lcnt_reg_4_ ( .ip(n1492), .ck(pclk), .rb(1'b1), .s(n485), .q(
        hcr_ic_ss_lcnt[4]) );
  drsp_1 r_ic_hs_lcnt_reg_4_ ( .ip(n1428), .ck(pclk), .rb(1'b1), .s(n760), .q(
        hcr_ic_hs_lcnt[4]) );
  drsp_1 r_ic_fs_lcnt_reg_1_ ( .ip(n1463), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_fs_lcnt[1]) );
  drsp_1 r_ic_ss_hcnt_reg_8_ ( .ip(n1503), .ck(pclk), .rb(1'b1), .s(n1), .q(
        hcr_ic_ss_hcnt[8]) );
  drsp_1 r_ic_ss_hcnt_reg_7_ ( .ip(n1505), .ck(pclk), .rb(1'b1), .s(n485), .q(
        hcr_ic_ss_hcnt[7]) );
  drsp_1 r_ic_ss_hcnt_reg_4_ ( .ip(n1508), .ck(pclk), .rb(1'b1), .s(n760), .q(
        hcr_ic_ss_hcnt[4]) );
  drsp_1 r_ic_fs_hcnt_reg_3_ ( .ip(n1477), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_fs_hcnt[3]) );
  drsp_1 r_ic_fs_hcnt_reg_4_ ( .ip(n1476), .ck(pclk), .rb(1'b1), .s(n1), .q(
        ic_fs_hcnt[4]) );
  nor2_1 U3 ( .ip1(n35), .ip2(n208), .op(n668) );
  nand3_1 U4 ( .ip1(n515), .ip2(n514), .ip3(n513), .op(ic_hcnt[8]) );
  nand3_1 U5 ( .ip1(n503), .ip2(n502), .ip3(n501), .op(ic_hcnt[5]) );
  nand3_1 U6 ( .ip1(n500), .ip2(n499), .ip3(n498), .op(ic_hcnt[4]) );
  nand3_1 U7 ( .ip1(n509), .ip2(n508), .ip3(n507), .op(ic_hcnt[7]) );
  nand3_1 U8 ( .ip1(n530), .ip2(n529), .ip3(n528), .op(ic_hcnt[11]) );
  nand3_1 U9 ( .ip1(n512), .ip2(n511), .ip3(n510), .op(ic_hcnt[14]) );
  nand3_1 U10 ( .ip1(n518), .ip2(n517), .ip3(n516), .op(ic_hcnt[10]) );
  nand3_1 U11 ( .ip1(n506), .ip2(n505), .ip3(n504), .op(ic_hcnt[6]) );
  nand3_1 U12 ( .ip1(n527), .ip2(n526), .ip3(n525), .op(ic_hcnt[12]) );
  nand3_1 U13 ( .ip1(n524), .ip2(n523), .ip3(n522), .op(ic_hcnt[13]) );
  nand3_1 U14 ( .ip1(n478), .ip2(n477), .ip3(n476), .op(ic_hcnt[15]) );
  nand3_1 U15 ( .ip1(n597), .ip2(n22), .ip3(n21), .op(n602) );
  inv_1 U16 ( .ip(n13), .op(n614) );
  nand2_1 U17 ( .ip1(n23), .ip2(n50), .op(n35) );
  inv_1 U18 ( .ip(fifo_rst_n), .op(n112) );
  nand2_1 U19 ( .ip1(fifo_rst_n), .ip2(n474), .op(n473) );
  nand3_1 U20 ( .ip1(n536), .ip2(n535), .ip3(n534), .op(ic_lcnt[1]) );
  nand3_1 U21 ( .ip1(n491), .ip2(n490), .ip3(n489), .op(ic_hcnt[1]) );
  nand3_1 U22 ( .ip1(n542), .ip2(n541), .ip3(n540), .op(ic_lcnt[2]) );
  nand3_1 U23 ( .ip1(n539), .ip2(n538), .ip3(n537), .op(ic_lcnt[3]) );
  nand3_1 U24 ( .ip1(n545), .ip2(n544), .ip3(n543), .op(ic_lcnt[5]) );
  nand3_1 U25 ( .ip1(n533), .ip2(n532), .ip3(n531), .op(ic_lcnt[0]) );
  nand3_1 U26 ( .ip1(n497), .ip2(n496), .ip3(n495), .op(ic_hcnt[3]) );
  nand3_1 U27 ( .ip1(n494), .ip2(n493), .ip3(n492), .op(ic_hcnt[2]) );
  nand3_1 U28 ( .ip1(n569), .ip2(n568), .ip3(n567), .op(ic_lcnt[9]) );
  nand3_1 U29 ( .ip1(n548), .ip2(n547), .ip3(n546), .op(ic_lcnt[4]) );
  nand3_1 U30 ( .ip1(n554), .ip2(n553), .ip3(n552), .op(ic_lcnt[6]) );
  nand3_1 U31 ( .ip1(n551), .ip2(n550), .ip3(n549), .op(ic_lcnt[7]) );
  nand3_1 U32 ( .ip1(n566), .ip2(n565), .ip3(n564), .op(ic_lcnt[10]) );
  nand3_1 U33 ( .ip1(n573), .ip2(n572), .ip3(n571), .op(ic_lcnt[8]) );
  nand3_1 U34 ( .ip1(n560), .ip2(n559), .ip3(n558), .op(ic_lcnt[12]) );
  nand3_1 U35 ( .ip1(n563), .ip2(n562), .ip3(n561), .op(ic_lcnt[11]) );
  nand3_1 U36 ( .ip1(n521), .ip2(n520), .ip3(n519), .op(ic_hcnt[9]) );
  nand3_1 U37 ( .ip1(n557), .ip2(n556), .ip3(n555), .op(ic_lcnt[13]) );
  nand3_1 U38 ( .ip1(n481), .ip2(n480), .ip3(n479), .op(ic_lcnt[14]) );
  nand3_1 U39 ( .ip1(n484), .ip2(n483), .ip3(n482), .op(ic_lcnt[15]) );
  nor2_1 U40 ( .ip1(n57), .ip2(n47), .op(n650) );
  inv_1 U41 ( .ip(n602), .op(n590) );
  nand2_1 U42 ( .ip1(n118), .ip2(n117), .op(n161) );
  nor2_1 U43 ( .ip1(n242), .ip2(n241), .op(n86) );
  nand2_1 U44 ( .ip1(n42), .ip2(n50), .op(n110) );
  inv_1 U45 ( .ip(n23), .op(n43) );
  inv_1 U46 ( .ip(n42), .op(n49) );
  nor2_1 U47 ( .ip1(n242), .ip2(n208), .op(n632) );
  nand3_1 U48 ( .ip1(n33), .ip2(n34), .ip3(n32), .op(n58) );
  nor2_1 U49 ( .ip1(n43), .ip2(n48), .op(n651) );
  nor2_1 U50 ( .ip1(n242), .ip2(n58), .op(n619) );
  nor2_1 U51 ( .ip1(n65), .ip2(n208), .op(n633) );
  nor2_1 U52 ( .ip1(n49), .ip2(n48), .op(n649) );
  nor2_1 U53 ( .ip1(n111), .ip2(n110), .op(ic_clr_tx_abrt_en) );
  nor2_1 U54 ( .ip1(n35), .ip2(n4), .op(ic_clr_intr_en) );
  nand2_1 U55 ( .ip1(n660), .ip2(n625), .op(n628) );
  nand2_1 U56 ( .ip1(n619), .ip2(n625), .op(n623) );
  nand2_1 U57 ( .ip1(n442), .ip2(n689), .op(n606) );
  nor2_1 U58 ( .ip1(n441), .ip2(n606), .op(n607) );
  inv_1 U59 ( .ip(n610), .op(n689) );
  nand2_1 U60 ( .ip1(n676), .ip2(n625), .op(n624) );
  nand2_1 U61 ( .ip1(n650), .ip2(n625), .op(n627) );
  nand2_1 U62 ( .ip1(n659), .ip2(n625), .op(n630) );
  nor2_1 U63 ( .ip1(n161), .ip2(n630), .op(n141) );
  nor2_1 U64 ( .ip1(n590), .ip2(n24), .op(n29) );
  nand2_1 U65 ( .ip1(n632), .ip2(n625), .op(n605) );
  nor2_1 U66 ( .ip1(n161), .ip2(n605), .op(n192) );
  nand2_1 U67 ( .ip1(n641), .ip2(n625), .op(n603) );
  nand2_1 U68 ( .ip1(n651), .ip2(n625), .op(n621) );
  nand2_1 U69 ( .ip1(n11), .ip2(n473), .op(n683) );
  nor2_1 U70 ( .ip1(n6), .ip2(n680), .op(n615) );
  nor2_1 U71 ( .ip1(n13), .ip2(n10), .op(n474) );
  nor2_1 U72 ( .ip1(n456), .ip2(n3), .op(fifo_rst_n) );
  nor2_1 U73 ( .ip1(n242), .ip2(n198), .op(n677) );
  nor2_1 U74 ( .ip1(n65), .ip2(n72), .op(n648) );
  nor2_1 U75 ( .ip1(n110), .ip2(n208), .op(n641) );
  nor2_1 U76 ( .ip1(n43), .ip2(n57), .op(n652) );
  nor2_1 U77 ( .ip1(n207), .ip2(n198), .op(iprdata[29]) );
  nor2_1 U78 ( .ip1(n48), .ip2(n47), .op(n678) );
  nor2_1 U79 ( .ip1(n49), .ip2(n57), .op(n659) );
  nor2_1 U80 ( .ip1(n242), .ip2(n72), .op(n658) );
  nor2_1 U81 ( .ip1(n65), .ip2(n58), .op(n669) );
  nor2_1 U82 ( .ip1(n35), .ip2(n51), .op(n661) );
  nor2_1 U83 ( .ip1(n199), .ip2(n57), .op(n676) );
  nor2_1 U84 ( .ip1(n570), .ip2(n679), .op(ic_hs) );
  inv_1 U85 ( .ip(n7), .op(rx_pop) );
  inv_1 U86 ( .ip(n440), .op(tx_push) );
  nor2_1 U87 ( .ip1(n161), .ip2(n603), .op(n144) );
  nand2_1 U88 ( .ip1(n652), .ip2(n625), .op(n24) );
  nand2_1 U89 ( .ip1(n648), .ip2(n625), .op(n589) );
  nand2_1 U90 ( .ip1(n633), .ip2(n625), .op(n591) );
  nand2_1 U91 ( .ip1(n649), .ip2(n625), .op(n622) );
  nand2_1 U92 ( .ip1(n677), .ip2(n625), .op(n596) );
  buf_1 U93 ( .ip(n596), .op(n629) );
  nand2_1 U94 ( .ip1(n669), .ip2(n625), .op(n620) );
  inv_1 U95 ( .ip(presetn), .op(n1) );
  inv_1 U96 ( .ip(presetn), .op(n2) );
  inv_1 U148 ( .ip(ic_enable[0]), .op(n706) );
  inv_1 U149 ( .ip(fifo_rst_n_int), .op(n113) );
  nor3_4 U150 ( .ip1(slv_clr_leftover_flg_edg), .ip2(n706), .ip3(n113), .op(
        tx_fifo_rst_n) );
  inv_1 U151 ( .ip(reg_addr[3]), .op(n33) );
  nand3_1 U152 ( .ip1(reg_addr[4]), .ip2(reg_addr[2]), .ip3(n33), .op(n111) );
  nor2_1 U153 ( .ip1(reg_addr[0]), .ip2(reg_addr[5]), .op(n23) );
  inv_1 U154 ( .ip(reg_addr[1]), .op(n50) );
  nor2_1 U155 ( .ip1(n111), .ip2(n35), .op(ic_clr_rd_req_en) );
  inv_1 U156 ( .ip(reg_addr[2]), .op(n32) );
  nand3_1 U157 ( .ip1(reg_addr[4]), .ip2(reg_addr[3]), .ip3(n32), .op(n241) );
  nor2_1 U158 ( .ip1(n35), .ip2(n241), .op(ic_clr_stop_det_en) );
  inv_1 U159 ( .ip(reg_addr[0]), .op(n93) );
  nor2_1 U160 ( .ip1(reg_addr[5]), .ip2(n93), .op(n42) );
  nand2_1 U161 ( .ip1(reg_addr[1]), .ip2(n42), .op(n242) );
  nand2_1 U162 ( .ip1(n86), .ip2(wr_en), .op(n583) );
  nor2_1 U163 ( .ip1(ipwdata[0]), .ip2(n583), .op(n456) );
  inv_1 U164 ( .ip(tx_abrt_flg_edg), .op(n584) );
  nand2_1 U165 ( .ip1(n584), .ip2(ic_enable[0]), .op(n3) );
  nand2_1 U166 ( .ip1(reg_addr[0]), .ip2(reg_addr[5]), .op(n199) );
  nand3_1 U167 ( .ip1(reg_addr[3]), .ip2(reg_addr[4]), .ip3(reg_addr[2]), .op(
        n198) );
  nor3_1 U168 ( .ip1(n50), .ip2(n199), .ip3(n198), .op(iprdata[30]) );
  nand3_1 U169 ( .ip1(reg_addr[4]), .ip2(n33), .ip3(n32), .op(n4) );
  nand2_1 U170 ( .ip1(reg_addr[1]), .ip2(n23), .op(n65) );
  nor2_1 U171 ( .ip1(n65), .ip2(n4), .op(ic_clr_rx_over_en) );
  nor2_1 U172 ( .ip1(n242), .ip2(n4), .op(ic_clr_tx_over_en) );
  nor2_1 U173 ( .ip1(n65), .ip2(n241), .op(ic_clr_gen_call_en) );
  nor2_1 U174 ( .ip1(n242), .ip2(n111), .op(ic_clr_activity_en) );
  nor2_1 U175 ( .ip1(n111), .ip2(n65), .op(ic_clr_rx_done_en) );
  nor2_1 U176 ( .ip1(n110), .ip2(n4), .op(ic_clr_rx_under_en) );
  nor2_1 U177 ( .ip1(n110), .ip2(n241), .op(ic_clr_start_det_en) );
  inv_1 U178 ( .ip(ic_rxflr[1]), .op(n6) );
  inv_1 U179 ( .ip(rx_push_sync), .op(n5) );
  inv_1 U180 ( .ip(reg_addr[4]), .op(n34) );
  nand3_1 U181 ( .ip1(reg_addr[2]), .ip2(n33), .ip3(n34), .op(n208) );
  nand2_1 U182 ( .ip1(n668), .ip2(rd_en), .op(n7) );
  nor4_1 U183 ( .ip1(n112), .ip2(n5), .ip3(ic_rxflr[3]), .ip4(rx_pop), .op(n10) );
  nand2_1 U184 ( .ip1(ic_rxflr[0]), .ip2(n10), .op(n680) );
  nand2_1 U185 ( .ip1(ic_rxflr[2]), .ip2(n615), .op(n17) );
  nor4_1 U186 ( .ip1(ic_rxflr[0]), .ip2(ic_rxflr[3]), .ip3(ic_rxflr[1]), .ip4(
        ic_rxflr[2]), .op(n8) );
  nor4_1 U187 ( .ip1(rx_push_sync), .ip2(n8), .ip3(n112), .ip4(n7), .op(n13)
         );
  inv_1 U188 ( .ip(n10), .op(n9) );
  nor2_1 U189 ( .ip1(n9), .ip2(ic_rxflr[1]), .op(n12) );
  mux2_1 U190 ( .ip1(n9), .ip2(n614), .s(ic_rxflr[0]), .op(n11) );
  not_ab_or_c_or_d U191 ( .ip1(ic_rxflr[1]), .ip2(n13), .ip3(n12), .ip4(n683), 
        .op(n616) );
  nand2_1 U192 ( .ip1(ic_rxflr[2]), .ip2(n13), .op(n14) );
  nand2_1 U193 ( .ip1(n616), .ip2(n14), .op(n15) );
  nand2_1 U194 ( .ip1(ic_rxflr[3]), .ip2(n15), .op(n16) );
  nand2_1 U195 ( .ip1(n17), .ip2(n16), .op(n1547) );
  inv_1 U196 ( .ip(ipwdata[5]), .op(n19) );
  inv_1 U197 ( .ip(ipwdata[6]), .op(n18) );
  nand2_1 U198 ( .ip1(n19), .ip2(n18), .op(n20) );
  nor4_1 U199 ( .ip1(ipwdata[3]), .ip2(ipwdata[4]), .ip3(ipwdata[7]), .ip4(n20), .op(n597) );
  nor4_1 U200 ( .ip1(ipwdata[8]), .ip2(ipwdata[9]), .ip3(ipwdata[10]), .ip4(
        ipwdata[11]), .op(n22) );
  nor4_1 U201 ( .ip1(ipwdata[14]), .ip2(ipwdata[12]), .ip3(ipwdata[13]), .ip4(
        ipwdata[15]), .op(n21) );
  nand3_1 U202 ( .ip1(n34), .ip2(n32), .ip3(reg_addr[3]), .op(n72) );
  or2_1 U203 ( .ip1(n72), .ip2(reg_addr[1]), .op(n57) );
  and2_1 U204 ( .ip1(n706), .ip2(wr_en), .op(n625) );
  nand2_1 U205 ( .ip1(ipwdata[0]), .ip2(n29), .op(n26) );
  nand2_1 U206 ( .ip1(ic_fs_lcnt[0]), .ip2(n24), .op(n25) );
  nand2_1 U207 ( .ip1(n26), .ip2(n25), .op(n1464) );
  nand2_1 U208 ( .ip1(n29), .ip2(ipwdata[1]), .op(n28) );
  nand2_1 U209 ( .ip1(ic_fs_lcnt[1]), .ip2(n24), .op(n27) );
  nand2_1 U210 ( .ip1(n28), .ip2(n27), .op(n1463) );
  nand2_1 U211 ( .ip1(n29), .ip2(ipwdata[2]), .op(n31) );
  nand2_1 U212 ( .ip1(ic_fs_lcnt[2]), .ip2(n24), .op(n30) );
  nand2_1 U213 ( .ip1(n31), .ip2(n30), .op(n1462) );
  nand3_1 U214 ( .ip1(reg_addr[3]), .ip2(reg_addr[2]), .ip3(n34), .op(n51) );
  and2_1 U215 ( .ip1(n661), .ip2(ic_intr_mask[2]), .op(n41) );
  nand2_1 U216 ( .ip1(n668), .ip2(rx_pop_data[2]), .op(n39) );
  nor2_1 U217 ( .ip1(n110), .ip2(n51), .op(n638) );
  nand2_1 U218 ( .ip1(n638), .ip2(ic_raw_intr_stat[2]), .op(n38) );
  nor2_1 U219 ( .ip1(n65), .ip2(n198), .op(n639) );
  nand2_1 U220 ( .ip1(n639), .ip2(ic_rxflr[2]), .op(n37) );
  nor2_1 U221 ( .ip1(n35), .ip2(n198), .op(n404) );
  nand2_1 U222 ( .ip1(n404), .ip2(tx_empty), .op(n36) );
  nand4_1 U223 ( .ip1(n39), .ip2(n38), .ip3(n37), .ip4(n36), .op(n40) );
  not_ab_or_c_or_d U224 ( .ip1(n669), .ip2(ic_sar[2]), .ip3(n41), .ip4(n40), 
        .op(n76) );
  or2_1 U225 ( .ip1(n58), .ip2(reg_addr[1]), .op(n48) );
  nand2_1 U226 ( .ip1(reg_addr[5]), .ip2(n93), .op(n47) );
  nand2_1 U227 ( .ip1(n650), .ip2(ic_fs_spklen[2]), .op(n46) );
  nand2_1 U228 ( .ip1(n651), .ip2(ic_con_pre_2_), .op(n45) );
  nand2_1 U229 ( .ip1(n652), .ip2(ic_fs_lcnt[2]), .op(n44) );
  nand3_1 U230 ( .ip1(n46), .ip2(n45), .ip3(n44), .op(n71) );
  nor2_1 U231 ( .ip1(n65), .ip2(n51), .op(n578) );
  nor3_1 U232 ( .ip1(reg_addr[1]), .ip2(n199), .ip3(n198), .op(n657) );
  nand2_1 U233 ( .ip1(n678), .ip2(ic_tx_abrt_source[2]), .op(n55) );
  nand2_1 U234 ( .ip1(n659), .ip2(hcr_ic_hs_hcnt[2]), .op(n54) );
  nor3_1 U235 ( .ip1(n50), .ip2(n199), .ip3(n208), .op(n245) );
  nand2_1 U236 ( .ip1(n245), .ip2(slv_fifo_filled_and_flushed_sync), .op(n53)
         );
  nor2_1 U237 ( .ip1(n242), .ip2(n51), .op(n576) );
  nand2_1 U238 ( .ip1(n576), .ip2(ic_tx_tl_2_), .op(n52) );
  nand4_1 U239 ( .ip1(n55), .ip2(n54), .ip3(n53), .ip4(n52), .op(n56) );
  not_ab_or_c_or_d U240 ( .ip1(n578), .ip2(ic_rx_tl_int[2]), .ip3(n657), .ip4(
        n56), .op(n69) );
  and2_1 U241 ( .ip1(n632), .ip2(ic_fs_hcnt[2]), .op(n64) );
  nand2_1 U242 ( .ip1(n633), .ip2(hcr_ic_ss_lcnt[2]), .op(n62) );
  nand2_1 U243 ( .ip1(n677), .ip2(ic_sda_hold[2]), .op(n61) );
  nand2_1 U244 ( .ip1(n676), .ip2(ic_hs_spklen[2]), .op(n60) );
  nand2_1 U245 ( .ip1(n619), .ip2(ic_hs_maddr[2]), .op(n59) );
  nand4_1 U246 ( .ip1(n62), .ip2(n61), .ip3(n60), .ip4(n59), .op(n63) );
  not_ab_or_c_or_d U247 ( .ip1(hcr_ic_ss_hcnt[2]), .ip2(n641), .ip3(n64), 
        .ip4(n63), .op(n68) );
  nand2_1 U248 ( .ip1(n648), .ip2(hcr_ic_hs_lcnt[2]), .op(n67) );
  nor2_1 U249 ( .ip1(n110), .ip2(n198), .op(n640) );
  nand2_1 U250 ( .ip1(n640), .ip2(ic_txflr[2]), .op(n66) );
  nand4_1 U251 ( .ip1(n69), .ip2(n68), .ip3(n67), .ip4(n66), .op(n70) );
  not_ab_or_c_or_d U252 ( .ip1(n649), .ip2(ic_tar[2]), .ip3(n71), .ip4(n70), 
        .op(n75) );
  nor3_1 U253 ( .ip1(reg_addr[1]), .ip2(n199), .ip3(n208), .op(n660) );
  nand2_1 U254 ( .ip1(n660), .ip2(ic_sda_setup[2]), .op(n74) );
  nand2_1 U255 ( .ip1(n658), .ip2(ic_intr_stat[2]), .op(n73) );
  nand4_1 U256 ( .ip1(n76), .ip2(n75), .ip3(n74), .ip4(n73), .op(iprdata[2])
         );
  inv_1 U257 ( .ip(n404), .op(n637) );
  nor2_1 U258 ( .ip1(tx_full), .ip2(n637), .op(n82) );
  nand2_1 U259 ( .ip1(n668), .ip2(rx_pop_data[1]), .op(n80) );
  nand2_1 U260 ( .ip1(ic_raw_intr_stat[1]), .ip2(n638), .op(n79) );
  nand2_1 U261 ( .ip1(n640), .ip2(ic_txflr[1]), .op(n78) );
  nand2_1 U262 ( .ip1(n648), .ip2(hcr_ic_hs_lcnt[1]), .op(n77) );
  nand4_1 U263 ( .ip1(n80), .ip2(n79), .ip3(n78), .ip4(n77), .op(n81) );
  not_ab_or_c_or_d U264 ( .ip1(ic_rxflr[1]), .ip2(n639), .ip3(n82), .ip4(n81), 
        .op(n109) );
  nand2_1 U265 ( .ip1(n651), .ip2(ic_con_pre_1_), .op(n85) );
  nand2_1 U266 ( .ip1(n652), .ip2(ic_fs_lcnt[1]), .op(n84) );
  nand2_1 U267 ( .ip1(n678), .ip2(ic_tx_abrt_source[1]), .op(n83) );
  nand3_1 U268 ( .ip1(n85), .ip2(n84), .ip3(n83), .op(n105) );
  and2_1 U269 ( .ip1(n576), .ip2(ic_tx_tl_1_), .op(n92) );
  nand2_1 U270 ( .ip1(n578), .ip2(ic_rx_tl_int[1]), .op(n90) );
  nand2_1 U271 ( .ip1(n86), .ip2(ic_enable[1]), .op(n89) );
  nand2_1 U272 ( .ip1(n658), .ip2(ic_intr_stat[1]), .op(n88) );
  nand2_1 U273 ( .ip1(n660), .ip2(ic_sda_setup[1]), .op(n87) );
  nand4_1 U274 ( .ip1(n90), .ip2(n89), .ip3(n88), .ip4(n87), .op(n91) );
  not_ab_or_c_or_d U275 ( .ip1(slv_rx_aborted_sync), .ip2(n245), .ip3(n92), 
        .ip4(n91), .op(n103) );
  nand3_1 U276 ( .ip1(reg_addr[1]), .ip2(reg_addr[5]), .ip3(n93), .op(n207) );
  not_ab_or_c_or_d U277 ( .ip1(n619), .ip2(ic_hs_maddr[1]), .ip3(iprdata[29]), 
        .ip4(n657), .op(n102) );
  and2_1 U278 ( .ip1(n632), .ip2(ic_fs_hcnt[1]), .op(n99) );
  nand2_1 U279 ( .ip1(n633), .ip2(hcr_ic_ss_lcnt[1]), .op(n97) );
  nand2_1 U280 ( .ip1(n677), .ip2(ic_sda_hold[1]), .op(n96) );
  nand2_1 U281 ( .ip1(n676), .ip2(ic_hs_spklen[1]), .op(n95) );
  nand2_1 U282 ( .ip1(n650), .ip2(ic_fs_spklen[1]), .op(n94) );
  nand4_1 U283 ( .ip1(n97), .ip2(n96), .ip3(n95), .ip4(n94), .op(n98) );
  not_ab_or_c_or_d U284 ( .ip1(hcr_ic_ss_hcnt[1]), .ip2(n641), .ip3(n99), 
        .ip4(n98), .op(n101) );
  nand2_1 U285 ( .ip1(n659), .ip2(hcr_ic_hs_hcnt[1]), .op(n100) );
  nand4_1 U286 ( .ip1(n103), .ip2(n102), .ip3(n101), .ip4(n100), .op(n104) );
  not_ab_or_c_or_d U287 ( .ip1(n649), .ip2(ic_tar[1]), .ip3(n105), .ip4(n104), 
        .op(n108) );
  nand2_1 U288 ( .ip1(n661), .ip2(ic_intr_mask[1]), .op(n107) );
  nand2_1 U289 ( .ip1(n669), .ip2(ic_sar[1]), .op(n106) );
  nand4_1 U290 ( .ip1(n109), .ip2(n108), .ip3(n107), .ip4(n106), .op(
        iprdata[1]) );
  inv_1 U291 ( .ip(ic_clr_tx_abrt_en), .op(n238) );
  or2_1 U292 ( .ip1(n238), .ip2(n112), .op(n115) );
  or2_1 U293 ( .ip1(n113), .ip2(n112), .op(n114) );
  nand2_1 U294 ( .ip1(n115), .ip2(n114), .op(n116) );
  or2_1 U295 ( .ip1(n116), .ip2(n706), .op(fix_c) );
  or2_1 U296 ( .ip1(ipwdata[2]), .ip2(n602), .op(n118) );
  or2_1 U297 ( .ip1(ipwdata[1]), .ip2(n602), .op(n117) );
  nand2_1 U298 ( .ip1(ipwdata[15]), .ip2(n141), .op(n120) );
  nand2_1 U299 ( .ip1(hcr_ic_hs_hcnt[15]), .ip2(n630), .op(n119) );
  nand2_1 U300 ( .ip1(n120), .ip2(n119), .op(n1440) );
  nand2_1 U301 ( .ip1(ipwdata[13]), .ip2(n141), .op(n122) );
  nand2_1 U302 ( .ip1(hcr_ic_hs_hcnt[13]), .ip2(n630), .op(n121) );
  nand2_1 U303 ( .ip1(n122), .ip2(n121), .op(n1434) );
  nand2_1 U304 ( .ip1(ipwdata[12]), .ip2(n141), .op(n124) );
  nand2_1 U305 ( .ip1(hcr_ic_hs_hcnt[12]), .ip2(n630), .op(n123) );
  nand2_1 U306 ( .ip1(n124), .ip2(n123), .op(n1435) );
  nand2_1 U307 ( .ip1(ipwdata[14]), .ip2(n141), .op(n126) );
  nand2_1 U308 ( .ip1(hcr_ic_hs_hcnt[14]), .ip2(n630), .op(n125) );
  nand2_1 U309 ( .ip1(n126), .ip2(n125), .op(n1433) );
  nand2_1 U310 ( .ip1(ipwdata[11]), .ip2(n141), .op(n128) );
  nand2_1 U311 ( .ip1(hcr_ic_hs_hcnt[11]), .ip2(n630), .op(n127) );
  nand2_1 U312 ( .ip1(n128), .ip2(n127), .op(n1436) );
  nand2_1 U313 ( .ip1(ipwdata[10]), .ip2(n141), .op(n130) );
  nand2_1 U314 ( .ip1(hcr_ic_hs_hcnt[10]), .ip2(n630), .op(n129) );
  nand2_1 U315 ( .ip1(n130), .ip2(n129), .op(n1437) );
  nand2_1 U316 ( .ip1(ipwdata[9]), .ip2(n141), .op(n132) );
  nand2_1 U317 ( .ip1(hcr_ic_hs_hcnt[9]), .ip2(n630), .op(n131) );
  nand2_1 U318 ( .ip1(n132), .ip2(n131), .op(n1438) );
  nand2_1 U319 ( .ip1(ipwdata[8]), .ip2(n141), .op(n134) );
  nand2_1 U320 ( .ip1(hcr_ic_hs_hcnt[8]), .ip2(n630), .op(n133) );
  nand2_1 U321 ( .ip1(n134), .ip2(n133), .op(n1439) );
  nand2_1 U322 ( .ip1(ipwdata[7]), .ip2(n141), .op(n136) );
  nand2_1 U323 ( .ip1(hcr_ic_hs_hcnt[7]), .ip2(n630), .op(n135) );
  nand2_1 U324 ( .ip1(n136), .ip2(n135), .op(n1441) );
  nand2_1 U325 ( .ip1(ipwdata[3]), .ip2(n141), .op(n138) );
  nand2_1 U326 ( .ip1(hcr_ic_hs_hcnt[3]), .ip2(n630), .op(n137) );
  nand2_1 U327 ( .ip1(n138), .ip2(n137), .op(n1445) );
  nand2_1 U328 ( .ip1(ipwdata[4]), .ip2(n141), .op(n140) );
  nand2_1 U329 ( .ip1(hcr_ic_hs_hcnt[4]), .ip2(n630), .op(n139) );
  nand2_1 U330 ( .ip1(n140), .ip2(n139), .op(n1444) );
  nand2_1 U331 ( .ip1(ipwdata[0]), .ip2(n141), .op(n143) );
  nand2_1 U332 ( .ip1(hcr_ic_hs_hcnt[0]), .ip2(n630), .op(n142) );
  nand2_1 U333 ( .ip1(n143), .ip2(n142), .op(n1448) );
  nand2_1 U334 ( .ip1(ipwdata[12]), .ip2(n144), .op(n146) );
  nand2_1 U335 ( .ip1(hcr_ic_ss_hcnt[12]), .ip2(n603), .op(n145) );
  nand2_1 U336 ( .ip1(n146), .ip2(n145), .op(n1499) );
  nand2_1 U337 ( .ip1(ipwdata[13]), .ip2(n144), .op(n148) );
  nand2_1 U338 ( .ip1(hcr_ic_ss_hcnt[13]), .ip2(n603), .op(n147) );
  nand2_1 U339 ( .ip1(n148), .ip2(n147), .op(n1498) );
  nand2_1 U340 ( .ip1(ipwdata[15]), .ip2(n144), .op(n150) );
  nand2_1 U341 ( .ip1(hcr_ic_ss_hcnt[15]), .ip2(n603), .op(n149) );
  nand2_1 U342 ( .ip1(n150), .ip2(n149), .op(n1504) );
  nand2_1 U343 ( .ip1(ipwdata[14]), .ip2(n144), .op(n152) );
  nand2_1 U344 ( .ip1(hcr_ic_ss_hcnt[14]), .ip2(n603), .op(n151) );
  nand2_1 U345 ( .ip1(n152), .ip2(n151), .op(n1497) );
  nand2_1 U346 ( .ip1(ipwdata[11]), .ip2(n144), .op(n154) );
  nand2_1 U347 ( .ip1(hcr_ic_ss_hcnt[11]), .ip2(n603), .op(n153) );
  nand2_1 U348 ( .ip1(n154), .ip2(n153), .op(n1500) );
  nand2_1 U349 ( .ip1(ipwdata[10]), .ip2(n144), .op(n156) );
  nand2_1 U350 ( .ip1(hcr_ic_ss_hcnt[10]), .ip2(n603), .op(n155) );
  nand2_1 U351 ( .ip1(n156), .ip2(n155), .op(n1501) );
  nand2_1 U352 ( .ip1(ipwdata[9]), .ip2(n144), .op(n158) );
  nand2_1 U353 ( .ip1(hcr_ic_ss_hcnt[9]), .ip2(n603), .op(n157) );
  nand2_1 U354 ( .ip1(n158), .ip2(n157), .op(n1502) );
  nand2_1 U355 ( .ip1(ipwdata[8]), .ip2(n144), .op(n160) );
  nand2_1 U356 ( .ip1(hcr_ic_ss_hcnt[8]), .ip2(n603), .op(n159) );
  nand2_1 U357 ( .ip1(n160), .ip2(n159), .op(n1503) );
  nand2_1 U358 ( .ip1(ipwdata[12]), .ip2(n192), .op(n163) );
  nand2_1 U359 ( .ip1(ic_fs_hcnt[12]), .ip2(n605), .op(n162) );
  nand2_1 U360 ( .ip1(n163), .ip2(n162), .op(n1467) );
  nand2_1 U361 ( .ip1(ipwdata[13]), .ip2(n192), .op(n165) );
  nand2_1 U362 ( .ip1(ic_fs_hcnt[13]), .ip2(n605), .op(n164) );
  nand2_1 U363 ( .ip1(n165), .ip2(n164), .op(n1466) );
  nand2_1 U364 ( .ip1(ipwdata[15]), .ip2(n192), .op(n167) );
  nand2_1 U365 ( .ip1(ic_fs_hcnt[15]), .ip2(n605), .op(n166) );
  nand2_1 U366 ( .ip1(n167), .ip2(n166), .op(n1472) );
  nand2_1 U367 ( .ip1(ipwdata[14]), .ip2(n192), .op(n169) );
  nand2_1 U368 ( .ip1(ic_fs_hcnt[14]), .ip2(n605), .op(n168) );
  nand2_1 U369 ( .ip1(n169), .ip2(n168), .op(n1465) );
  nand2_1 U370 ( .ip1(ipwdata[7]), .ip2(n144), .op(n171) );
  nand2_1 U371 ( .ip1(hcr_ic_ss_hcnt[7]), .ip2(n603), .op(n170) );
  nand2_1 U372 ( .ip1(n171), .ip2(n170), .op(n1505) );
  nand2_1 U373 ( .ip1(ipwdata[10]), .ip2(n192), .op(n173) );
  nand2_1 U374 ( .ip1(ic_fs_hcnt[10]), .ip2(n605), .op(n172) );
  nand2_1 U375 ( .ip1(n173), .ip2(n172), .op(n1469) );
  nand2_1 U376 ( .ip1(ipwdata[3]), .ip2(n144), .op(n175) );
  nand2_1 U377 ( .ip1(hcr_ic_ss_hcnt[3]), .ip2(n603), .op(n174) );
  nand2_1 U378 ( .ip1(n175), .ip2(n174), .op(n1509) );
  nand2_1 U379 ( .ip1(ipwdata[11]), .ip2(n192), .op(n177) );
  nand2_1 U380 ( .ip1(ic_fs_hcnt[11]), .ip2(n605), .op(n176) );
  nand2_1 U381 ( .ip1(n177), .ip2(n176), .op(n1468) );
  nand2_1 U382 ( .ip1(ipwdata[4]), .ip2(n144), .op(n179) );
  nand2_1 U383 ( .ip1(hcr_ic_ss_hcnt[4]), .ip2(n603), .op(n178) );
  nand2_1 U384 ( .ip1(n179), .ip2(n178), .op(n1508) );
  nand2_1 U385 ( .ip1(ipwdata[9]), .ip2(n192), .op(n181) );
  nand2_1 U386 ( .ip1(ic_fs_hcnt[9]), .ip2(n605), .op(n180) );
  nand2_1 U387 ( .ip1(n181), .ip2(n180), .op(n1470) );
  nand2_1 U388 ( .ip1(ipwdata[0]), .ip2(n144), .op(n183) );
  nand2_1 U389 ( .ip1(hcr_ic_ss_hcnt[0]), .ip2(n603), .op(n182) );
  nand2_1 U390 ( .ip1(n183), .ip2(n182), .op(n1512) );
  nand2_1 U391 ( .ip1(ipwdata[8]), .ip2(n192), .op(n185) );
  nand2_1 U392 ( .ip1(ic_fs_hcnt[8]), .ip2(n605), .op(n184) );
  nand2_1 U393 ( .ip1(n185), .ip2(n184), .op(n1471) );
  nand2_1 U394 ( .ip1(ipwdata[7]), .ip2(n192), .op(n187) );
  nand2_1 U395 ( .ip1(ic_fs_hcnt[7]), .ip2(n605), .op(n186) );
  nand2_1 U396 ( .ip1(n187), .ip2(n186), .op(n1473) );
  nand2_1 U397 ( .ip1(ipwdata[3]), .ip2(n192), .op(n189) );
  nand2_1 U398 ( .ip1(ic_fs_hcnt[3]), .ip2(n605), .op(n188) );
  nand2_1 U399 ( .ip1(n189), .ip2(n188), .op(n1477) );
  nand2_1 U400 ( .ip1(ipwdata[4]), .ip2(n192), .op(n191) );
  nand2_1 U401 ( .ip1(ic_fs_hcnt[4]), .ip2(n605), .op(n190) );
  nand2_1 U402 ( .ip1(n191), .ip2(n190), .op(n1476) );
  nand2_1 U403 ( .ip1(ipwdata[0]), .ip2(n192), .op(n194) );
  nand2_1 U404 ( .ip1(ic_fs_hcnt[0]), .ip2(n605), .op(n193) );
  nand2_1 U405 ( .ip1(n194), .ip2(n193), .op(n1480) );
  inv_1 U406 ( .ip(iprdata[29]), .op(n355) );
  nand2_1 U407 ( .ip1(n678), .ip2(ic_txflr_flushed[1]), .op(n195) );
  nand2_1 U408 ( .ip1(n355), .ip2(n195), .op(iprdata[24]) );
  nand2_1 U409 ( .ip1(n677), .ip2(ic_sda_hold[21]), .op(n196) );
  nand2_1 U410 ( .ip1(n355), .ip2(n196), .op(iprdata[21]) );
  nand2_1 U411 ( .ip1(ic_sda_hold[20]), .ip2(n677), .op(n197) );
  inv_1 U412 ( .ip(iprdata[30]), .op(n450) );
  nand3_1 U413 ( .ip1(n197), .ip2(n450), .ip3(n355), .op(iprdata[20]) );
  nand2_1 U414 ( .ip1(ic_sda_hold[17]), .ip2(n677), .op(n200) );
  or2_1 U415 ( .ip1(n199), .ip2(n198), .op(n454) );
  nand3_1 U416 ( .ip1(n200), .ip2(n454), .ip3(n355), .op(iprdata[17]) );
  nand2_1 U417 ( .ip1(n678), .ip2(ic_txflr_flushed[3]), .op(n201) );
  nand2_1 U418 ( .ip1(n450), .ip2(n201), .op(iprdata[26]) );
  nand2_1 U419 ( .ip1(ic_clr_stop_det_en), .ip2(ic_raw_intr_stat[9]), .op(n205) );
  inv_1 U420 ( .ip(ic_clr_start_det_en), .op(n203) );
  nor2_1 U421 ( .ip1(ic_raw_intr_stat[10]), .ip2(n203), .op(n202) );
  or2_1 U422 ( .ip1(n203), .ip2(n202), .op(n204) );
  nand2_1 U423 ( .ip1(n205), .ip2(n204), .op(n213) );
  nand2_1 U424 ( .ip1(n649), .ip2(ic_tar[0]), .op(n211) );
  or2_1 U425 ( .ip1(n638), .ip2(ic_clr_rx_under_en), .op(n206) );
  nand2_1 U426 ( .ip1(ic_raw_intr_stat[0]), .ip2(n206), .op(n210) );
  nor2_1 U427 ( .ip1(n208), .ip2(n207), .op(n574) );
  nand2_1 U428 ( .ip1(ic_ack_general_call), .ip2(n574), .op(n209) );
  nand3_1 U429 ( .ip1(n211), .ip2(n210), .ip3(n209), .op(n212) );
  not_ab_or_c_or_d U430 ( .ip1(n676), .ip2(ic_hs_spklen[0]), .ip3(n213), .ip4(
        n212), .op(n260) );
  nand2_1 U431 ( .ip1(ic_txflr[0]), .ip2(n640), .op(n217) );
  nand2_1 U432 ( .ip1(n648), .ip2(hcr_ic_hs_lcnt[0]), .op(n216) );
  nand2_1 U433 ( .ip1(n641), .ip2(hcr_ic_ss_hcnt[0]), .op(n215) );
  nand2_1 U434 ( .ip1(n632), .ip2(ic_fs_hcnt[0]), .op(n214) );
  nand4_1 U435 ( .ip1(n217), .ip2(n216), .ip3(n215), .ip4(n214), .op(n222) );
  nand2_1 U436 ( .ip1(n633), .ip2(hcr_ic_ss_lcnt[0]), .op(n220) );
  nand2_1 U437 ( .ip1(ic_sda_hold[0]), .ip2(n677), .op(n219) );
  nand2_1 U438 ( .ip1(ic_hs_maddr[0]), .ip2(n619), .op(n218) );
  nand3_1 U439 ( .ip1(n220), .ip2(n219), .ip3(n218), .op(n221) );
  not_ab_or_c_or_d U440 ( .ip1(ic_clr_gen_call_en), .ip2(ic_raw_intr_stat[11]), 
        .ip3(n222), .ip4(n221), .op(n259) );
  nand2_1 U441 ( .ip1(n660), .ip2(ic_sda_setup[0]), .op(n226) );
  nand2_1 U442 ( .ip1(n658), .ip2(ic_intr_stat[0]), .op(n225) );
  nand2_1 U443 ( .ip1(n661), .ip2(ic_intr_mask[0]), .op(n224) );
  nand2_1 U444 ( .ip1(n669), .ip2(ic_sar[0]), .op(n223) );
  nand4_1 U445 ( .ip1(n226), .ip2(n225), .ip3(n224), .ip4(n223), .op(n231) );
  nand2_1 U446 ( .ip1(n668), .ip2(rx_pop_data[0]), .op(n229) );
  nand2_1 U447 ( .ip1(ic_rxflr[0]), .ip2(n639), .op(n228) );
  nand2_1 U448 ( .ip1(n404), .ip2(activity_r), .op(n227) );
  nand3_1 U449 ( .ip1(n229), .ip2(n228), .ip3(n227), .op(n230) );
  not_ab_or_c_or_d U450 ( .ip1(ic_clr_activity_en), .ip2(ic_raw_intr_stat[8]), 
        .ip3(n231), .ip4(n230), .op(n258) );
  nand2_1 U451 ( .ip1(ic_fs_spklen[0]), .ip2(n650), .op(n235) );
  nand2_1 U452 ( .ip1(ic_master), .ip2(n651), .op(n234) );
  nand2_1 U453 ( .ip1(n652), .ip2(ic_fs_lcnt[0]), .op(n233) );
  nand2_1 U454 ( .ip1(n678), .ip2(ic_tx_abrt_source[0]), .op(n232) );
  nand4_1 U455 ( .ip1(n235), .ip2(n234), .ip3(n233), .ip4(n232), .op(n256) );
  and2_1 U456 ( .ip1(ic_clr_rx_over_en), .ip2(ic_raw_intr_stat[1]), .op(n236)
         );
  mux2_1 U457 ( .ip1(n236), .ip2(ic_raw_intr_stat[3]), .s(ic_clr_tx_over_en), 
        .op(n237) );
  mux2_1 U458 ( .ip1(n237), .ip2(ic_raw_intr_stat[5]), .s(ic_clr_rd_req_en), 
        .op(n239) );
  mux2_1 U459 ( .ip1(ic_raw_intr_stat[6]), .ip2(n239), .s(n238), .op(n240) );
  mux2_1 U460 ( .ip1(n240), .ip2(ic_raw_intr_stat[7]), .s(ic_clr_rx_done_en), 
        .op(n255) );
  nor3_1 U461 ( .ip1(n242), .ip2(n241), .ip3(n706), .op(n244) );
  and2_1 U462 ( .ip1(ic_tx_tl_0_), .ip2(n576), .op(n243) );
  not_ab_or_c_or_d U463 ( .ip1(n245), .ip2(ic_en), .ip3(n244), .ip4(n243), 
        .op(n253) );
  nand2_1 U464 ( .ip1(n659), .ip2(hcr_ic_hs_hcnt[0]), .op(n252) );
  nor4_1 U465 ( .ip1(ic_raw_intr_stat[1]), .ip2(ic_raw_intr_stat[3]), .ip3(
        ic_raw_intr_stat[0]), .ip4(ic_raw_intr_stat[2]), .op(n248) );
  nor4_1 U466 ( .ip1(ic_raw_intr_stat[9]), .ip2(ic_raw_intr_stat[10]), .ip3(
        ic_raw_intr_stat[11]), .ip4(ic_raw_intr_stat[4]), .op(n247) );
  nor4_1 U467 ( .ip1(ic_raw_intr_stat[5]), .ip2(ic_raw_intr_stat[6]), .ip3(
        ic_raw_intr_stat[7]), .ip4(ic_raw_intr_stat[8]), .op(n246) );
  nand3_1 U468 ( .ip1(n248), .ip2(n247), .ip3(n246), .op(n249) );
  nand2_1 U469 ( .ip1(ic_clr_intr_en), .ip2(n249), .op(n251) );
  nand2_1 U470 ( .ip1(ic_rx_tl_int[0]), .ip2(n578), .op(n250) );
  nand4_1 U471 ( .ip1(n253), .ip2(n252), .ip3(n251), .ip4(n250), .op(n254) );
  nor3_1 U472 ( .ip1(n256), .ip2(n255), .ip3(n254), .op(n257) );
  nand4_1 U473 ( .ip1(n260), .ip2(n259), .ip3(n258), .ip4(n257), .op(
        iprdata[0]) );
  nand2_1 U474 ( .ip1(ic_raw_intr_stat[7]), .ip2(n638), .op(n264) );
  nand2_1 U475 ( .ip1(n641), .ip2(hcr_ic_ss_hcnt[7]), .op(n263) );
  nand2_1 U476 ( .ip1(n648), .ip2(hcr_ic_hs_lcnt[7]), .op(n262) );
  nand2_1 U477 ( .ip1(n632), .ip2(ic_fs_hcnt[7]), .op(n261) );
  and4_1 U478 ( .ip1(n264), .ip2(n263), .ip3(n262), .ip4(n261), .op(n282) );
  nand2_1 U479 ( .ip1(n660), .ip2(ic_sda_setup[7]), .op(n268) );
  nand2_1 U480 ( .ip1(n661), .ip2(ic_intr_mask[7]), .op(n267) );
  nand2_1 U481 ( .ip1(n669), .ip2(ic_sar[7]), .op(n266) );
  nand2_1 U482 ( .ip1(n668), .ip2(rx_pop_data[7]), .op(n265) );
  nand4_1 U483 ( .ip1(n268), .ip2(n267), .ip3(n266), .ip4(n265), .op(n269) );
  not_ab_or_c_or_d U484 ( .ip1(n658), .ip2(ic_intr_stat[7]), .ip3(n657), .ip4(
        n269), .op(n281) );
  nand2_1 U485 ( .ip1(n650), .ip2(ic_fs_spklen[7]), .op(n272) );
  nand2_1 U486 ( .ip1(n633), .ip2(hcr_ic_ss_lcnt[7]), .op(n271) );
  nand2_1 U487 ( .ip1(n677), .ip2(ic_sda_hold[7]), .op(n270) );
  nand3_1 U488 ( .ip1(n272), .ip2(n271), .ip3(n270), .op(n278) );
  nand2_1 U489 ( .ip1(n651), .ip2(p_det_ifaddr), .op(n276) );
  nand2_1 U490 ( .ip1(n649), .ip2(ic_tar[7]), .op(n275) );
  nand2_1 U491 ( .ip1(n652), .ip2(ic_fs_lcnt[7]), .op(n274) );
  nand2_1 U492 ( .ip1(n678), .ip2(ic_tx_abrt_source[7]), .op(n273) );
  nand4_1 U493 ( .ip1(n276), .ip2(n275), .ip3(n274), .ip4(n273), .op(n277) );
  not_ab_or_c_or_d U494 ( .ip1(n676), .ip2(ic_hs_spklen[7]), .ip3(n278), .ip4(
        n277), .op(n280) );
  nand2_1 U495 ( .ip1(n659), .ip2(hcr_ic_hs_hcnt[7]), .op(n279) );
  nand4_1 U496 ( .ip1(n282), .ip2(n281), .ip3(n280), .ip4(n279), .op(
        iprdata[7]) );
  nand2_1 U497 ( .ip1(n641), .ip2(hcr_ic_ss_hcnt[4]), .op(n286) );
  nand2_1 U498 ( .ip1(n404), .ip2(rx_full), .op(n285) );
  nand2_1 U499 ( .ip1(n648), .ip2(hcr_ic_hs_lcnt[4]), .op(n284) );
  nand2_1 U500 ( .ip1(n632), .ip2(ic_fs_hcnt[4]), .op(n283) );
  and4_1 U501 ( .ip1(n286), .ip2(n285), .ip3(n284), .ip4(n283), .op(n305) );
  and2_1 U502 ( .ip1(n661), .ip2(ic_intr_mask[4]), .op(n292) );
  nand2_1 U503 ( .ip1(n658), .ip2(ic_intr_stat[4]), .op(n290) );
  nand2_1 U504 ( .ip1(n660), .ip2(ic_sda_setup[4]), .op(n289) );
  nand2_1 U505 ( .ip1(n668), .ip2(rx_pop_data[4]), .op(n288) );
  nand2_1 U506 ( .ip1(n638), .ip2(ic_raw_intr_stat[4]), .op(n287) );
  nand4_1 U507 ( .ip1(n290), .ip2(n289), .ip3(n288), .ip4(n287), .op(n291) );
  not_ab_or_c_or_d U508 ( .ip1(n669), .ip2(ic_sar[4]), .ip3(n292), .ip4(n291), 
        .op(n304) );
  nand2_1 U509 ( .ip1(n650), .ip2(ic_fs_spklen[4]), .op(n295) );
  nand2_1 U510 ( .ip1(n633), .ip2(hcr_ic_ss_lcnt[4]), .op(n294) );
  nand2_1 U511 ( .ip1(n677), .ip2(ic_sda_hold[4]), .op(n293) );
  nand3_1 U512 ( .ip1(n295), .ip2(n294), .ip3(n293), .op(n301) );
  nand2_1 U513 ( .ip1(n651), .ip2(ic_10bit_mst), .op(n299) );
  nand2_1 U514 ( .ip1(n649), .ip2(ic_tar[4]), .op(n298) );
  nand2_1 U515 ( .ip1(n652), .ip2(ic_fs_lcnt[4]), .op(n297) );
  nand2_1 U516 ( .ip1(n678), .ip2(ic_tx_abrt_source[4]), .op(n296) );
  nand4_1 U517 ( .ip1(n299), .ip2(n298), .ip3(n297), .ip4(n296), .op(n300) );
  not_ab_or_c_or_d U518 ( .ip1(n676), .ip2(ic_hs_spklen[4]), .ip3(n301), .ip4(
        n300), .op(n303) );
  nand2_1 U519 ( .ip1(n659), .ip2(hcr_ic_hs_hcnt[4]), .op(n302) );
  nand4_1 U520 ( .ip1(n305), .ip2(n304), .ip3(n303), .ip4(n302), .op(
        iprdata[4]) );
  and2_1 U521 ( .ip1(n658), .ip2(ic_intr_stat[10]), .op(n306) );
  not_ab_or_c_or_d U522 ( .ip1(n678), .ip2(ic_tx_abrt_source[10]), .ip3(n306), 
        .ip4(n657), .op(n319) );
  nand2_1 U523 ( .ip1(n661), .ip2(ic_intr_mask[10]), .op(n310) );
  nand2_1 U524 ( .ip1(ic_raw_intr_stat[10]), .ip2(n638), .op(n309) );
  nand2_1 U525 ( .ip1(n641), .ip2(hcr_ic_ss_hcnt[10]), .op(n308) );
  nand2_1 U526 ( .ip1(n648), .ip2(hcr_ic_hs_lcnt[10]), .op(n307) );
  nand4_1 U527 ( .ip1(n310), .ip2(n309), .ip3(n308), .ip4(n307), .op(n315) );
  nand2_1 U528 ( .ip1(ic_fs_hcnt[10]), .ip2(n632), .op(n313) );
  nand2_1 U529 ( .ip1(n633), .ip2(hcr_ic_ss_lcnt[10]), .op(n312) );
  nand2_1 U530 ( .ip1(n677), .ip2(ic_sda_hold[10]), .op(n311) );
  nand3_1 U531 ( .ip1(n313), .ip2(n312), .ip3(n311), .op(n314) );
  not_ab_or_c_or_d U532 ( .ip1(n649), .ip2(ic_tar[10]), .ip3(n315), .ip4(n314), 
        .op(n318) );
  nand2_1 U533 ( .ip1(n652), .ip2(ic_fs_lcnt[10]), .op(n317) );
  nand2_1 U534 ( .ip1(n659), .ip2(hcr_ic_hs_hcnt[10]), .op(n316) );
  nand4_1 U535 ( .ip1(n319), .ip2(n318), .ip3(n317), .ip4(n316), .op(
        iprdata[10]) );
  nand2_1 U536 ( .ip1(n648), .ip2(hcr_ic_hs_lcnt[15]), .op(n328) );
  and2_1 U537 ( .ip1(n632), .ip2(ic_fs_hcnt[15]), .op(n325) );
  nand2_1 U538 ( .ip1(n652), .ip2(ic_fs_lcnt[15]), .op(n323) );
  nand2_1 U539 ( .ip1(n677), .ip2(ic_sda_hold[15]), .op(n322) );
  nand2_1 U540 ( .ip1(n678), .ip2(ic_tx_abrt_source[15]), .op(n321) );
  nand2_1 U541 ( .ip1(n659), .ip2(hcr_ic_hs_hcnt[15]), .op(n320) );
  nand4_1 U542 ( .ip1(n323), .ip2(n322), .ip3(n321), .ip4(n320), .op(n324) );
  not_ab_or_c_or_d U543 ( .ip1(n633), .ip2(hcr_ic_ss_lcnt[15]), .ip3(n325), 
        .ip4(n324), .op(n327) );
  nand2_1 U544 ( .ip1(n641), .ip2(hcr_ic_ss_hcnt[15]), .op(n326) );
  nand3_1 U545 ( .ip1(n328), .ip2(n327), .ip3(n326), .op(iprdata[15]) );
  nand2_1 U546 ( .ip1(n648), .ip2(hcr_ic_hs_lcnt[14]), .op(n337) );
  and2_1 U547 ( .ip1(n632), .ip2(ic_fs_hcnt[14]), .op(n334) );
  nand2_1 U548 ( .ip1(n652), .ip2(ic_fs_lcnt[14]), .op(n332) );
  nand2_1 U549 ( .ip1(n677), .ip2(ic_sda_hold[14]), .op(n331) );
  nand2_1 U550 ( .ip1(n678), .ip2(ic_tx_abrt_source[14]), .op(n330) );
  nand2_1 U551 ( .ip1(n659), .ip2(hcr_ic_hs_hcnt[14]), .op(n329) );
  nand4_1 U552 ( .ip1(n332), .ip2(n331), .ip3(n330), .ip4(n329), .op(n333) );
  not_ab_or_c_or_d U553 ( .ip1(n633), .ip2(hcr_ic_ss_lcnt[14]), .ip3(n334), 
        .ip4(n333), .op(n336) );
  nand2_1 U554 ( .ip1(n641), .ip2(hcr_ic_ss_hcnt[14]), .op(n335) );
  nand3_1 U555 ( .ip1(n337), .ip2(n336), .ip3(n335), .op(iprdata[14]) );
  and2_1 U556 ( .ip1(n632), .ip2(ic_fs_hcnt[13]), .op(n343) );
  nand2_1 U557 ( .ip1(n633), .ip2(hcr_ic_ss_lcnt[13]), .op(n341) );
  nand2_1 U558 ( .ip1(n677), .ip2(ic_sda_hold[13]), .op(n340) );
  nand2_1 U559 ( .ip1(n652), .ip2(ic_fs_lcnt[13]), .op(n339) );
  nand2_1 U560 ( .ip1(n678), .ip2(ic_tx_abrt_source[13]), .op(n338) );
  nand4_1 U561 ( .ip1(n341), .ip2(n340), .ip3(n339), .ip4(n338), .op(n342) );
  not_ab_or_c_or_d U562 ( .ip1(hcr_ic_hs_lcnt[13]), .ip2(n648), .ip3(n343), 
        .ip4(n342), .op(n346) );
  nand2_1 U563 ( .ip1(n641), .ip2(hcr_ic_ss_hcnt[13]), .op(n345) );
  nand2_1 U564 ( .ip1(n659), .ip2(hcr_ic_hs_hcnt[13]), .op(n344) );
  nand4_1 U565 ( .ip1(n346), .ip2(n355), .ip3(n345), .ip4(n344), .op(
        iprdata[13]) );
  and2_1 U566 ( .ip1(n632), .ip2(ic_fs_hcnt[12]), .op(n352) );
  nand2_1 U567 ( .ip1(n633), .ip2(hcr_ic_ss_lcnt[12]), .op(n350) );
  nand2_1 U568 ( .ip1(n677), .ip2(ic_sda_hold[12]), .op(n349) );
  nand2_1 U569 ( .ip1(n652), .ip2(ic_fs_lcnt[12]), .op(n348) );
  nand2_1 U570 ( .ip1(n678), .ip2(ic_tx_abrt_source[12]), .op(n347) );
  nand4_1 U571 ( .ip1(n350), .ip2(n349), .ip3(n348), .ip4(n347), .op(n351) );
  not_ab_or_c_or_d U572 ( .ip1(hcr_ic_hs_lcnt[12]), .ip2(n648), .ip3(n352), 
        .ip4(n351), .op(n356) );
  nand2_1 U573 ( .ip1(n641), .ip2(hcr_ic_ss_hcnt[12]), .op(n354) );
  nand2_1 U574 ( .ip1(n659), .ip2(hcr_ic_hs_hcnt[12]), .op(n353) );
  nand4_1 U575 ( .ip1(n356), .ip2(n355), .ip3(n354), .ip4(n353), .op(
        iprdata[12]) );
  nand2_1 U576 ( .ip1(n661), .ip2(ic_intr_mask[8]), .op(n360) );
  nand2_1 U577 ( .ip1(n669), .ip2(ic_sar[8]), .op(n359) );
  nand2_1 U578 ( .ip1(n638), .ip2(ic_raw_intr_stat[8]), .op(n358) );
  nand2_1 U579 ( .ip1(n648), .ip2(hcr_ic_hs_lcnt[8]), .op(n357) );
  nand4_1 U580 ( .ip1(n360), .ip2(n359), .ip3(n358), .ip4(n357), .op(n371) );
  nand2_1 U581 ( .ip1(n641), .ip2(hcr_ic_ss_hcnt[8]), .op(n364) );
  nand2_1 U582 ( .ip1(n632), .ip2(ic_fs_hcnt[8]), .op(n363) );
  nand2_1 U583 ( .ip1(n633), .ip2(hcr_ic_ss_lcnt[8]), .op(n362) );
  nand2_1 U584 ( .ip1(n677), .ip2(ic_sda_hold[8]), .op(n361) );
  nand4_1 U585 ( .ip1(n364), .ip2(n363), .ip3(n362), .ip4(n361), .op(n370) );
  nand2_1 U586 ( .ip1(n651), .ip2(tx_empty_ctrl), .op(n368) );
  nand2_1 U587 ( .ip1(n649), .ip2(ic_tar[8]), .op(n367) );
  nand2_1 U588 ( .ip1(n652), .ip2(ic_fs_lcnt[8]), .op(n366) );
  nand2_1 U589 ( .ip1(n659), .ip2(hcr_ic_hs_hcnt[8]), .op(n365) );
  nand4_1 U590 ( .ip1(n368), .ip2(n367), .ip3(n366), .ip4(n365), .op(n369) );
  nor3_1 U591 ( .ip1(n371), .ip2(n370), .ip3(n369), .op(n374) );
  nand2_1 U592 ( .ip1(n658), .ip2(ic_intr_stat[8]), .op(n373) );
  nand2_1 U593 ( .ip1(n678), .ip2(ic_tx_abrt_source[8]), .op(n372) );
  nand4_1 U594 ( .ip1(n374), .ip2(n454), .ip3(n373), .ip4(n372), .op(
        iprdata[8]) );
  nand2_1 U595 ( .ip1(n669), .ip2(ic_sar[5]), .op(n378) );
  nand2_1 U596 ( .ip1(n668), .ip2(rx_pop_data[5]), .op(n377) );
  nand2_1 U597 ( .ip1(ic_raw_intr_stat[5]), .ip2(n638), .op(n376) );
  nand2_1 U598 ( .ip1(n648), .ip2(hcr_ic_hs_lcnt[5]), .op(n375) );
  nand4_1 U599 ( .ip1(n378), .ip2(n377), .ip3(n376), .ip4(n375), .op(n379) );
  not_ab_or_c_or_d U600 ( .ip1(n658), .ip2(ic_intr_stat[5]), .ip3(iprdata[29]), 
        .ip4(n379), .op(n398) );
  nand2_1 U601 ( .ip1(n404), .ip2(mst_activity_r), .op(n383) );
  nand2_1 U602 ( .ip1(n641), .ip2(hcr_ic_ss_hcnt[5]), .op(n382) );
  nand2_1 U603 ( .ip1(n677), .ip2(ic_sda_hold[5]), .op(n381) );
  nand2_1 U604 ( .ip1(n632), .ip2(ic_fs_hcnt[5]), .op(n380) );
  nand4_1 U605 ( .ip1(n383), .ip2(n382), .ip3(n381), .ip4(n380), .op(n394) );
  nand2_1 U606 ( .ip1(n676), .ip2(ic_hs_spklen[5]), .op(n387) );
  nand2_1 U607 ( .ip1(n650), .ip2(ic_fs_spklen[5]), .op(n386) );
  nand2_1 U608 ( .ip1(n651), .ip2(ic_rstrt_en), .op(n385) );
  nand2_1 U609 ( .ip1(n633), .ip2(hcr_ic_ss_lcnt[5]), .op(n384) );
  nand4_1 U610 ( .ip1(n387), .ip2(n386), .ip3(n385), .ip4(n384), .op(n393) );
  nand2_1 U611 ( .ip1(n649), .ip2(ic_tar[5]), .op(n391) );
  nand2_1 U612 ( .ip1(n652), .ip2(ic_fs_lcnt[5]), .op(n390) );
  nand2_1 U613 ( .ip1(n678), .ip2(ic_tx_abrt_source[5]), .op(n389) );
  nand2_1 U614 ( .ip1(n659), .ip2(hcr_ic_hs_hcnt[5]), .op(n388) );
  nand4_1 U615 ( .ip1(n391), .ip2(n390), .ip3(n389), .ip4(n388), .op(n392) );
  nor3_1 U616 ( .ip1(n394), .ip2(n393), .ip3(n392), .op(n397) );
  nand2_1 U617 ( .ip1(n660), .ip2(ic_sda_setup[5]), .op(n396) );
  nand2_1 U618 ( .ip1(n661), .ip2(ic_intr_mask[5]), .op(n395) );
  nand4_1 U619 ( .ip1(n398), .ip2(n397), .ip3(n396), .ip4(n395), .op(
        iprdata[5]) );
  nand2_1 U620 ( .ip1(n669), .ip2(ic_sar[6]), .op(n402) );
  nand2_1 U621 ( .ip1(n668), .ip2(rx_pop_data[6]), .op(n401) );
  nand2_1 U622 ( .ip1(ic_raw_intr_stat[6]), .ip2(n638), .op(n400) );
  nand2_1 U623 ( .ip1(n648), .ip2(hcr_ic_hs_lcnt[6]), .op(n399) );
  nand4_1 U624 ( .ip1(n402), .ip2(n401), .ip3(n400), .ip4(n399), .op(n403) );
  not_ab_or_c_or_d U625 ( .ip1(n658), .ip2(ic_intr_stat[6]), .ip3(iprdata[30]), 
        .ip4(n403), .op(n423) );
  nand2_1 U626 ( .ip1(n404), .ip2(slv_activity_r), .op(n408) );
  nand2_1 U627 ( .ip1(n641), .ip2(hcr_ic_ss_hcnt[6]), .op(n407) );
  nand2_1 U628 ( .ip1(n677), .ip2(ic_sda_hold[6]), .op(n406) );
  nand2_1 U629 ( .ip1(n632), .ip2(ic_fs_hcnt[6]), .op(n405) );
  nand4_1 U630 ( .ip1(n408), .ip2(n407), .ip3(n406), .ip4(n405), .op(n419) );
  nand2_1 U631 ( .ip1(n676), .ip2(ic_hs_spklen[6]), .op(n412) );
  nand2_1 U632 ( .ip1(n650), .ip2(ic_fs_spklen[6]), .op(n411) );
  nand2_1 U633 ( .ip1(n651), .ip2(ic_con_pre_6_), .op(n410) );
  nand2_1 U634 ( .ip1(n633), .ip2(hcr_ic_ss_lcnt[6]), .op(n409) );
  nand4_1 U635 ( .ip1(n412), .ip2(n411), .ip3(n410), .ip4(n409), .op(n418) );
  nand2_1 U636 ( .ip1(n649), .ip2(ic_tar[6]), .op(n416) );
  nand2_1 U637 ( .ip1(n652), .ip2(ic_fs_lcnt[6]), .op(n415) );
  nand2_1 U638 ( .ip1(n678), .ip2(ic_tx_abrt_source[6]), .op(n414) );
  nand2_1 U639 ( .ip1(n659), .ip2(hcr_ic_hs_hcnt[6]), .op(n413) );
  nand4_1 U640 ( .ip1(n416), .ip2(n415), .ip3(n414), .ip4(n413), .op(n417) );
  nor3_1 U641 ( .ip1(n419), .ip2(n418), .ip3(n417), .op(n422) );
  nand2_1 U642 ( .ip1(n660), .ip2(ic_sda_setup[6]), .op(n421) );
  nand2_1 U643 ( .ip1(n661), .ip2(ic_intr_mask[6]), .op(n420) );
  nand4_1 U644 ( .ip1(n423), .ip2(n422), .ip3(n421), .ip4(n420), .op(
        iprdata[6]) );
  not_ab_or_c_or_d U645 ( .ip1(n669), .ip2(ic_sar[9]), .ip3(iprdata[29]), 
        .ip4(n657), .op(n438) );
  nand2_1 U646 ( .ip1(n652), .ip2(ic_fs_lcnt[9]), .op(n426) );
  nand2_1 U647 ( .ip1(n633), .ip2(hcr_ic_ss_lcnt[9]), .op(n425) );
  nand2_1 U648 ( .ip1(n677), .ip2(ic_sda_hold[9]), .op(n424) );
  nand3_1 U649 ( .ip1(n426), .ip2(n425), .ip3(n424), .op(n434) );
  and2_1 U650 ( .ip1(n641), .ip2(hcr_ic_ss_hcnt[9]), .op(n428) );
  and2_1 U651 ( .ip1(n632), .ip2(ic_fs_hcnt[9]), .op(n427) );
  not_ab_or_c_or_d U652 ( .ip1(n648), .ip2(hcr_ic_hs_lcnt[9]), .ip3(n428), 
        .ip4(n427), .op(n432) );
  nand2_1 U653 ( .ip1(n659), .ip2(hcr_ic_hs_hcnt[9]), .op(n431) );
  nand2_1 U654 ( .ip1(n678), .ip2(ic_tx_abrt_source[9]), .op(n430) );
  nand2_1 U655 ( .ip1(ic_raw_intr_stat[9]), .ip2(n638), .op(n429) );
  nand4_1 U656 ( .ip1(n432), .ip2(n431), .ip3(n430), .ip4(n429), .op(n433) );
  not_ab_or_c_or_d U657 ( .ip1(n649), .ip2(ic_tar[9]), .ip3(n434), .ip4(n433), 
        .op(n437) );
  nand2_1 U658 ( .ip1(n658), .ip2(ic_intr_stat[9]), .op(n436) );
  nand2_1 U659 ( .ip1(n661), .ip2(ic_intr_mask[9]), .op(n435) );
  nand4_1 U660 ( .ip1(n438), .ip2(n437), .ip3(n436), .ip4(n435), .op(
        iprdata[9]) );
  inv_1 U661 ( .ip(tx_fifo_rst_n), .op(n441) );
  nor3_1 U662 ( .ip1(ic_txflr[0]), .ip2(ic_txflr[1]), .ip3(ic_txflr[2]), .op(
        n692) );
  inv_1 U663 ( .ip(ic_txflr[3]), .op(n701) );
  nand2_1 U664 ( .ip1(n668), .ip2(wr_en), .op(n440) );
  nand2_1 U665 ( .ip1(tx_fifo_rst_n), .ip2(tx_pop_sync), .op(n439) );
  not_ab_or_c_or_d U666 ( .ip1(n692), .ip2(n701), .ip3(tx_push), .ip4(n439), 
        .op(n693) );
  inv_1 U667 ( .ip(n693), .op(n442) );
  nor4_1 U668 ( .ip1(n441), .ip2(n440), .ip3(ic_txflr[3]), .ip4(tx_pop_sync), 
        .op(n610) );
  nor2_1 U669 ( .ip1(n442), .ip2(n692), .op(n443) );
  or2_1 U670 ( .ip1(n607), .ip2(n443), .op(n444) );
  nand2_1 U671 ( .ip1(ic_txflr[3]), .ip2(n444), .op(n447) );
  nand3_1 U672 ( .ip1(ic_txflr[0]), .ip2(ic_txflr[1]), .ip3(ic_txflr[2]), .op(
        n445) );
  mux2_1 U673 ( .ip1(ic_txflr[3]), .ip2(n701), .s(n445), .op(n700) );
  or2_1 U674 ( .ip1(n689), .ip2(n700), .op(n446) );
  nand2_1 U675 ( .ip1(n447), .ip2(n446), .op(n1364) );
  nand2_1 U676 ( .ip1(n677), .ip2(ic_sda_hold[18]), .op(n448) );
  nand2_1 U677 ( .ip1(n454), .ip2(n448), .op(iprdata[18]) );
  nand2_1 U678 ( .ip1(n677), .ip2(ic_sda_hold[22]), .op(n449) );
  nand2_1 U679 ( .ip1(n450), .ip2(n449), .op(iprdata[22]) );
  nand2_1 U680 ( .ip1(ic_sda_hold[23]), .ip2(n677), .op(n452) );
  nand2_1 U681 ( .ip1(ic_txflr_flushed[0]), .ip2(n678), .op(n451) );
  nand2_1 U682 ( .ip1(n452), .ip2(n451), .op(iprdata[23]) );
  nand2_1 U683 ( .ip1(ic_tx_abrt_source[16]), .ip2(n678), .op(n455) );
  nand2_1 U684 ( .ip1(n677), .ip2(ic_sda_hold[16]), .op(n453) );
  nand3_1 U685 ( .ip1(n455), .ip2(n454), .ip3(n453), .op(iprdata[16]) );
  or2_1 U686 ( .ip1(n706), .ip2(n456), .op(n458) );
  or2_1 U687 ( .ip1(n583), .ip2(n456), .op(n457) );
  nand2_1 U688 ( .ip1(n458), .ip2(n457), .op(n1549) );
  nand2_1 U689 ( .ip1(n658), .ip2(ic_intr_stat[11]), .op(n462) );
  nand2_1 U690 ( .ip1(n661), .ip2(ic_intr_mask[11]), .op(n461) );
  nand2_1 U691 ( .ip1(n638), .ip2(ic_raw_intr_stat[11]), .op(n460) );
  nand2_1 U692 ( .ip1(n641), .ip2(hcr_ic_ss_hcnt[11]), .op(n459) );
  and4_1 U693 ( .ip1(n462), .ip2(n461), .ip3(n460), .ip4(n459), .op(n472) );
  and2_1 U694 ( .ip1(n652), .ip2(ic_fs_lcnt[11]), .op(n468) );
  nand2_1 U695 ( .ip1(n648), .ip2(hcr_ic_hs_lcnt[11]), .op(n466) );
  nand2_1 U696 ( .ip1(n633), .ip2(hcr_ic_ss_lcnt[11]), .op(n465) );
  nand2_1 U697 ( .ip1(n632), .ip2(ic_fs_hcnt[11]), .op(n464) );
  nand2_1 U698 ( .ip1(n677), .ip2(ic_sda_hold[11]), .op(n463) );
  nand4_1 U699 ( .ip1(n466), .ip2(n465), .ip3(n464), .ip4(n463), .op(n467) );
  not_ab_or_c_or_d U700 ( .ip1(ic_tar[11]), .ip2(n649), .ip3(n468), .ip4(n467), 
        .op(n471) );
  nand2_1 U701 ( .ip1(n659), .ip2(hcr_ic_hs_hcnt[11]), .op(n470) );
  nand2_1 U702 ( .ip1(n678), .ip2(ic_tx_abrt_source[11]), .op(n469) );
  nand4_1 U703 ( .ip1(n472), .ip2(n471), .ip3(n470), .ip4(n469), .op(
        iprdata[11]) );
  mux2_1 U704 ( .ip1(n474), .ip2(n473), .s(ic_rxflr[0]), .op(n475) );
  inv_1 U705 ( .ip(n475), .op(n1546) );
  inv_1 U706 ( .ip(presetn), .op(n760) );
  inv_1 U707 ( .ip(presetn), .op(n485) );
  inv_1 U708 ( .ip(ic_con_pre_1_), .op(n570) );
  nand2_1 U709 ( .ip1(n570), .ip2(ic_fs_hcnt[15]), .op(n478) );
  inv_1 U710 ( .ip(ic_con_pre_2_), .op(n679) );
  nand2_1 U711 ( .ip1(hcr_ic_hs_hcnt[15]), .ip2(ic_hs), .op(n477) );
  nor2_1 U712 ( .ip1(ic_con_pre_2_), .ip2(n570), .op(ic_ss) );
  nand2_1 U713 ( .ip1(hcr_ic_ss_hcnt[15]), .ip2(ic_ss), .op(n476) );
  nand2_1 U714 ( .ip1(n570), .ip2(ic_fs_lcnt[14]), .op(n481) );
  nand2_1 U715 ( .ip1(hcr_ic_hs_lcnt[14]), .ip2(ic_hs), .op(n480) );
  nand2_1 U716 ( .ip1(hcr_ic_ss_lcnt[14]), .ip2(ic_ss), .op(n479) );
  nand2_1 U717 ( .ip1(n570), .ip2(ic_fs_lcnt[15]), .op(n484) );
  nand2_1 U718 ( .ip1(hcr_ic_hs_lcnt[15]), .ip2(ic_hs), .op(n483) );
  nand2_1 U719 ( .ip1(hcr_ic_ss_lcnt[15]), .ip2(ic_ss), .op(n482) );
  nand2_1 U720 ( .ip1(hcr_ic_hs_hcnt[0]), .ip2(ic_hs), .op(n488) );
  nand2_1 U721 ( .ip1(ic_fs_hcnt[0]), .ip2(n570), .op(n487) );
  nand2_1 U722 ( .ip1(hcr_ic_ss_hcnt[0]), .ip2(ic_ss), .op(n486) );
  nand3_1 U723 ( .ip1(n488), .ip2(n487), .ip3(n486), .op(ic_hcnt[0]) );
  nand2_1 U724 ( .ip1(n570), .ip2(ic_fs_hcnt[1]), .op(n491) );
  nand2_1 U725 ( .ip1(hcr_ic_hs_hcnt[1]), .ip2(ic_hs), .op(n490) );
  nand2_1 U726 ( .ip1(hcr_ic_ss_hcnt[1]), .ip2(ic_ss), .op(n489) );
  nand2_1 U727 ( .ip1(n570), .ip2(ic_fs_hcnt[2]), .op(n494) );
  nand2_1 U728 ( .ip1(hcr_ic_hs_hcnt[2]), .ip2(ic_hs), .op(n493) );
  nand2_1 U729 ( .ip1(hcr_ic_ss_hcnt[2]), .ip2(ic_ss), .op(n492) );
  nand2_1 U730 ( .ip1(n570), .ip2(ic_fs_hcnt[3]), .op(n497) );
  nand2_1 U731 ( .ip1(hcr_ic_hs_hcnt[3]), .ip2(ic_hs), .op(n496) );
  nand2_1 U732 ( .ip1(hcr_ic_ss_hcnt[3]), .ip2(ic_ss), .op(n495) );
  nand2_1 U733 ( .ip1(n570), .ip2(ic_fs_hcnt[4]), .op(n500) );
  nand2_1 U734 ( .ip1(hcr_ic_hs_hcnt[4]), .ip2(ic_hs), .op(n499) );
  nand2_1 U735 ( .ip1(hcr_ic_ss_hcnt[4]), .ip2(ic_ss), .op(n498) );
  nand2_1 U736 ( .ip1(n570), .ip2(ic_fs_hcnt[5]), .op(n503) );
  nand2_1 U737 ( .ip1(hcr_ic_hs_hcnt[5]), .ip2(ic_hs), .op(n502) );
  nand2_1 U738 ( .ip1(hcr_ic_ss_hcnt[5]), .ip2(ic_ss), .op(n501) );
  nand2_1 U739 ( .ip1(n570), .ip2(ic_fs_hcnt[6]), .op(n506) );
  nand2_1 U740 ( .ip1(hcr_ic_hs_hcnt[6]), .ip2(ic_hs), .op(n505) );
  nand2_1 U741 ( .ip1(hcr_ic_ss_hcnt[6]), .ip2(ic_ss), .op(n504) );
  nand2_1 U742 ( .ip1(n570), .ip2(ic_fs_hcnt[7]), .op(n509) );
  nand2_1 U743 ( .ip1(hcr_ic_hs_hcnt[7]), .ip2(ic_hs), .op(n508) );
  nand2_1 U744 ( .ip1(hcr_ic_ss_hcnt[7]), .ip2(ic_ss), .op(n507) );
  nand2_1 U745 ( .ip1(n570), .ip2(ic_fs_hcnt[14]), .op(n512) );
  nand2_1 U746 ( .ip1(hcr_ic_hs_hcnt[14]), .ip2(ic_hs), .op(n511) );
  nand2_1 U747 ( .ip1(hcr_ic_ss_hcnt[14]), .ip2(ic_ss), .op(n510) );
  nand2_1 U748 ( .ip1(n570), .ip2(ic_fs_hcnt[8]), .op(n515) );
  nand2_1 U749 ( .ip1(hcr_ic_hs_hcnt[8]), .ip2(ic_hs), .op(n514) );
  nand2_1 U750 ( .ip1(hcr_ic_ss_hcnt[8]), .ip2(ic_ss), .op(n513) );
  nand2_1 U751 ( .ip1(n570), .ip2(ic_fs_hcnt[10]), .op(n518) );
  nand2_1 U752 ( .ip1(hcr_ic_hs_hcnt[10]), .ip2(ic_hs), .op(n517) );
  nand2_1 U753 ( .ip1(hcr_ic_ss_hcnt[10]), .ip2(ic_ss), .op(n516) );
  nand2_1 U754 ( .ip1(n570), .ip2(ic_fs_hcnt[9]), .op(n521) );
  nand2_1 U755 ( .ip1(hcr_ic_hs_hcnt[9]), .ip2(ic_hs), .op(n520) );
  nand2_1 U756 ( .ip1(hcr_ic_ss_hcnt[9]), .ip2(ic_ss), .op(n519) );
  nand2_1 U757 ( .ip1(n570), .ip2(ic_fs_hcnt[13]), .op(n524) );
  nand2_1 U758 ( .ip1(hcr_ic_hs_hcnt[13]), .ip2(ic_hs), .op(n523) );
  nand2_1 U759 ( .ip1(hcr_ic_ss_hcnt[13]), .ip2(ic_ss), .op(n522) );
  nand2_1 U760 ( .ip1(n570), .ip2(ic_fs_hcnt[12]), .op(n527) );
  nand2_1 U761 ( .ip1(hcr_ic_hs_hcnt[12]), .ip2(ic_hs), .op(n526) );
  nand2_1 U762 ( .ip1(hcr_ic_ss_hcnt[12]), .ip2(ic_ss), .op(n525) );
  nand2_1 U763 ( .ip1(n570), .ip2(ic_fs_hcnt[11]), .op(n530) );
  nand2_1 U764 ( .ip1(hcr_ic_hs_hcnt[11]), .ip2(ic_hs), .op(n529) );
  nand2_1 U765 ( .ip1(hcr_ic_ss_hcnt[11]), .ip2(ic_ss), .op(n528) );
  nand2_1 U766 ( .ip1(n570), .ip2(ic_fs_lcnt[0]), .op(n533) );
  nand2_1 U767 ( .ip1(hcr_ic_ss_lcnt[0]), .ip2(ic_ss), .op(n532) );
  nand2_1 U768 ( .ip1(hcr_ic_hs_lcnt[0]), .ip2(ic_hs), .op(n531) );
  nand2_1 U769 ( .ip1(n570), .ip2(ic_fs_lcnt[1]), .op(n536) );
  nand2_1 U770 ( .ip1(hcr_ic_hs_lcnt[1]), .ip2(ic_hs), .op(n535) );
  nand2_1 U771 ( .ip1(hcr_ic_ss_lcnt[1]), .ip2(ic_ss), .op(n534) );
  nand2_1 U772 ( .ip1(n570), .ip2(ic_fs_lcnt[3]), .op(n539) );
  nand2_1 U773 ( .ip1(hcr_ic_hs_lcnt[3]), .ip2(ic_hs), .op(n538) );
  nand2_1 U774 ( .ip1(hcr_ic_ss_lcnt[3]), .ip2(ic_ss), .op(n537) );
  nand2_1 U775 ( .ip1(n570), .ip2(ic_fs_lcnt[2]), .op(n542) );
  nand2_1 U776 ( .ip1(hcr_ic_hs_lcnt[2]), .ip2(ic_hs), .op(n541) );
  nand2_1 U777 ( .ip1(hcr_ic_ss_lcnt[2]), .ip2(ic_ss), .op(n540) );
  nand2_1 U778 ( .ip1(n570), .ip2(ic_fs_lcnt[5]), .op(n545) );
  nand2_1 U779 ( .ip1(hcr_ic_hs_lcnt[5]), .ip2(ic_hs), .op(n544) );
  nand2_1 U780 ( .ip1(hcr_ic_ss_lcnt[5]), .ip2(ic_ss), .op(n543) );
  nand2_1 U781 ( .ip1(n570), .ip2(ic_fs_lcnt[4]), .op(n548) );
  nand2_1 U782 ( .ip1(hcr_ic_hs_lcnt[4]), .ip2(ic_hs), .op(n547) );
  nand2_1 U783 ( .ip1(hcr_ic_ss_lcnt[4]), .ip2(ic_ss), .op(n546) );
  nand2_1 U784 ( .ip1(n570), .ip2(ic_fs_lcnt[7]), .op(n551) );
  nand2_1 U785 ( .ip1(hcr_ic_hs_lcnt[7]), .ip2(ic_hs), .op(n550) );
  nand2_1 U786 ( .ip1(hcr_ic_ss_lcnt[7]), .ip2(ic_ss), .op(n549) );
  nand2_1 U787 ( .ip1(n570), .ip2(ic_fs_lcnt[6]), .op(n554) );
  nand2_1 U788 ( .ip1(hcr_ic_hs_lcnt[6]), .ip2(ic_hs), .op(n553) );
  nand2_1 U789 ( .ip1(hcr_ic_ss_lcnt[6]), .ip2(ic_ss), .op(n552) );
  nand2_1 U790 ( .ip1(n570), .ip2(ic_fs_lcnt[13]), .op(n557) );
  nand2_1 U791 ( .ip1(hcr_ic_hs_lcnt[13]), .ip2(ic_hs), .op(n556) );
  nand2_1 U792 ( .ip1(hcr_ic_ss_lcnt[13]), .ip2(ic_ss), .op(n555) );
  nand2_1 U793 ( .ip1(n570), .ip2(ic_fs_lcnt[12]), .op(n560) );
  nand2_1 U794 ( .ip1(hcr_ic_hs_lcnt[12]), .ip2(ic_hs), .op(n559) );
  nand2_1 U795 ( .ip1(hcr_ic_ss_lcnt[12]), .ip2(ic_ss), .op(n558) );
  nand2_1 U796 ( .ip1(n570), .ip2(ic_fs_lcnt[11]), .op(n563) );
  nand2_1 U797 ( .ip1(hcr_ic_hs_lcnt[11]), .ip2(ic_hs), .op(n562) );
  nand2_1 U798 ( .ip1(hcr_ic_ss_lcnt[11]), .ip2(ic_ss), .op(n561) );
  nand2_1 U799 ( .ip1(n570), .ip2(ic_fs_lcnt[10]), .op(n566) );
  nand2_1 U800 ( .ip1(hcr_ic_hs_lcnt[10]), .ip2(ic_hs), .op(n565) );
  nand2_1 U801 ( .ip1(hcr_ic_ss_lcnt[10]), .ip2(ic_ss), .op(n564) );
  nand2_1 U802 ( .ip1(n570), .ip2(ic_fs_lcnt[9]), .op(n569) );
  nand2_1 U803 ( .ip1(hcr_ic_hs_lcnt[9]), .ip2(ic_hs), .op(n568) );
  nand2_1 U804 ( .ip1(hcr_ic_ss_lcnt[9]), .ip2(ic_ss), .op(n567) );
  nand2_1 U805 ( .ip1(n570), .ip2(ic_fs_lcnt[8]), .op(n573) );
  nand2_1 U806 ( .ip1(hcr_ic_hs_lcnt[8]), .ip2(ic_hs), .op(n572) );
  nand2_1 U807 ( .ip1(hcr_ic_ss_lcnt[8]), .ip2(ic_ss), .op(n571) );
  nand2_1 U808 ( .ip1(n574), .ip2(wr_en), .op(n575) );
  mux2_1 U809 ( .ip1(ipwdata[0]), .ip2(ic_ack_general_call), .s(n575), .op(
        n1105) );
  inv_1 U810 ( .ip(ipwdata[0]), .op(n598) );
  nand2_1 U811 ( .ip1(n597), .ip2(n598), .op(n582) );
  and2_1 U812 ( .ip1(n576), .ip2(wr_en), .op(n577) );
  mux2_1 U813 ( .ip1(ic_tx_tl_0_), .ip2(n582), .s(n577), .op(n1133) );
  inv_1 U814 ( .ip(ipwdata[2]), .op(n601) );
  nand2_1 U815 ( .ip1(n597), .ip2(n601), .op(n579) );
  mux2_1 U816 ( .ip1(ic_tx_tl_2_), .ip2(n579), .s(n577), .op(n1137) );
  inv_1 U817 ( .ip(ipwdata[1]), .op(n600) );
  nand2_1 U818 ( .ip1(n597), .ip2(n600), .op(n580) );
  mux2_1 U819 ( .ip1(ic_tx_tl_1_), .ip2(n580), .s(n577), .op(n1135) );
  nand2_1 U820 ( .ip1(n578), .ip2(wr_en), .op(n581) );
  mux2_1 U821 ( .ip1(n579), .ip2(ic_rx_tl_int[2]), .s(n581), .op(n1153) );
  mux2_1 U822 ( .ip1(n580), .ip2(ic_rx_tl_int[1]), .s(n581), .op(n1151) );
  mux2_1 U823 ( .ip1(n582), .ip2(ic_rx_tl_int[0]), .s(n581), .op(n1149) );
  and2_1 U824 ( .ip1(n661), .ip2(wr_en), .op(n586) );
  mux2_1 U825 ( .ip1(ic_intr_mask[9]), .ip2(ipwdata[9]), .s(n586), .op(n1399)
         );
  mux2_1 U826 ( .ip1(ic_intr_mask[10]), .ip2(ipwdata[10]), .s(n586), .op(n1398) );
  mux2_1 U827 ( .ip1(ic_intr_mask[8]), .ip2(ipwdata[8]), .s(n586), .op(n1400)
         );
  nor3_1 U828 ( .ip1(n706), .ip2(n583), .ip3(n600), .op(n585) );
  mux2_1 U829 ( .ip1(n585), .ip2(n584), .s(ic_enable[1]), .op(n1548) );
  mux2_1 U830 ( .ip1(ic_intr_mask[11]), .ip2(ipwdata[11]), .s(n586), .op(n1397) );
  mux2_1 U831 ( .ip1(ic_intr_mask[7]), .ip2(ipwdata[7]), .s(n586), .op(n1389)
         );
  mux2_1 U832 ( .ip1(ic_intr_mask[1]), .ip2(ipwdata[1]), .s(n586), .op(n1395)
         );
  mux2_1 U833 ( .ip1(ic_intr_mask[3]), .ip2(ipwdata[3]), .s(n586), .op(n1393)
         );
  mux2_1 U834 ( .ip1(ic_intr_mask[6]), .ip2(ipwdata[6]), .s(n586), .op(n1390)
         );
  mux2_1 U835 ( .ip1(ic_intr_mask[5]), .ip2(ipwdata[5]), .s(n586), .op(n1391)
         );
  mux2_1 U836 ( .ip1(ic_intr_mask[4]), .ip2(ipwdata[4]), .s(n586), .op(n1392)
         );
  mux2_1 U837 ( .ip1(ic_intr_mask[2]), .ip2(ipwdata[2]), .s(n586), .op(n1394)
         );
  mux2_1 U838 ( .ip1(ic_intr_mask[0]), .ip2(ipwdata[0]), .s(n586), .op(n1396)
         );
  nand2_1 U839 ( .ip1(ipwdata[2]), .ip2(n600), .op(n587) );
  mux2_1 U840 ( .ip1(n587), .ip2(ic_con_pre_1_), .s(n621), .op(n1536) );
  nand2_1 U841 ( .ip1(ipwdata[1]), .ip2(n601), .op(n588) );
  mux2_1 U842 ( .ip1(n588), .ip2(ic_con_pre_2_), .s(n621), .op(n1537) );
  or2_1 U843 ( .ip1(ipwdata[3]), .ip2(n590), .op(n593) );
  mux2_1 U844 ( .ip1(n593), .ip2(ic_fs_lcnt[3]), .s(n24), .op(n1461) );
  nor2_1 U845 ( .ip1(n590), .ip2(n601), .op(n595) );
  mux2_1 U846 ( .ip1(n595), .ip2(hcr_ic_hs_lcnt[2]), .s(n589), .op(n1430) );
  nor2_1 U847 ( .ip1(n590), .ip2(n598), .op(n592) );
  mux2_1 U848 ( .ip1(n592), .ip2(hcr_ic_hs_lcnt[0]), .s(n589), .op(n1432) );
  mux2_1 U849 ( .ip1(n593), .ip2(hcr_ic_hs_lcnt[3]), .s(n589), .op(n1429) );
  nor2_1 U850 ( .ip1(n590), .ip2(n600), .op(n594) );
  mux2_1 U851 ( .ip1(n594), .ip2(hcr_ic_hs_lcnt[1]), .s(n589), .op(n1431) );
  mux2_1 U852 ( .ip1(n592), .ip2(hcr_ic_ss_lcnt[0]), .s(n591), .op(n1496) );
  mux2_1 U853 ( .ip1(n593), .ip2(hcr_ic_ss_lcnt[3]), .s(n591), .op(n1493) );
  mux2_1 U854 ( .ip1(n594), .ip2(hcr_ic_ss_lcnt[1]), .s(n591), .op(n1495) );
  mux2_1 U855 ( .ip1(n595), .ip2(hcr_ic_ss_lcnt[2]), .s(n591), .op(n1494) );
  mux2_1 U856 ( .ip1(ipwdata[9]), .ip2(ic_sda_hold[9]), .s(n629), .op(n1374)
         );
  mux2_1 U857 ( .ip1(ipwdata[10]), .ip2(ic_sda_hold[10]), .s(n629), .op(n1375)
         );
  mux2_1 U858 ( .ip1(ipwdata[14]), .ip2(ic_sda_hold[14]), .s(n629), .op(n1379)
         );
  mux2_1 U859 ( .ip1(ipwdata[12]), .ip2(ic_sda_hold[12]), .s(n596), .op(n1377)
         );
  mux2_1 U860 ( .ip1(ipwdata[15]), .ip2(ic_sda_hold[15]), .s(n629), .op(n1380)
         );
  mux2_1 U861 ( .ip1(ipwdata[13]), .ip2(ic_sda_hold[13]), .s(n596), .op(n1378)
         );
  mux2_1 U862 ( .ip1(ipwdata[11]), .ip2(ic_sda_hold[11]), .s(n629), .op(n1376)
         );
  nand3_1 U863 ( .ip1(n601), .ip2(n597), .ip3(n600), .op(n599) );
  nand2_1 U864 ( .ip1(n599), .ip2(n598), .op(n626) );
  mux2_1 U865 ( .ip1(n626), .ip2(ic_hs_spklen[0]), .s(n624), .op(n1401) );
  nand2_1 U866 ( .ip1(n602), .ip2(n600), .op(n604) );
  mux2_1 U867 ( .ip1(n604), .ip2(hcr_ic_ss_hcnt[1]), .s(n603), .op(n1511) );
  nand2_1 U868 ( .ip1(n602), .ip2(n601), .op(n631) );
  mux2_1 U869 ( .ip1(n631), .ip2(hcr_ic_ss_hcnt[2]), .s(n603), .op(n1510) );
  mux2_1 U870 ( .ip1(ipwdata[6]), .ip2(hcr_ic_ss_hcnt[6]), .s(n603), .op(n1506) );
  mux2_1 U871 ( .ip1(ipwdata[5]), .ip2(hcr_ic_ss_hcnt[5]), .s(n603), .op(n1507) );
  mux2_1 U872 ( .ip1(n604), .ip2(ic_fs_hcnt[1]), .s(n605), .op(n1479) );
  mux2_1 U873 ( .ip1(ipwdata[6]), .ip2(ic_fs_hcnt[6]), .s(n605), .op(n1474) );
  mux2_1 U874 ( .ip1(n604), .ip2(hcr_ic_hs_hcnt[1]), .s(n630), .op(n1447) );
  mux2_1 U875 ( .ip1(n631), .ip2(ic_fs_hcnt[2]), .s(n605), .op(n1478) );
  mux2_1 U876 ( .ip1(ipwdata[5]), .ip2(ic_fs_hcnt[5]), .s(n605), .op(n1475) );
  inv_1 U877 ( .ip(ic_txflr[0]), .op(n694) );
  mux2_1 U878 ( .ip1(n607), .ip2(n606), .s(n694), .op(n1363) );
  mux2_1 U879 ( .ip1(n610), .ip2(n693), .s(n694), .op(n613) );
  or2_1 U880 ( .ip1(n693), .ip2(n607), .op(n609) );
  or2_1 U881 ( .ip1(ic_txflr[0]), .ip2(n607), .op(n608) );
  nand2_1 U882 ( .ip1(n609), .ip2(n608), .op(n684) );
  nand2_1 U883 ( .ip1(n610), .ip2(n694), .op(n611) );
  nand2_1 U884 ( .ip1(n684), .ip2(n611), .op(n612) );
  mux2_1 U885 ( .ip1(n613), .ip2(n612), .s(ic_txflr[1]), .op(n1362) );
  nor3_1 U886 ( .ip1(ic_rxflr[0]), .ip2(ic_rxflr[1]), .ip3(n614), .op(n682) );
  or2_1 U887 ( .ip1(n615), .ip2(n682), .op(n618) );
  inv_1 U888 ( .ip(n616), .op(n617) );
  mux2_1 U889 ( .ip1(n618), .ip2(n617), .s(ic_rxflr[2]), .op(n1544) );
  mux2_1 U890 ( .ip1(ipwdata[8]), .ip2(tx_empty_ctrl), .s(n621), .op(n1543) );
  mux2_1 U891 ( .ip1(ipwdata[7]), .ip2(p_det_ifaddr), .s(n621), .op(n1542) );
  mux2_1 U892 ( .ip1(ipwdata[1]), .ip2(ic_hs_maddr[1]), .s(n623), .op(n1165)
         );
  mux2_1 U893 ( .ip1(ipwdata[2]), .ip2(ic_hs_maddr[2]), .s(n623), .op(n1167)
         );
  mux2_1 U894 ( .ip1(ipwdata[9]), .ip2(ic_sar[9]), .s(n620), .op(n1533) );
  mux2_1 U895 ( .ip1(ipwdata[8]), .ip2(ic_sar[8]), .s(n620), .op(n1534) );
  mux2_1 U896 ( .ip1(ipwdata[6]), .ip2(ic_con_pre_6_), .s(n621), .op(n1541) );
  mux2_1 U897 ( .ip1(ipwdata[5]), .ip2(ic_rstrt_en), .s(n621), .op(n1540) );
  mux2_1 U898 ( .ip1(ipwdata[4]), .ip2(ic_10bit_mst), .s(n621), .op(n1539) );
  mux2_1 U899 ( .ip1(ipwdata[3]), .ip2(ic_10bit_slv), .s(n621), .op(n1538) );
  mux2_1 U900 ( .ip1(ipwdata[0]), .ip2(ic_master), .s(n621), .op(n1535) );
  mux2_1 U901 ( .ip1(ipwdata[3]), .ip2(ic_sar[3]), .s(n620), .op(n1525) );
  mux2_1 U902 ( .ip1(ipwdata[5]), .ip2(ic_sar[5]), .s(n620), .op(n1523) );
  mux2_1 U903 ( .ip1(ipwdata[7]), .ip2(ic_sar[7]), .s(n620), .op(n1521) );
  mux2_1 U904 ( .ip1(ipwdata[1]), .ip2(ic_sar[1]), .s(n620), .op(n1527) );
  mux2_1 U905 ( .ip1(ipwdata[11]), .ip2(ic_tar[11]), .s(n622), .op(n1529) );
  mux2_1 U906 ( .ip1(ipwdata[10]), .ip2(ic_tar[10]), .s(n622), .op(n1530) );
  mux2_1 U907 ( .ip1(ipwdata[9]), .ip2(ic_tar[9]), .s(n622), .op(n1531) );
  mux2_1 U908 ( .ip1(ipwdata[8]), .ip2(ic_tar[8]), .s(n622), .op(n1532) );
  mux2_1 U909 ( .ip1(ipwdata[7]), .ip2(ic_tar[7]), .s(n622), .op(n1513) );
  mux2_1 U910 ( .ip1(ipwdata[3]), .ip2(ic_tar[3]), .s(n622), .op(n1517) );
  mux2_1 U911 ( .ip1(ipwdata[1]), .ip2(ic_tar[1]), .s(n622), .op(n1519) );
  mux2_1 U912 ( .ip1(ipwdata[5]), .ip2(ic_tar[5]), .s(n622), .op(n1515) );
  mux2_1 U913 ( .ip1(ipwdata[0]), .ip2(ic_hs_maddr[0]), .s(n623), .op(n1113)
         );
  mux2_1 U914 ( .ip1(ipwdata[12]), .ip2(ic_fs_lcnt[12]), .s(n24), .op(n1451)
         );
  mux2_1 U915 ( .ip1(ipwdata[14]), .ip2(ic_fs_lcnt[14]), .s(n24), .op(n1449)
         );
  mux2_1 U916 ( .ip1(ipwdata[13]), .ip2(ic_fs_lcnt[13]), .s(n24), .op(n1450)
         );
  mux2_1 U917 ( .ip1(ipwdata[15]), .ip2(ic_fs_lcnt[15]), .s(n24), .op(n1456)
         );
  mux2_1 U918 ( .ip1(ipwdata[10]), .ip2(ic_fs_lcnt[10]), .s(n24), .op(n1453)
         );
  mux2_1 U919 ( .ip1(ipwdata[11]), .ip2(ic_fs_lcnt[11]), .s(n24), .op(n1452)
         );
  mux2_1 U920 ( .ip1(ipwdata[9]), .ip2(ic_fs_lcnt[9]), .s(n24), .op(n1454) );
  mux2_1 U921 ( .ip1(ipwdata[8]), .ip2(ic_fs_lcnt[8]), .s(n24), .op(n1455) );
  mux2_1 U922 ( .ip1(ipwdata[6]), .ip2(ic_fs_lcnt[6]), .s(n24), .op(n1458) );
  mux2_1 U923 ( .ip1(ipwdata[5]), .ip2(ic_fs_lcnt[5]), .s(n24), .op(n1459) );
  mux2_1 U924 ( .ip1(ipwdata[4]), .ip2(ic_fs_lcnt[4]), .s(n24), .op(n1460) );
  mux2_1 U925 ( .ip1(ipwdata[14]), .ip2(hcr_ic_hs_lcnt[14]), .s(n589), .op(
        n1417) );
  mux2_1 U926 ( .ip1(ipwdata[13]), .ip2(hcr_ic_hs_lcnt[13]), .s(n589), .op(
        n1418) );
  mux2_1 U927 ( .ip1(ipwdata[15]), .ip2(hcr_ic_hs_lcnt[15]), .s(n589), .op(
        n1424) );
  mux2_1 U928 ( .ip1(ipwdata[12]), .ip2(hcr_ic_hs_lcnt[12]), .s(n589), .op(
        n1419) );
  mux2_1 U929 ( .ip1(ipwdata[9]), .ip2(hcr_ic_hs_lcnt[9]), .s(n589), .op(n1422) );
  mux2_1 U930 ( .ip1(ipwdata[11]), .ip2(hcr_ic_hs_lcnt[11]), .s(n589), .op(
        n1420) );
  mux2_1 U931 ( .ip1(ipwdata[10]), .ip2(hcr_ic_hs_lcnt[10]), .s(n589), .op(
        n1421) );
  mux2_1 U932 ( .ip1(ipwdata[8]), .ip2(hcr_ic_hs_lcnt[8]), .s(n589), .op(n1423) );
  mux2_1 U933 ( .ip1(ipwdata[6]), .ip2(hcr_ic_hs_lcnt[6]), .s(n589), .op(n1426) );
  mux2_1 U934 ( .ip1(ipwdata[5]), .ip2(hcr_ic_hs_lcnt[5]), .s(n589), .op(n1427) );
  mux2_1 U935 ( .ip1(ipwdata[7]), .ip2(hcr_ic_hs_lcnt[7]), .s(n589), .op(n1425) );
  mux2_1 U936 ( .ip1(ipwdata[15]), .ip2(hcr_ic_ss_lcnt[15]), .s(n591), .op(
        n1488) );
  mux2_1 U937 ( .ip1(ipwdata[12]), .ip2(hcr_ic_ss_lcnt[12]), .s(n591), .op(
        n1483) );
  mux2_1 U938 ( .ip1(ipwdata[14]), .ip2(hcr_ic_ss_lcnt[14]), .s(n591), .op(
        n1481) );
  mux2_1 U939 ( .ip1(ipwdata[13]), .ip2(hcr_ic_ss_lcnt[13]), .s(n591), .op(
        n1482) );
  mux2_1 U940 ( .ip1(ipwdata[9]), .ip2(hcr_ic_ss_lcnt[9]), .s(n591), .op(n1486) );
  mux2_1 U941 ( .ip1(ipwdata[11]), .ip2(hcr_ic_ss_lcnt[11]), .s(n591), .op(
        n1484) );
  mux2_1 U942 ( .ip1(ipwdata[10]), .ip2(hcr_ic_ss_lcnt[10]), .s(n591), .op(
        n1485) );
  mux2_1 U943 ( .ip1(ipwdata[5]), .ip2(hcr_ic_ss_lcnt[5]), .s(n591), .op(n1491) );
  mux2_1 U944 ( .ip1(ipwdata[6]), .ip2(ic_sar[6]), .s(n620), .op(n1522) );
  mux2_1 U945 ( .ip1(ipwdata[4]), .ip2(ic_sar[4]), .s(n620), .op(n1524) );
  mux2_1 U946 ( .ip1(ipwdata[2]), .ip2(ic_sar[2]), .s(n620), .op(n1526) );
  mux2_1 U947 ( .ip1(ipwdata[0]), .ip2(ic_sar[0]), .s(n620), .op(n1528) );
  mux2_1 U948 ( .ip1(ipwdata[4]), .ip2(ic_tar[4]), .s(n622), .op(n1516) );
  mux2_1 U949 ( .ip1(ipwdata[6]), .ip2(ic_tar[6]), .s(n622), .op(n1514) );
  mux2_1 U950 ( .ip1(ipwdata[2]), .ip2(ic_tar[2]), .s(n622), .op(n1518) );
  mux2_1 U951 ( .ip1(ipwdata[0]), .ip2(ic_tar[0]), .s(n622), .op(n1520) );
  mux2_1 U952 ( .ip1(ipwdata[7]), .ip2(ic_fs_lcnt[7]), .s(n24), .op(n1457) );
  mux2_1 U953 ( .ip1(ipwdata[4]), .ip2(hcr_ic_hs_lcnt[4]), .s(n589), .op(n1428) );
  mux2_1 U954 ( .ip1(ipwdata[8]), .ip2(hcr_ic_ss_lcnt[8]), .s(n591), .op(n1487) );
  mux2_1 U955 ( .ip1(ipwdata[7]), .ip2(hcr_ic_ss_lcnt[7]), .s(n591), .op(n1489) );
  mux2_1 U956 ( .ip1(ipwdata[4]), .ip2(hcr_ic_ss_lcnt[4]), .s(n591), .op(n1492) );
  mux2_1 U957 ( .ip1(ipwdata[6]), .ip2(hcr_ic_ss_lcnt[6]), .s(n591), .op(n1490) );
  mux2_1 U958 ( .ip1(ipwdata[3]), .ip2(ic_fs_spklen[3]), .s(n627), .op(n1412)
         );
  mux2_1 U959 ( .ip1(ipwdata[7]), .ip2(ic_fs_spklen[7]), .s(n627), .op(n1416)
         );
  mux2_1 U960 ( .ip1(ipwdata[6]), .ip2(ic_fs_spklen[6]), .s(n627), .op(n1415)
         );
  mux2_1 U961 ( .ip1(ipwdata[7]), .ip2(ic_hs_spklen[7]), .s(n624), .op(n1408)
         );
  mux2_1 U962 ( .ip1(ipwdata[4]), .ip2(ic_fs_spklen[4]), .s(n627), .op(n1413)
         );
  mux2_1 U963 ( .ip1(ipwdata[6]), .ip2(ic_hs_spklen[6]), .s(n624), .op(n1407)
         );
  mux2_1 U964 ( .ip1(ipwdata[3]), .ip2(ic_hs_spklen[3]), .s(n624), .op(n1404)
         );
  mux2_1 U965 ( .ip1(ipwdata[4]), .ip2(ic_hs_spklen[4]), .s(n624), .op(n1405)
         );
  mux2_1 U966 ( .ip1(ipwdata[1]), .ip2(ic_fs_spklen[1]), .s(n627), .op(n1410)
         );
  mux2_1 U967 ( .ip1(ipwdata[5]), .ip2(ic_fs_spklen[5]), .s(n627), .op(n1414)
         );
  mux2_1 U968 ( .ip1(ipwdata[5]), .ip2(ic_hs_spklen[5]), .s(n624), .op(n1406)
         );
  mux2_1 U969 ( .ip1(ipwdata[1]), .ip2(ic_hs_spklen[1]), .s(n624), .op(n1402)
         );
  mux2_1 U970 ( .ip1(ipwdata[2]), .ip2(ic_hs_spklen[2]), .s(n624), .op(n1403)
         );
  mux2_1 U971 ( .ip1(ipwdata[7]), .ip2(ic_sda_setup[7]), .s(n628), .op(n1131)
         );
  mux2_1 U972 ( .ip1(ipwdata[1]), .ip2(ic_sda_setup[1]), .s(n628), .op(n1125)
         );
  mux2_1 U973 ( .ip1(ipwdata[4]), .ip2(ic_sda_setup[4]), .s(n628), .op(n1129)
         );
  mux2_1 U974 ( .ip1(ipwdata[3]), .ip2(ic_sda_setup[3]), .s(n628), .op(n1127)
         );
  mux2_1 U975 ( .ip1(ipwdata[0]), .ip2(ic_sda_setup[0]), .s(n628), .op(n1123)
         );
  mux2_1 U976 ( .ip1(ipwdata[8]), .ip2(ic_sda_hold[8]), .s(n629), .op(n1373)
         );
  mux2_1 U977 ( .ip1(ipwdata[3]), .ip2(ic_sda_hold[3]), .s(n629), .op(n1368)
         );
  mux2_1 U978 ( .ip1(ipwdata[6]), .ip2(ic_sda_hold[6]), .s(n629), .op(n1371)
         );
  mux2_1 U979 ( .ip1(ipwdata[7]), .ip2(ic_sda_hold[7]), .s(n629), .op(n1372)
         );
  mux2_1 U980 ( .ip1(ipwdata[1]), .ip2(ic_sda_hold[1]), .s(n629), .op(n1366)
         );
  mux2_1 U981 ( .ip1(ipwdata[5]), .ip2(ic_sda_hold[5]), .s(n629), .op(n1370)
         );
  mux2_1 U982 ( .ip1(ipwdata[4]), .ip2(ic_sda_hold[4]), .s(n629), .op(n1369)
         );
  mux2_1 U983 ( .ip1(ipwdata[2]), .ip2(ic_sda_hold[2]), .s(n629), .op(n1367)
         );
  mux2_1 U984 ( .ip1(ipwdata[20]), .ip2(ic_sda_hold[20]), .s(n596), .op(n1385)
         );
  mux2_1 U985 ( .ip1(ipwdata[19]), .ip2(ic_sda_hold[19]), .s(n596), .op(n1384)
         );
  mux2_1 U986 ( .ip1(ipwdata[23]), .ip2(ic_sda_hold[23]), .s(n596), .op(n1388)
         );
  mux2_1 U987 ( .ip1(ipwdata[21]), .ip2(ic_sda_hold[21]), .s(n596), .op(n1386)
         );
  mux2_1 U988 ( .ip1(ipwdata[16]), .ip2(ic_sda_hold[16]), .s(n596), .op(n1381)
         );
  mux2_1 U989 ( .ip1(ipwdata[17]), .ip2(ic_sda_hold[17]), .s(n596), .op(n1382)
         );
  mux2_1 U990 ( .ip1(ipwdata[18]), .ip2(ic_sda_hold[18]), .s(n596), .op(n1383)
         );
  mux2_1 U991 ( .ip1(ipwdata[22]), .ip2(ic_sda_hold[22]), .s(n596), .op(n1387)
         );
  mux2_1 U992 ( .ip1(n626), .ip2(ic_fs_spklen[0]), .s(n627), .op(n1409) );
  mux2_1 U993 ( .ip1(ipwdata[2]), .ip2(ic_fs_spklen[2]), .s(n627), .op(n1411)
         );
  mux2_1 U994 ( .ip1(ipwdata[6]), .ip2(ic_sda_setup[6]), .s(n628), .op(n1111)
         );
  mux2_1 U995 ( .ip1(ipwdata[5]), .ip2(ic_sda_setup[5]), .s(n628), .op(n1109)
         );
  mux2_1 U996 ( .ip1(ipwdata[2]), .ip2(ic_sda_setup[2]), .s(n628), .op(n1107)
         );
  mux2_1 U997 ( .ip1(ipwdata[0]), .ip2(ic_sda_hold[0]), .s(n629), .op(n1365)
         );
  mux2_1 U998 ( .ip1(ipwdata[6]), .ip2(hcr_ic_hs_hcnt[6]), .s(n630), .op(n1442) );
  mux2_1 U999 ( .ip1(ipwdata[5]), .ip2(hcr_ic_hs_hcnt[5]), .s(n630), .op(n1443) );
  mux2_1 U1000 ( .ip1(n631), .ip2(hcr_ic_hs_hcnt[2]), .s(n630), .op(n1446) );
  nand2_1 U1001 ( .ip1(n632), .ip2(ic_fs_hcnt[3]), .op(n636) );
  nand2_1 U1002 ( .ip1(n633), .ip2(hcr_ic_ss_lcnt[3]), .op(n635) );
  nand2_1 U1003 ( .ip1(n677), .ip2(ic_sda_hold[3]), .op(n634) );
  nand3_1 U1004 ( .ip1(n636), .ip2(n635), .ip3(n634), .op(n675) );
  nor2_1 U1005 ( .ip1(rx_empty), .ip2(n637), .op(n647) );
  nand2_1 U1006 ( .ip1(ic_raw_intr_stat[3]), .ip2(n638), .op(n645) );
  nand2_1 U1007 ( .ip1(n639), .ip2(ic_rxflr[3]), .op(n644) );
  nand2_1 U1008 ( .ip1(n640), .ip2(ic_txflr[3]), .op(n643) );
  nand2_1 U1009 ( .ip1(n641), .ip2(hcr_ic_ss_hcnt[3]), .op(n642) );
  nand4_1 U1010 ( .ip1(n645), .ip2(n644), .ip3(n643), .ip4(n642), .op(n646) );
  not_ab_or_c_or_d U1011 ( .ip1(hcr_ic_hs_lcnt[3]), .ip2(n648), .ip3(n647), 
        .ip4(n646), .op(n673) );
  nand2_1 U1012 ( .ip1(n649), .ip2(ic_tar[3]), .op(n656) );
  nand2_1 U1013 ( .ip1(n650), .ip2(ic_fs_spklen[3]), .op(n655) );
  nand2_1 U1014 ( .ip1(n651), .ip2(ic_10bit_slv), .op(n654) );
  nand2_1 U1015 ( .ip1(n652), .ip2(ic_fs_lcnt[3]), .op(n653) );
  nand4_1 U1016 ( .ip1(n656), .ip2(n655), .ip3(n654), .ip4(n653), .op(n667) );
  not_ab_or_c_or_d U1017 ( .ip1(n658), .ip2(ic_intr_stat[3]), .ip3(iprdata[29]), .ip4(n657), .op(n665) );
  nand2_1 U1018 ( .ip1(n659), .ip2(hcr_ic_hs_hcnt[3]), .op(n664) );
  nand2_1 U1019 ( .ip1(n660), .ip2(ic_sda_setup[3]), .op(n663) );
  nand2_1 U1020 ( .ip1(n661), .ip2(ic_intr_mask[3]), .op(n662) );
  nand4_1 U1021 ( .ip1(n665), .ip2(n664), .ip3(n663), .ip4(n662), .op(n666) );
  not_ab_or_c_or_d U1022 ( .ip1(n678), .ip2(ic_tx_abrt_source[3]), .ip3(n667), 
        .ip4(n666), .op(n672) );
  nand2_1 U1023 ( .ip1(n668), .ip2(rx_pop_data[3]), .op(n671) );
  nand2_1 U1024 ( .ip1(n669), .ip2(ic_sar[3]), .op(n670) );
  nand4_1 U1025 ( .ip1(n673), .ip2(n672), .ip3(n671), .ip4(n670), .op(n674) );
  ab_or_c_or_d U1026 ( .ip1(n676), .ip2(ic_hs_spklen[3]), .ip3(n675), .ip4(
        n674), .op(iprdata[3]) );
  inv_1 U1027 ( .ip(ic_con_pre_6_), .op(ic_slave_en) );
  and2_1 U1028 ( .ip1(n677), .ip2(ic_sda_hold[19]), .op(iprdata[19]) );
  and2_1 U1029 ( .ip1(n678), .ip2(ic_txflr_flushed[2]), .op(iprdata[25]) );
  nor2_1 U1030 ( .ip1(ic_con_pre_1_), .ip2(n679), .op(ic_fs) );
  nor2_1 U1031 ( .ip1(ic_rxflr[1]), .ip2(n680), .op(n681) );
  ab_or_c_or_d U1032 ( .ip1(ic_rxflr[1]), .ip2(n683), .ip3(n682), .ip4(n681), 
        .op(n1545) );
  inv_1 U1033 ( .ip(ic_txflr[2]), .op(n705) );
  or2_1 U1034 ( .ip1(n684), .ip2(n705), .op(n687) );
  nand2_1 U1035 ( .ip1(ic_txflr[1]), .ip2(n693), .op(n685) );
  or2_1 U1036 ( .ip1(n685), .ip2(n705), .op(n686) );
  nand2_1 U1037 ( .ip1(n687), .ip2(n686), .op(n691) );
  nand2_1 U1038 ( .ip1(ic_txflr[0]), .ip2(ic_txflr[1]), .op(n688) );
  mux2_1 U1039 ( .ip1(ic_txflr[2]), .ip2(n705), .s(n688), .op(n704) );
  nor2_1 U1040 ( .ip1(n689), .ip2(n704), .op(n690) );
  ab_or_c_or_d U1041 ( .ip1(n693), .ip2(n692), .ip3(n691), .ip4(n690), .op(
        n1361) );
  mux2_1 U1042 ( .ip1(n694), .ip2(ic_txflr[0]), .s(abrt_in_rcve_trns), .op(
        n696) );
  nor2_1 U1043 ( .ip1(ic_txflr_flushed[0]), .ip2(tx_abrt_flg_edg), .op(n695)
         );
  not_ab_or_c_or_d U1044 ( .ip1(tx_abrt_flg_edg), .ip2(n696), .ip3(n695), 
        .ip4(n706), .op(n1121) );
  nand2_1 U1045 ( .ip1(abrt_in_rcve_trns), .ip2(ic_txflr[0]), .op(n697) );
  xor2_1 U1046 ( .ip1(ic_txflr[1]), .ip2(n697), .op(n699) );
  nor2_1 U1047 ( .ip1(ic_txflr_flushed[1]), .ip2(tx_abrt_flg_edg), .op(n698)
         );
  not_ab_or_c_or_d U1048 ( .ip1(tx_abrt_flg_edg), .ip2(n699), .ip3(n698), 
        .ip4(n706), .op(n1119) );
  mux2_1 U1049 ( .ip1(n701), .ip2(n700), .s(abrt_in_rcve_trns), .op(n703) );
  nor2_1 U1050 ( .ip1(ic_txflr_flushed[3]), .ip2(tx_abrt_flg_edg), .op(n702)
         );
  not_ab_or_c_or_d U1051 ( .ip1(tx_abrt_flg_edg), .ip2(n703), .ip3(n702), 
        .ip4(n706), .op(n1117) );
  mux2_1 U1052 ( .ip1(n705), .ip2(n704), .s(abrt_in_rcve_trns), .op(n708) );
  nor2_1 U1053 ( .ip1(ic_txflr_flushed[2]), .ip2(tx_abrt_flg_edg), .op(n707)
         );
  not_ab_or_c_or_d U1054 ( .ip1(tx_abrt_flg_edg), .ip2(n708), .ip3(n707), 
        .ip4(n706), .op(n1115) );
endmodule


module interconnect_ip ( HCLK_hclk, HRESETn_hresetn, PCLK_pclk, 
        PRESETn_presetn, ex_i_ahb_AHB_MASTER_CORTEXM0_haddr, 
        ex_i_ahb_AHB_MASTER_CORTEXM0_hburst, 
        ex_i_ahb_AHB_MASTER_CORTEXM0_hlock, ex_i_ahb_AHB_MASTER_CORTEXM0_hprot, 
        ex_i_ahb_AHB_MASTER_CORTEXM0_hsize, 
        ex_i_ahb_AHB_MASTER_CORTEXM0_htrans, 
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata, 
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite, 
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata, 
        ex_i_ahb_AHB_MASTER_CORTEXM0_hready, 
        ex_i_ahb_AHB_MASTER_CORTEXM0_hresp, ex_i_ahb_AHB_Slave_PID_hrdata, 
        ex_i_ahb_AHB_Slave_PID_hready_resp, ex_i_ahb_AHB_Slave_PID_hresp, 
        ex_i_ahb_AHB_Slave_PID_haddr, ex_i_ahb_AHB_Slave_PID_hburst, 
        ex_i_ahb_AHB_Slave_PID_hmastlock, ex_i_ahb_AHB_Slave_PID_hprot, 
        ex_i_ahb_AHB_Slave_PID_hready, ex_i_ahb_AHB_Slave_PID_hsel, 
        ex_i_ahb_AHB_Slave_PID_hsize, ex_i_ahb_AHB_Slave_PID_htrans, 
        ex_i_ahb_AHB_Slave_PID_hwdata, ex_i_ahb_AHB_Slave_PID_hwrite, 
        ex_i_ahb_AHB_Slave_PWM_hrdata, ex_i_ahb_AHB_Slave_PWM_hready_resp, 
        ex_i_ahb_AHB_Slave_PWM_hresp, ex_i_ahb_AHB_Slave_PWM_haddr, 
        ex_i_ahb_AHB_Slave_PWM_hburst, ex_i_ahb_AHB_Slave_PWM_hmastlock, 
        ex_i_ahb_AHB_Slave_PWM_hprot, ex_i_ahb_AHB_Slave_PWM_hready, 
        ex_i_ahb_AHB_Slave_PWM_hsel, ex_i_ahb_AHB_Slave_PWM_hsize, 
        ex_i_ahb_AHB_Slave_PWM_htrans, ex_i_ahb_AHB_Slave_PWM_hwdata, 
        ex_i_ahb_AHB_Slave_PWM_hwrite, ex_i_ahb_AHB_Slave_RAM_hrdata, 
        ex_i_ahb_AHB_Slave_RAM_hready_resp, ex_i_ahb_AHB_Slave_RAM_hresp, 
        ex_i_ahb_AHB_Slave_RAM_haddr, ex_i_ahb_AHB_Slave_RAM_hburst, 
        ex_i_ahb_AHB_Slave_RAM_hmastlock, ex_i_ahb_AHB_Slave_RAM_hprot, 
        ex_i_ahb_AHB_Slave_RAM_hready, ex_i_ahb_AHB_Slave_RAM_hsel, 
        ex_i_ahb_AHB_Slave_RAM_hsize, ex_i_ahb_AHB_Slave_RAM_htrans, 
        ex_i_ahb_AHB_Slave_RAM_hwdata, ex_i_ahb_AHB_Slave_RAM_hwrite, 
        i_apb_pclk_en, i_i2c_ic_clk, i_i2c_ic_clk_in_a, i_i2c_ic_data_in_a, 
        i_i2c_ic_rst_n, i_ssi_rxd, i_ssi_ss_in_n, i_ssi_ssi_clk, 
        i_ssi_ssi_rst_n, i_ahb_hmaster_data, i_i2c_debug_addr, 
        i_i2c_debug_addr_10bit, i_i2c_debug_data, i_i2c_debug_hs, 
        i_i2c_debug_master_act, i_i2c_debug_mst_cstate, i_i2c_debug_p_gen, 
        i_i2c_debug_rd, i_i2c_debug_s_gen, i_i2c_debug_slave_act, 
        i_i2c_debug_slv_cstate, i_i2c_debug_wr, i_i2c_ic_activity_intr, 
        i_i2c_ic_clk_oe, i_i2c_ic_current_src_en, i_i2c_ic_data_oe, 
        i_i2c_ic_en, i_i2c_ic_gen_call_intr, i_i2c_ic_rd_req_intr, 
        i_i2c_ic_rx_done_intr, i_i2c_ic_rx_full_intr, i_i2c_ic_rx_over_intr, 
        i_i2c_ic_rx_under_intr, i_i2c_ic_start_det_intr, 
        i_i2c_ic_stop_det_intr, i_i2c_ic_tx_abrt_intr, i_i2c_ic_tx_empty_intr, 
        i_i2c_ic_tx_over_intr, i_ssi_sclk_out, i_ssi_ss_0_n, 
        i_ssi_ssi_mst_intr_n, i_ssi_ssi_oe_n, i_ssi_ssi_rxf_intr_n, 
        i_ssi_ssi_rxo_intr_n, i_ssi_ssi_rxu_intr_n, i_ssi_ssi_sleep, 
        i_ssi_ssi_txe_intr_n, i_ssi_ssi_txo_intr_n, i_ssi_txd );
  input [31:0] ex_i_ahb_AHB_MASTER_CORTEXM0_haddr;
  input [2:0] ex_i_ahb_AHB_MASTER_CORTEXM0_hburst;
  input [3:0] ex_i_ahb_AHB_MASTER_CORTEXM0_hprot;
  input [2:0] ex_i_ahb_AHB_MASTER_CORTEXM0_hsize;
  input [1:0] ex_i_ahb_AHB_MASTER_CORTEXM0_htrans;
  input [31:0] ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata;
  output [31:0] ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata;
  output [1:0] ex_i_ahb_AHB_MASTER_CORTEXM0_hresp;
  input [31:0] ex_i_ahb_AHB_Slave_PID_hrdata;
  input [1:0] ex_i_ahb_AHB_Slave_PID_hresp;
  output [31:0] ex_i_ahb_AHB_Slave_PID_haddr;
  output [2:0] ex_i_ahb_AHB_Slave_PID_hburst;
  output [3:0] ex_i_ahb_AHB_Slave_PID_hprot;
  output [2:0] ex_i_ahb_AHB_Slave_PID_hsize;
  output [1:0] ex_i_ahb_AHB_Slave_PID_htrans;
  output [31:0] ex_i_ahb_AHB_Slave_PID_hwdata;
  input [31:0] ex_i_ahb_AHB_Slave_PWM_hrdata;
  input [1:0] ex_i_ahb_AHB_Slave_PWM_hresp;
  output [31:0] ex_i_ahb_AHB_Slave_PWM_haddr;
  output [2:0] ex_i_ahb_AHB_Slave_PWM_hburst;
  output [3:0] ex_i_ahb_AHB_Slave_PWM_hprot;
  output [2:0] ex_i_ahb_AHB_Slave_PWM_hsize;
  output [1:0] ex_i_ahb_AHB_Slave_PWM_htrans;
  output [31:0] ex_i_ahb_AHB_Slave_PWM_hwdata;
  input [31:0] ex_i_ahb_AHB_Slave_RAM_hrdata;
  input [1:0] ex_i_ahb_AHB_Slave_RAM_hresp;
  output [31:0] ex_i_ahb_AHB_Slave_RAM_haddr;
  output [2:0] ex_i_ahb_AHB_Slave_RAM_hburst;
  output [3:0] ex_i_ahb_AHB_Slave_RAM_hprot;
  output [2:0] ex_i_ahb_AHB_Slave_RAM_hsize;
  output [1:0] ex_i_ahb_AHB_Slave_RAM_htrans;
  output [31:0] ex_i_ahb_AHB_Slave_RAM_hwdata;
  output [3:0] i_ahb_hmaster_data;
  output [4:0] i_i2c_debug_mst_cstate;
  output [3:0] i_i2c_debug_slv_cstate;
  input HCLK_hclk, HRESETn_hresetn, PCLK_pclk, PRESETn_presetn,
         ex_i_ahb_AHB_MASTER_CORTEXM0_hlock,
         ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite,
         ex_i_ahb_AHB_Slave_PID_hready_resp,
         ex_i_ahb_AHB_Slave_PWM_hready_resp,
         ex_i_ahb_AHB_Slave_RAM_hready_resp, i_apb_pclk_en, i_i2c_ic_clk,
         i_i2c_ic_clk_in_a, i_i2c_ic_data_in_a, i_i2c_ic_rst_n, i_ssi_rxd,
         i_ssi_ss_in_n, i_ssi_ssi_clk, i_ssi_ssi_rst_n;
  output ex_i_ahb_AHB_MASTER_CORTEXM0_hready, ex_i_ahb_AHB_Slave_PID_hmastlock,
         ex_i_ahb_AHB_Slave_PID_hready, ex_i_ahb_AHB_Slave_PID_hsel,
         ex_i_ahb_AHB_Slave_PID_hwrite, ex_i_ahb_AHB_Slave_PWM_hmastlock,
         ex_i_ahb_AHB_Slave_PWM_hready, ex_i_ahb_AHB_Slave_PWM_hsel,
         ex_i_ahb_AHB_Slave_PWM_hwrite, ex_i_ahb_AHB_Slave_RAM_hmastlock,
         ex_i_ahb_AHB_Slave_RAM_hready, ex_i_ahb_AHB_Slave_RAM_hsel,
         ex_i_ahb_AHB_Slave_RAM_hwrite, i_i2c_debug_addr,
         i_i2c_debug_addr_10bit, i_i2c_debug_data, i_i2c_debug_hs,
         i_i2c_debug_master_act, i_i2c_debug_p_gen, i_i2c_debug_rd,
         i_i2c_debug_s_gen, i_i2c_debug_slave_act, i_i2c_debug_wr,
         i_i2c_ic_activity_intr, i_i2c_ic_clk_oe, i_i2c_ic_current_src_en,
         i_i2c_ic_data_oe, i_i2c_ic_en, i_i2c_ic_gen_call_intr,
         i_i2c_ic_rd_req_intr, i_i2c_ic_rx_done_intr, i_i2c_ic_rx_full_intr,
         i_i2c_ic_rx_over_intr, i_i2c_ic_rx_under_intr,
         i_i2c_ic_start_det_intr, i_i2c_ic_stop_det_intr,
         i_i2c_ic_tx_abrt_intr, i_i2c_ic_tx_empty_intr, i_i2c_ic_tx_over_intr,
         i_ssi_sclk_out, i_ssi_ss_0_n, i_ssi_ssi_mst_intr_n, i_ssi_ssi_oe_n,
         i_ssi_ssi_rxf_intr_n, i_ssi_ssi_rxo_intr_n, i_ssi_ssi_rxu_intr_n,
         i_ssi_ssi_sleep, i_ssi_ssi_txe_intr_n, i_ssi_ssi_txo_intr_n,
         i_ssi_txd;
  wire   ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite, ex_i_ahb_AHB_Slave_PID_hmastlock,
         i_apb_hready_resp, i_apb_penable, i_apb_pwrite, i_ahb_hresp_none_0_,
         i_apb_psel_en, i_i2c_tx_full, i_i2c_rx_full, i_i2c_tx_push,
         i_i2c_rx_pop, i_i2c_rx_push_sync, i_i2c_tx_pop_sync,
         i_i2c_tx_fifo_rst_n, i_i2c_fifo_rst_n, i_i2c_abrt_in_rcve_trns,
         i_i2c_split_start_en, i_i2c_ack_det, i_i2c_ic_bus_idle,
         i_i2c_slv_addressed, i_i2c_slv_ack_det, i_i2c_p_det, i_i2c_wr_en,
         i_i2c_sda_vld, i_i2c_sda_int, i_i2c_slv_rx_2addr, i_i2c_rx_hs_mcode,
         i_i2c_rx_addr_match, i_i2c_slv_rxbyte_rdy, i_i2c_rx_slv_read,
         i_i2c_mst_rxbyte_rdy, i_i2c_slv_rx_ack_vld, i_i2c_mst_rx_bwen,
         i_i2c_rx_scl_hcnt_en, i_i2c_rx_scl_lcnt_en, i_i2c_mst_rx_data_scl,
         i_i2c_mst_rx_ack_vld, i_i2c_slv_tx_ack_vld, i_i2c_mst_tx_ack_vld,
         i_i2c_scl_p_setup_cmplt, i_i2c_scl_s_setup_cmplt,
         i_i2c_scl_s_hld_cmplt, i_i2c_scl_lcnt_cmplt, i_i2c_scl_p_setup_en,
         i_i2c_scl_s_setup_en, i_i2c_scl_hcnt_en, i_i2c_slv_tx_cmplt,
         i_i2c_slv_tx_ready_unconn, i_i2c_scl_hld_low_en, i_i2c_byte_wait_scl,
         i_i2c_slv_fifo_filled_and_flushed_sync, i_i2c_slv_rx_aborted_sync,
         i_i2c_activity, i_i2c_slv_activity_sync, i_i2c_mst_activity_sync,
         i_i2c_slv_clr_leftover_flg_edg, i_i2c_tx_abrt_flg_edg,
         i_i2c_ic_clr_gen_call_en, i_i2c_ic_clr_start_det_en,
         i_i2c_ic_clr_stop_det_en, i_i2c_ic_clr_activity_en,
         i_i2c_ic_clr_rx_done_en, i_i2c_ic_clr_tx_abrt_en,
         i_i2c_ic_clr_rd_req_en, i_i2c_ic_clr_tx_over_en,
         i_i2c_ic_clr_rx_over_en, i_i2c_ic_clr_rx_under_en,
         i_i2c_ic_clr_intr_en, i_i2c_tx_empty_ctrl,
         i_i2c_slv_fifo_filled_and_flushed, i_i2c_slv_rx_aborted,
         i_i2c_ic_ack_general_call_sync, i_i2c_ic_slave_en_sync,
         i_i2c_p_det_ifaddr_sync, i_i2c_ic_ss_sync, i_i2c_ic_fs_sync,
         i_i2c_ic_abort_sync, i_i2c_ic_ack_general_call, i_i2c_p_det_ifaddr,
         i_i2c_ic_slave_en, i_i2c_ic_rstrt_en, i_i2c_ic_10bit_slv, i_i2c_ic_ss,
         i_i2c_ic_fs, i_i2c_ic_hs, i_i2c_ic_10bit_mst, i_i2c_ic_master,
         i_i2c_set_tx_empty_en_flg, i_i2c_slv_clr_leftover_flg,
         i_i2c_rx_push_flg, i_i2c_tx_pop_flg, i_i2c_rx_gen_call_flg,
         i_i2c_s_det_flg, i_i2c_p_det_flg, i_i2c_ic_rd_req_flg,
         i_i2c_rx_done_flg, i_i2c_tx_abrt_flg, i_i2c_rx_addr_10bit,
         i_i2c_hs_mcode_en, i_i2c_ic_enable_sync, i_i2c_re_start_en,
         i_i2c_start_en, i_i2c_rx_current_src_en, i_i2c_tx_current_src_en,
         i_i2c_set_tx_empty_en, i_i2c_rx_push, i_i2c_tx_pop, i_i2c_rx_gen_call,
         i_i2c_s_det, i_i2c_p_det_intr, i_i2c_slv_activity, i_i2c_mst_activity,
         i_ssi_mst_contention, i_ssi_load_start_bit, i_ssi_rx_push,
         i_ssi_tx_pop, i_ssi_sclk_fe, i_ssi_sclk_re, i_ssi_start_xfer,
         i_ssi_baud2, i_ssi_ser_0_, i_ssi_sclk_active, i_ssi_fsm_multi_mst,
         i_ssi_ssi_en_int, i_ssi_rx_full, i_ssi_tx_full, i_ssi_tx_pop_sync,
         i_ssi_fsm_busy, i_ssi_fsm_sleep, i_ahb_U_dfltslv_N4,
         i_ahb_U_dfltslv_next_state, i_ahb_U_dfltslv_current_state,
         i_apb_U_DW_apb_ahbsif_N727, i_apb_U_DW_apb_ahbsif_use_saved_c,
         i_apb_U_DW_apb_ahbsif_piped_hwrite_c,
         i_apb_U_DW_apb_ahbsif_pipeline_c,
         i_apb_U_DW_apb_ahbsif_use_saved_data, i_i2c_U_DW_apb_i2c_toggle_N33,
         i_i2c_U_DW_apb_i2c_toggle_N32, i_i2c_U_DW_apb_i2c_toggle_N31,
         i_i2c_U_DW_apb_i2c_toggle_N30, i_i2c_U_DW_apb_i2c_toggle_N29,
         i_i2c_U_DW_apb_i2c_toggle_rx_gen_call_r,
         i_i2c_U_DW_apb_i2c_toggle_tx_abrt_r,
         i_i2c_U_DW_apb_i2c_toggle_tx_abrt,
         i_i2c_U_DW_apb_i2c_sync_tx_empty_sync_r,
         i_i2c_U_DW_apb_i2c_sync_ic_rstrt_en_sync_inv,
         i_i2c_U_DW_apb_i2c_sync_ic_10bit_slv_sync_inv,
         i_i2c_U_DW_apb_i2c_sync_tx_empty_int_inv,
         i_i2c_U_DW_apb_i2c_sync_ic_10bit_mst_sync_inv,
         i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv,
         i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv,
         i_i2c_U_DW_apb_i2c_intctl_N4,
         i_i2c_U_DW_apb_i2c_intctl_set_tx_empty_en_flg_sync_q,
         i_i2c_U_DW_apb_i2c_intctl_slv_clr_leftover_flg_sync_q,
         i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync_q,
         i_i2c_U_DW_apb_i2c_intctl_s_det_flg_sync_q,
         i_i2c_U_DW_apb_i2c_intctl_p_det_flg_sync_q,
         i_i2c_U_DW_apb_i2c_intctl_ic_rd_req_flg_sync_q,
         i_i2c_U_DW_apb_i2c_intctl_rx_done_flg_sync_q,
         i_i2c_U_DW_apb_i2c_intctl_tx_abrt_flg_sync_q,
         i_i2c_U_DW_apb_i2c_intctl_set_tx_empty_en_flg_sync,
         i_i2c_U_DW_apb_i2c_intctl_slv_clr_leftover_flg_sync,
         i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync,
         i_i2c_U_DW_apb_i2c_intctl_s_det_flg_sync,
         i_i2c_U_DW_apb_i2c_intctl_p_det_flg_sync,
         i_i2c_U_DW_apb_i2c_intctl_ic_rd_req_flg_sync,
         i_i2c_U_DW_apb_i2c_intctl_rx_done_flg_sync,
         i_i2c_U_DW_apb_i2c_intctl_tx_abrt_flg_sync,
         i_i2c_U_DW_apb_i2c_tx_shift_N403, i_i2c_U_DW_apb_i2c_tx_shift_N402,
         i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly2,
         i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly1,
         i_i2c_U_DW_apb_i2c_tx_shift_N281,
         i_i2c_U_DW_apb_i2c_tx_shift_stop_sda_gate_r,
         i_i2c_U_DW_apb_i2c_tx_shift_N272,
         i_i2c_U_DW_apb_i2c_tx_shift_start_sda_gate_r,
         i_i2c_U_DW_apb_i2c_tx_shift_slv_data_sda,
         i_i2c_U_DW_apb_i2c_tx_shift_data_sda,
         i_i2c_U_DW_apb_i2c_tx_shift_data_sda_prev_r,
         i_i2c_U_DW_apb_i2c_tx_shift_stop_sda,
         i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda,
         i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda_r,
         i_i2c_U_DW_apb_i2c_tx_shift_start_sda,
         i_i2c_U_DW_apb_i2c_tx_shift_byte_wait_en,
         i_i2c_U_DW_apb_i2c_tx_shift_mst_tx_bwen,
         i_i2c_U_DW_apb_i2c_tx_shift_N90,
         i_i2c_U_DW_apb_i2c_tx_shift_data_scl_lcnt_en,
         i_i2c_U_DW_apb_i2c_tx_shift_re_scl_s_hld_en,
         i_i2c_U_DW_apb_i2c_tx_shift_st_scl_s_hld_en,
         i_i2c_U_DW_apb_i2c_tx_shift_N85,
         i_i2c_U_DW_apb_i2c_tx_shift_mst_slv_ack_ext_r,
         i_i2c_U_DW_apb_i2c_tx_shift_mst_slv_ack_ext,
         i_i2c_U_DW_apb_i2c_tx_shift_N74,
         i_i2c_U_DW_apb_i2c_tx_shift_ic_data_oe_early,
         i_i2c_U_DW_apb_i2c_tx_shift_scl_hld_low_en_r,
         i_i2c_U_DW_apb_i2c_tx_shift_stop_scl_lcnt_en,
         i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl_lcnt_en,
         i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl,
         i_i2c_U_DW_apb_i2c_tx_shift_stop_scl,
         i_i2c_U_DW_apb_i2c_tx_shift_data_scl,
         i_i2c_U_DW_apb_i2c_rx_shift_rx_slv_read_s,
         i_i2c_U_DW_apb_i2c_rx_shift_N30,
         i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_3_,
         i_i2c_U_DW_apb_i2c_slvfsm_N284,
         i_i2c_U_DW_apb_i2c_slvfsm_ic_enable_sync_vld,
         i_i2c_U_DW_apb_i2c_slvfsm_slv_tx_flush, i_i2c_U_DW_apb_i2c_slvfsm_N39,
         i_i2c_U_DW_apb_i2c_slvfsm_N38, i_i2c_U_DW_apb_i2c_slvfsm_N37,
         i_i2c_U_DW_apb_i2c_slvfsm_N36, i_i2c_U_DW_apb_i2c_mstfsm_N487,
         i_i2c_U_DW_apb_i2c_mstfsm_mst_gen_ack_en_r,
         i_i2c_U_DW_apb_i2c_mstfsm_N421, i_i2c_U_DW_apb_i2c_mstfsm_N382,
         i_i2c_U_DW_apb_i2c_mstfsm_N252,
         i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_sync_d,
         i_i2c_U_DW_apb_i2c_mstfsm_delay_stop_en,
         i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_chk_win,
         i_i2c_U_DW_apb_i2c_mstfsm_tx_empty_hld,
         i_i2c_U_DW_apb_i2c_mstfsm_abrt_in_idle,
         i_i2c_U_DW_apb_i2c_mstfsm_mst_tx_flush,
         i_i2c_U_DW_apb_i2c_mstfsm_byte_waiting_q,
         i_i2c_U_DW_apb_i2c_mstfsm_old_is_read, i_i2c_U_DW_apb_i2c_mstfsm_N76,
         i_i2c_U_DW_apb_i2c_mstfsm_N75, i_i2c_U_DW_apb_i2c_mstfsm_N74,
         i_i2c_U_DW_apb_i2c_mstfsm_N73, i_i2c_U_DW_apb_i2c_mstfsm_N72,
         i_i2c_U_DW_apb_i2c_mstfsm_addr_1byte_sent,
         i_i2c_U_DW_apb_i2c_mstfsm_addr_2byte_sent,
         i_i2c_U_DW_apb_i2c_rx_filter_N241,
         i_i2c_U_DW_apb_i2c_rx_filter_slv_arb_lost,
         i_i2c_U_DW_apb_i2c_rx_filter_mst_arb_lost,
         i_i2c_U_DW_apb_i2c_rx_filter_N207,
         i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_q,
         i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_qq,
         i_i2c_U_DW_apb_i2c_rx_filter_sda_post_hold_done,
         i_i2c_U_DW_apb_i2c_rx_filter_N130, i_i2c_U_DW_apb_i2c_rx_filter_N129,
         i_i2c_U_DW_apb_i2c_rx_filter_N128, i_i2c_U_DW_apb_i2c_rx_filter_N127,
         i_i2c_U_DW_apb_i2c_rx_filter_N126, i_i2c_U_DW_apb_i2c_rx_filter_N125,
         i_i2c_U_DW_apb_i2c_rx_filter_N124, i_i2c_U_DW_apb_i2c_rx_filter_N123,
         i_i2c_U_DW_apb_i2c_rx_filter_sda_data_int,
         i_i2c_U_DW_apb_i2c_rx_filter_N89, i_i2c_U_DW_apb_i2c_rx_filter_N88,
         i_i2c_U_DW_apb_i2c_rx_filter_N87, i_i2c_U_DW_apb_i2c_rx_filter_N86,
         i_i2c_U_DW_apb_i2c_rx_filter_N85, i_i2c_U_DW_apb_i2c_rx_filter_N84,
         i_i2c_U_DW_apb_i2c_rx_filter_N83, i_i2c_U_DW_apb_i2c_rx_filter_N82,
         i_i2c_U_DW_apb_i2c_rx_filter_scl_clk_int,
         i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r,
         i_i2c_U_DW_apb_i2c_rx_filter_ic_hs, i_i2c_U_DW_apb_i2c_rx_filter_N50,
         i_i2c_U_DW_apb_i2c_rx_filter_hs_mcode_fed_dtctd_r,
         i_i2c_U_DW_apb_i2c_rx_filter_hs_mcode_en_r,
         i_i2c_U_DW_apb_i2c_rx_filter_rx_hs_mcode_r,
         i_i2c_U_DW_apb_i2c_rx_filter_scl_edg_hl_q,
         i_i2c_U_DW_apb_i2c_rx_filter_s_det_int,
         i_i2c_U_DW_apb_i2c_rx_filter_sda_int_q,
         i_i2c_U_DW_apb_i2c_rx_filter_scl_int_q,
         i_i2c_U_DW_apb_i2c_clk_gen_scl_int_d,
         i_i2c_U_DW_apb_i2c_clk_gen_scl_hcnt_cmplt_int,
         i_i2c_U_DW_apb_i2c_clk_gen_N77, i_i2c_U_DW_apb_i2c_clk_gen_N76,
         i_i2c_U_DW_apb_i2c_clk_gen_N75, i_i2c_U_DW_apb_i2c_clk_gen_N74,
         i_i2c_U_DW_apb_i2c_clk_gen_N73, i_i2c_U_DW_apb_i2c_clk_gen_N72,
         i_i2c_U_DW_apb_i2c_clk_gen_N71, i_i2c_U_DW_apb_i2c_clk_gen_N70,
         i_i2c_U_DW_apb_i2c_clk_gen_N69, i_i2c_U_DW_apb_i2c_clk_gen_N68,
         i_i2c_U_DW_apb_i2c_clk_gen_N67, i_i2c_U_DW_apb_i2c_clk_gen_N66,
         i_i2c_U_DW_apb_i2c_clk_gen_N65, i_i2c_U_DW_apb_i2c_clk_gen_N64,
         i_i2c_U_DW_apb_i2c_clk_gen_N63, i_i2c_U_DW_apb_i2c_clk_gen_N62,
         i_i2c_U_DW_apb_i2c_clk_gen_N51, i_i2c_U_DW_apb_i2c_clk_gen_count_en,
         i_i2c_U_DW_apb_i2c_fifo_i_rx_almost_full,
         i_i2c_U_DW_apb_i2c_fifo_rx_error_ir,
         i_i2c_U_DW_apb_i2c_fifo_tx_error_ir,
         i_i2c_U_DW_apb_i2c_fifo_rx_push_sync_dly,
         i_i2c_U_DW_apb_i2c_fifo_rx_pop_dly,
         i_i2c_U_DW_apb_i2c_fifo_tx_pop_sync_dly,
         i_i2c_U_DW_apb_i2c_fifo_tx_push_dly,
         i_i2c_U_DW_apb_i2c_fifo_rx_push_flg_sync_q,
         i_i2c_U_DW_apb_i2c_fifo_tx_pop_flg_sync_q,
         i_i2c_U_DW_apb_i2c_fifo_rx_push_flg_sync,
         i_i2c_U_DW_apb_i2c_fifo_tx_pop_flg_sync, i_ssi_U_regfile_N452,
         i_ssi_U_regfile_N451, i_ssi_U_regfile_multi_mst_edge,
         i_ssi_U_regfile_sr_6_, i_ssi_U_regfile_ctrlr0_ir_int_7,
         i_ssi_U_sclkgen_N75, i_ssi_U_sclkgen_N74, i_ssi_U_sclkgen_N55,
         i_ssi_U_sclkgen_N54, i_ssi_U_sclkgen_N53, i_ssi_U_sclkgen_N52,
         i_ssi_U_sclkgen_N51, i_ssi_U_sclkgen_N50, i_ssi_U_sclkgen_N49,
         i_ssi_U_sclkgen_N48, i_ssi_U_sclkgen_N47, i_ssi_U_sclkgen_N46,
         i_ssi_U_sclkgen_N45, i_ssi_U_sclkgen_N44, i_ssi_U_sclkgen_N43,
         i_ssi_U_sclkgen_N42, i_ssi_U_sclkgen_N41,
         i_ssi_U_fifo_switch_almost_full, i_ssi_U_fifo_rx_push_edge,
         i_ssi_U_fifo_tx_pop_edge, i_ssi_U_fifo_rx_error_ir,
         i_ssi_U_fifo_tx_error_ir, i_ssi_U_fifo_rx_push_sync_dly,
         i_ssi_U_fifo_rx_pop_dly, i_ssi_U_fifo_tx_pop_sync_dly,
         i_ssi_U_fifo_tx_push_dly, i_ssi_U_mstfsm_abort_ir,
         i_ssi_U_mstfsm_N223, i_ssi_U_mstfsm_N222, i_ssi_U_mstfsm_N221,
         i_ssi_U_mstfsm_N220, i_ssi_U_mstfsm_last_frame,
         i_ssi_U_mstfsm_spi1_control, i_ssi_U_mstfsm_spi0_control,
         i_ssi_U_mstfsm_c_done_ir, i_ssi_U_mstfsm_ss_in_n_sync,
         i_ssi_U_mstfsm_tx_load_en_int, i_ssi_U_intctl_N33, i_ssi_U_intctl_N2,
         i_i2c_U_DW_apb_i2c_sync_U_ic_enable_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_abort_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_gen_call_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_master_1_sync_N2,
         i_i2c_U_DW_apb_i2c_sync_U_ic_master_1_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_hs_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_fs_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_ss_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_mst_1_sync_N2,
         i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_mst_1_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_tx_empty_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_slv_1_sync_N2,
         i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_slv_1_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_rstrt_en_1_sync_N2,
         i_i2c_U_DW_apb_i2c_sync_U_ic_rstrt_en_1_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_slave_en_1_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_p_det_ifaddr_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_rx_done_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_ic_rd_req_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_p_det_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_s_det_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_rx_gen_call_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_slv_clr_leftover_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_set_tx_empty_en_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_mst_activity_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_slv_activity_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_slv_rx_aborted_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_slv_fifo_filled_and_flushed_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_data_d_int_0_,
         i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_data_d_int_0_,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_pop_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_push_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N49,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N48,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N47,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N46,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N45,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N44,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N43,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N42,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N41,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N40,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N39,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N38,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N37,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N34,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N33,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_almost_empty_n,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_rd_addr_at_max,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_wr_addr_at_max,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_empty_n,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N49,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N48,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N47,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N46,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N45,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N44,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N43,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N42,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N41,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N40,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N39,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N38,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N37,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N36,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N33,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_rd_addr_at_max,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_wr_addr_at_max,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_empty_n, i_ssi_U_fifo_U_tx_fifo_N48,
         i_ssi_U_fifo_U_tx_fifo_N47, i_ssi_U_fifo_U_tx_fifo_N46,
         i_ssi_U_fifo_U_tx_fifo_N45, i_ssi_U_fifo_U_tx_fifo_N43,
         i_ssi_U_fifo_U_tx_fifo_N42, i_ssi_U_fifo_U_tx_fifo_N41,
         i_ssi_U_fifo_U_tx_fifo_N40, i_ssi_U_fifo_U_tx_fifo_N39,
         i_ssi_U_fifo_U_tx_fifo_N38, i_ssi_U_fifo_U_tx_fifo_N37,
         i_ssi_U_fifo_U_tx_fifo_N34, i_ssi_U_fifo_U_tx_fifo_N33,
         i_ssi_U_fifo_U_tx_fifo_almost_empty_n,
         i_ssi_U_fifo_U_tx_fifo_rd_addr_at_max,
         i_ssi_U_fifo_U_tx_fifo_wr_addr_at_max, i_ssi_U_fifo_U_tx_fifo_empty_n,
         i_ssi_U_fifo_U_rx_fifo_N49, i_ssi_U_fifo_U_rx_fifo_N48,
         i_ssi_U_fifo_U_rx_fifo_N47, i_ssi_U_fifo_U_rx_fifo_N46,
         i_ssi_U_fifo_U_rx_fifo_N45, i_ssi_U_fifo_U_rx_fifo_N43,
         i_ssi_U_fifo_U_rx_fifo_N42, i_ssi_U_fifo_U_rx_fifo_N41,
         i_ssi_U_fifo_U_rx_fifo_N40, i_ssi_U_fifo_U_rx_fifo_N39,
         i_ssi_U_fifo_U_rx_fifo_N38, i_ssi_U_fifo_U_rx_fifo_N36,
         i_ssi_U_fifo_U_rx_fifo_N33, i_ssi_U_fifo_U_rx_fifo_rd_addr_at_max,
         i_ssi_U_fifo_U_rx_fifo_wr_addr_at_max, i_ssi_U_fifo_U_rx_fifo_empty_n,
         i_ssi_U_shift_U_tx_shifter_load_start_bit_ir,
         i_ssi_U_mstfsm_U_ss_in_n_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_U_SYNC_N2,
         i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_U_SYNC_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_U_SYNC_N2,
         i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_U_SYNC_next_sample_syncm1_0_,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4824, n4825, n4826, n4841, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5241, n5242, n5245, n5246, n5247, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11726, n11747, n11748, n11759, n11760, n11761, n11762,
         n11763, n11764, ex_i_ahb_AHB_Slave_PID_hready, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14;
  wire   [31:12] i_apb_paddr;
  wire   [31:0] i_ssi_prdata;
  wire   [30:0] i_i2c_prdata;
  wire   [23:0] i_apb_pwdata_int;
  wire   [2:0] i_i2c_rx_rd_addr;
  wire   [2:0] i_i2c_rx_wr_addr;
  wire   [2:0] i_i2c_tx_rd_addr;
  wire   [2:0] i_i2c_tx_wr_addr;
  wire   [7:0] i_i2c_rx_pop_data;
  wire   [2:0] i_i2c_ic_tx_tl;
  wire   [2:0] i_i2c_ic_rx_tl;
  wire   [15:0] i_i2c_ic_fs_hcnt;
  wire   [15:0] i_i2c_ic_fs_lcnt;
  wire   [15:0] i_i2c_ic_lcnt;
  wire   [15:0] i_i2c_ic_hcnt;
  wire   [7:0] i_i2c_ic_fs_spklen;
  wire   [7:0] i_i2c_ic_hs_spklen;
  wire   [10:0] i_i2c_ic_tar;
  wire   [2:0] i_i2c_ic_hs_maddr;
  wire   [7:0] i_i2c_ic_sda_setup;
  wire   [30:0] i_i2c_iprdata;
  wire   [7:0] i_i2c_rx_push_data;
  wire   [9:0] i_i2c_ic_sar;
  wire   [3:0] i_i2c_mst_rx_bit_count;
  wire   [8:0] i_i2c_tx_fifo_data_buf;
  wire   [16:0] i_i2c_ic_tx_abrt_source;
  wire   [11:0] i_i2c_ic_raw_intr_stat;
  wire   [11:0] i_i2c_ic_intr_stat;
  wire   [11:0] i_i2c_ic_intr_mask;
  wire   [7:0] i_i2c_ic_sda_rx_hold_sync;
  wire   [15:0] i_i2c_ic_sda_tx_hold_sync;
  wire   [23:0] i_i2c_ic_sda_hold;
  wire   [1:0] i_i2c_ic_enable;
  wire   [16:0] i_i2c_tx_abrt_source;
  wire   [3:0] i_i2c_slv_debug_cstate;
  wire   [4:0] i_i2c_mst_debug_cstate;
  wire   [15:0] i_ssi_rx_push_data;
  wire   [2:0] i_ssi_rx_rd_addr;
  wire   [2:0] i_ssi_rx_wr_addr;
  wire   [2:0] i_ssi_tx_rd_addr;
  wire   [2:0] i_ssi_tx_wr_addr;
  wire   [2:0] i_ssi_rxftlr;
  wire   [2:0] i_ssi_txftlr;
  wire   [15:1] i_ssi_baudr;
  wire   [2:0] i_ssi_mwcr;
  wire   [5:0] i_ssi_imr;
  wire   [5:0] i_ssi_risr;
  wire   [5:0] i_ssi_reg_addr;
  wire   [3:0] i_ssi_cfs;
  wire   [1:0] i_ssi_tmod;
  wire   [11:10] i_ssi_ctrlr0;
  wire   [3:0] i_ssi_dfs;
  wire   [4:1] i_ahb_U_mux_hsel_prev;
  wire   [23:0] i_apb_U_DW_apb_ahbsif_saved_hwdata32_c;
  wire   [31:2] i_apb_U_DW_apb_ahbsif_saved_haddr_c;
  wire   [17:2] i_apb_U_DW_apb_ahbsif_piped_haddr_c;
  wire   [2:0] i_apb_U_DW_apb_ahbsif_nextstate;
  wire   [2:0] i_apb_U_DW_apb_ahbsif_state;
  wire   [16:0] i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q;
  wire   [16:0] i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync;
  wire   [15:0] i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r;
  wire   [7:0] i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf;
  wire   [3:0] i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count;
  wire   [3:0] i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count;
  wire   [3:0] i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr;
  wire   [7:0] i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg;
  wire   [7:0] i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg;
  wire   [2:0] i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0;
  wire   [7:0] i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count;
  wire  
         [3:0] i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en
;
  wire   [1:0] i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt;
  wire   [7:0] i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt;
  wire   [7:0] i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt;
  wire   [7:0] i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt;
  wire   [15:0] i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr;
  wire   [15:0] i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr;
  wire   [15:0] i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr;
  wire   [15:0] i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr;
  wire   [15:0] i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr;
  wire   [15:0] i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr;
  wire   [15:0] i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr;
  wire   [2:0] i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn;
  wire   [2:0] i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn;
  wire   [7:0] i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr;
  wire   [63:0] i_i2c_U_dff_rx_mem;
  wire   [71:0] i_i2c_U_dff_tx_mem;
  wire   [3:0] i_ssi_U_regfile_rxflr;
  wire   [3:0] i_ssi_U_regfile_txflr;
  wire   [15:0] i_ssi_U_regfile_ctrlr1_int;
  wire   [5:4] i_ssi_U_regfile_ctrlr0_ir_int;
  wire   [15:0] i_ssi_U_sclkgen_ssi_cnt;
  wire   [2:0] i_ssi_U_fifo_unconnected_rx_wrd_count;
  wire   [2:0] i_ssi_U_fifo_unconnected_tx_wrd_count;
  wire   [16:0] i_ssi_U_mstfsm_frame_cnt;
  wire   [3:0] i_ssi_U_mstfsm_c_state;
  wire   [3:0] i_ssi_U_mstfsm_ctrl_cnt;
  wire   [4:0] i_ssi_U_mstfsm_bit_cnt;
  wire   [127:0] i_ssi_U_dff_rx_mem;
  wire   [127:0] i_ssi_U_dff_tx_mem;
  wire   [23:0] i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1;
  wire  
         [16:0] i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1
;
  wire   [15:0] i_ssi_U_shift_U_tx_shifter_tx_buffer;
  wire   [15:0] i_ssi_U_shift_U_tx_shifter_tx_shift_reg;
  wire   [15:0] i_ssi_U_shift_U_rx_shifter_rx_shift_reg;
  assign ex_i_ahb_AHB_Slave_RAM_haddr[31] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[31];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[31] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[31];
  assign ex_i_ahb_AHB_Slave_PID_haddr[31] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[31];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[30] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[30];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[30] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[30];
  assign ex_i_ahb_AHB_Slave_PID_haddr[30] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[30];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[29] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[29];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[29] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[29];
  assign ex_i_ahb_AHB_Slave_PID_haddr[29] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[29];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[28] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[28];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[28] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[28];
  assign ex_i_ahb_AHB_Slave_PID_haddr[28] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[28];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[27] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[27];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[27] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[27];
  assign ex_i_ahb_AHB_Slave_PID_haddr[27] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[27];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[26] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[26];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[26] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[26];
  assign ex_i_ahb_AHB_Slave_PID_haddr[26] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[26];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[25] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[25];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[25] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[25];
  assign ex_i_ahb_AHB_Slave_PID_haddr[25] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[25];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[24] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[24];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[24] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[24];
  assign ex_i_ahb_AHB_Slave_PID_haddr[24] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[24];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[23] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[23];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[23] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[23];
  assign ex_i_ahb_AHB_Slave_PID_haddr[23] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[23];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[22] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[22];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[22] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[22];
  assign ex_i_ahb_AHB_Slave_PID_haddr[22] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[22];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[21] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[21];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[21] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[21];
  assign ex_i_ahb_AHB_Slave_PID_haddr[21] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[21];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[20] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[20];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[20] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[20];
  assign ex_i_ahb_AHB_Slave_PID_haddr[20] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[20];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[19] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[19];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[19] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[19];
  assign ex_i_ahb_AHB_Slave_PID_haddr[19] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[19];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[18] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[18];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[18] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[18];
  assign ex_i_ahb_AHB_Slave_PID_haddr[18] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[18];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[17] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[17];
  assign ex_i_ahb_AHB_Slave_PID_haddr[17] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[17];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[17] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[17];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[16] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[16];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[16] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[16];
  assign ex_i_ahb_AHB_Slave_PID_haddr[16] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[16];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[15] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[15];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[15] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[15];
  assign ex_i_ahb_AHB_Slave_PID_haddr[15] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[15];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[14] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[14];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[14] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[14];
  assign ex_i_ahb_AHB_Slave_PID_haddr[14] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[14];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[13] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[13];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[13] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[13];
  assign ex_i_ahb_AHB_Slave_PID_haddr[13] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[13];
  assign ex_i_ahb_AHB_Slave_PID_haddr[12] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[12];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[12] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[12];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[12] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[12];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[11] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[11];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[11] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[11];
  assign ex_i_ahb_AHB_Slave_PID_haddr[11] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[11];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[10] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[10];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[10] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[10];
  assign ex_i_ahb_AHB_Slave_PID_haddr[10] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[10];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[9] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[9];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[9] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[9];
  assign ex_i_ahb_AHB_Slave_PID_haddr[9] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[9];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[8] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[8];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[8] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[8];
  assign ex_i_ahb_AHB_Slave_PID_haddr[8] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[8];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[7] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[7];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[7] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[7];
  assign ex_i_ahb_AHB_Slave_PID_haddr[7] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[7];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[6] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[6];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[6] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[6];
  assign ex_i_ahb_AHB_Slave_PID_haddr[6] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[6];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[5] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[5];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[5] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[5];
  assign ex_i_ahb_AHB_Slave_PID_haddr[5] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[5];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[4] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[4];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[4] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[4];
  assign ex_i_ahb_AHB_Slave_PID_haddr[4] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[4];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[3] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[3];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[3] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[3];
  assign ex_i_ahb_AHB_Slave_PID_haddr[3] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[3];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[2];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[2];
  assign ex_i_ahb_AHB_Slave_PID_haddr[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[2];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[1];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[1];
  assign ex_i_ahb_AHB_Slave_PID_haddr[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[1];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[0];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[0];
  assign ex_i_ahb_AHB_Slave_PID_haddr[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[0];
  assign ex_i_ahb_AHB_Slave_RAM_hburst[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hburst[2];
  assign ex_i_ahb_AHB_Slave_PWM_hburst[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hburst[2];
  assign ex_i_ahb_AHB_Slave_PID_hburst[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hburst[2];
  assign ex_i_ahb_AHB_Slave_RAM_hburst[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hburst[1];
  assign ex_i_ahb_AHB_Slave_PWM_hburst[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hburst[1];
  assign ex_i_ahb_AHB_Slave_PID_hburst[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hburst[1];
  assign ex_i_ahb_AHB_Slave_RAM_hburst[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hburst[0];
  assign ex_i_ahb_AHB_Slave_PWM_hburst[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hburst[0];
  assign ex_i_ahb_AHB_Slave_PID_hburst[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hburst[0];
  assign ex_i_ahb_AHB_Slave_RAM_hprot[3] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[3];
  assign ex_i_ahb_AHB_Slave_PWM_hprot[3] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[3];
  assign ex_i_ahb_AHB_Slave_PID_hprot[3] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[3];
  assign ex_i_ahb_AHB_Slave_RAM_hprot[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[2];
  assign ex_i_ahb_AHB_Slave_PWM_hprot[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[2];
  assign ex_i_ahb_AHB_Slave_PID_hprot[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[2];
  assign ex_i_ahb_AHB_Slave_RAM_hprot[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[1];
  assign ex_i_ahb_AHB_Slave_PWM_hprot[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[1];
  assign ex_i_ahb_AHB_Slave_PID_hprot[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[1];
  assign ex_i_ahb_AHB_Slave_RAM_hprot[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[0];
  assign ex_i_ahb_AHB_Slave_PWM_hprot[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[0];
  assign ex_i_ahb_AHB_Slave_PID_hprot[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[0];
  assign ex_i_ahb_AHB_Slave_RAM_hsize[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hsize[2];
  assign ex_i_ahb_AHB_Slave_PWM_hsize[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hsize[2];
  assign ex_i_ahb_AHB_Slave_PID_hsize[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hsize[2];
  assign ex_i_ahb_AHB_Slave_RAM_hsize[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hsize[1];
  assign ex_i_ahb_AHB_Slave_PWM_hsize[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hsize[1];
  assign ex_i_ahb_AHB_Slave_PID_hsize[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hsize[1];
  assign ex_i_ahb_AHB_Slave_RAM_hsize[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hsize[0];
  assign ex_i_ahb_AHB_Slave_PWM_hsize[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hsize[0];
  assign ex_i_ahb_AHB_Slave_PID_hsize[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hsize[0];
  assign ex_i_ahb_AHB_Slave_RAM_htrans[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_htrans[1];
  assign ex_i_ahb_AHB_Slave_PWM_htrans[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_htrans[1];
  assign ex_i_ahb_AHB_Slave_PID_htrans[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_htrans[1];
  assign ex_i_ahb_AHB_Slave_RAM_htrans[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_htrans[0];
  assign ex_i_ahb_AHB_Slave_PWM_htrans[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_htrans[0];
  assign ex_i_ahb_AHB_Slave_PID_htrans[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_htrans[0];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[31] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[31];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[31] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[31];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[31] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[31];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[30] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[30];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[30] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[30];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[30] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[30];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[29] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[29];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[29] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[29];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[29] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[29];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[28] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[28];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[28] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[28];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[28] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[28];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[27] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[27];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[27] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[27];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[27] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[27];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[26] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[26];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[26] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[26];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[26] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[26];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[25] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[25];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[25] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[25];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[25] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[25];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[24] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[24];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[24] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[24];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[24] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[24];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[23] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[23];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[23] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[23];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[23] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[23];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[22] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[22];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[22] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[22];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[22] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[22];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[21] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[21];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[21] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[21];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[21] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[21];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[20] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[20];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[20] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[20];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[20] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[20];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[19] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[19];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[19] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[19];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[19] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[19];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[18] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[18];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[18] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[18];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[18] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[18];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[17] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[17];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[17] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[17];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[17] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[17];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[16] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[16];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[16] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[16];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[16] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[16];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[15] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[15];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[15] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[15];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[15] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[15];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[14] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[14];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[14] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[14];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[14] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[14];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[13] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[13];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[13] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[13];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[13] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[13];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[12] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[12];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[12] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[12];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[12] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[12];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[11] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[11];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[11] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[11];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[11] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[11];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[10] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[10];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[10] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[10];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[10] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[10];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[9] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[9];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[9] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[9];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[9] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[9];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[8] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[8];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[8] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[8];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[8] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[8];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[7] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[7];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[7] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[7];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[7] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[7];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[6] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[6];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[6] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[6];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[6] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[6];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[5] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[5];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[5] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[5];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[5] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[5];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[4] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[4];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[4] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[4];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[4] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[4];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[3] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[3];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[3] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[3];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[3] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[3];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[2];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[2];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[2];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[1];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[1];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[1];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[0];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[0];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[0];
  assign ex_i_ahb_AHB_Slave_PID_hwrite = ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite;
  assign ex_i_ahb_AHB_Slave_RAM_hwrite = ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite;
  assign ex_i_ahb_AHB_Slave_PWM_hwrite = ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite;
  assign ex_i_ahb_AHB_Slave_RAM_hmastlock = ex_i_ahb_AHB_Slave_PID_hmastlock;
  assign ex_i_ahb_AHB_Slave_PWM_hmastlock = ex_i_ahb_AHB_Slave_PID_hmastlock;
  assign i_ahb_hmaster_data[0] = 1'b1;
  assign i_ahb_hmaster_data[3] = 1'b0;
  assign i_ahb_hmaster_data[2] = 1'b0;
  assign i_ahb_hmaster_data[1] = 1'b0;
  assign ex_i_ahb_AHB_Slave_RAM_hready = ex_i_ahb_AHB_Slave_PID_hready;
  assign ex_i_ahb_AHB_MASTER_CORTEXM0_hready = ex_i_ahb_AHB_Slave_PID_hready;
  assign ex_i_ahb_AHB_Slave_PWM_hready = ex_i_ahb_AHB_Slave_PID_hready;

  i_i2c_DW_apb_i2c_regfile i_i2c_U_DW_apb_i2c_regfile ( .pclk(PCLK_pclk), 
        .presetn(PRESETn_presetn), .wr_en(i_i2c_wr_en), .rd_en(n11762), 
        .byte_en({1'b1, 1'b1, 1'b1, 1'b1}), .reg_addr(i_ssi_reg_addr), 
        .ipwdata({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        i_apb_pwdata_int}), .iprdata({SYNOPSYS_UNCONNECTED_1, 
        i_i2c_iprdata[30:29], SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        i_i2c_iprdata[26:0]}), .ic_clr_intr_en(i_i2c_ic_clr_intr_en), 
        .ic_clr_rx_under_en(i_i2c_ic_clr_rx_under_en), .ic_clr_rx_over_en(
        i_i2c_ic_clr_rx_over_en), .ic_clr_tx_over_en(i_i2c_ic_clr_tx_over_en), 
        .ic_clr_rd_req_en(i_i2c_ic_clr_rd_req_en), .ic_clr_tx_abrt_en(
        i_i2c_ic_clr_tx_abrt_en), .ic_clr_rx_done_en(i_i2c_ic_clr_rx_done_en), 
        .ic_clr_activity_en(i_i2c_ic_clr_activity_en), .ic_clr_stop_det_en(
        i_i2c_ic_clr_stop_det_en), .ic_clr_start_det_en(
        i_i2c_ic_clr_start_det_en), .ic_clr_gen_call_en(
        i_i2c_ic_clr_gen_call_en), .mst_activity(i_i2c_mst_activity_sync), 
        .slv_activity(i_i2c_slv_activity_sync), .activity(i_i2c_activity), 
        .ic_tx_abrt_source(i_i2c_ic_tx_abrt_source), .ic_en(i_i2c_ic_en), 
        .slv_rx_aborted_sync(i_i2c_slv_rx_aborted_sync), 
        .slv_fifo_filled_and_flushed_sync(
        i_i2c_slv_fifo_filled_and_flushed_sync), .ic_tar({
        i_i2c_U_DW_apb_i2c_mstfsm_N252, i_i2c_ic_tar}), .ic_sar(i_i2c_ic_sar), 
        .ic_hs_maddr(i_i2c_ic_hs_maddr), .ic_fs_hcnt(i_i2c_ic_fs_hcnt), 
        .ic_fs_lcnt(i_i2c_ic_fs_lcnt), .ic_intr_mask({SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, i_i2c_ic_intr_mask}), .ic_rx_tl_int(
        i_i2c_ic_rx_tl), .ic_enable(i_i2c_ic_enable), .ic_hcnt(i_i2c_ic_hcnt), 
        .ic_lcnt(i_i2c_ic_lcnt), .ic_fs_spklen(i_i2c_ic_fs_spklen), 
        .ic_hs_spklen(i_i2c_ic_hs_spklen), .ic_intr_stat({1'b0, 1'b0, 
        i_i2c_ic_intr_stat}), .ic_raw_intr_stat({1'b0, 1'b0, 
        i_i2c_ic_raw_intr_stat}), .ic_hs(i_i2c_ic_hs), .ic_fs(i_i2c_ic_fs), 
        .ic_ss(i_i2c_ic_ss), .ic_master(i_i2c_ic_master), .ic_10bit_mst(
        i_i2c_ic_10bit_mst), .ic_10bit_slv(i_i2c_ic_10bit_slv), .ic_slave_en(
        i_i2c_ic_slave_en), .p_det_ifaddr(i_i2c_p_det_ifaddr), .tx_empty_ctrl(
        i_i2c_tx_empty_ctrl), .rx_pop_data(i_i2c_rx_pop_data), .tx_push_data({
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14}), .fifo_rst_n(
        i_i2c_fifo_rst_n), .tx_fifo_rst_n(i_i2c_tx_fifo_rst_n), .tx_pop_sync(
        i_i2c_tx_pop_sync), .rx_push_sync(i_i2c_rx_push_sync), .rx_pop(
        i_i2c_rx_pop), .tx_push(i_i2c_tx_push), .tx_empty(n5246), .rx_full(
        i_i2c_rx_full), .tx_full(i_i2c_tx_full), .rx_empty(n5247), 
        .tx_abrt_flg_edg(i_i2c_tx_abrt_flg_edg), .abrt_in_rcve_trns(
        i_i2c_abrt_in_rcve_trns), .slv_clr_leftover_flg_edg(
        i_i2c_slv_clr_leftover_flg_edg), .ic_rstrt_en(i_i2c_ic_rstrt_en), 
        .ic_sda_setup(i_i2c_ic_sda_setup), .ic_sda_hold(i_i2c_ic_sda_hold), 
        .ic_ack_general_call(i_i2c_ic_ack_general_call), .ic_tx_tl_2_(
        i_i2c_ic_tx_tl[2]), .ic_tx_tl_1_(i_i2c_ic_tx_tl[1]), .ic_tx_tl_0_(
        i_i2c_ic_tx_tl[0]) );
  drsp_1 i_ssi_U_mstfsm_tx_load_en_reg ( .ip(n4586), .ck(i_ssi_ssi_clk), .rb(
        1'b1), .s(n11764), .q(i_ssi_U_mstfsm_tx_load_en_int) );
  drsp_1 i_ssi_U_sclkgen_sclk_out_reg ( .ip(n4249), .ck(i_ssi_ssi_clk), .rb(
        1'b1), .s(n11764), .q(i_ssi_sclk_out) );
  drp_1 i_ahb_U_dfltslv_current_state_reg ( .ip(i_ahb_U_dfltslv_next_state), 
        .ck(HCLK_hclk), .rb(HRESETn_hresetn), .q(i_ahb_U_dfltslv_current_state) );
  drp_1 i_ahb_U_dfltslv_hresp_none_reg_0_ ( .ip(i_ahb_U_dfltslv_N4), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(i_ahb_hresp_none_0_) );
  drp_1 i_ahb_U_mux_hsel_prev_reg_4_ ( .ip(n4859), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ahb_U_mux_hsel_prev[4]) );
  drp_1 i_ahb_U_mux_hsel_prev_reg_3_ ( .ip(n4858), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ahb_U_mux_hsel_prev[3]) );
  drp_1 i_ahb_U_mux_hsel_prev_reg_2_ ( .ip(n4857), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ahb_U_mux_hsel_prev[2]) );
  drp_1 i_ahb_U_mux_hsel_prev_reg_1_ ( .ip(n4856), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ahb_U_mux_hsel_prev[1]) );
  drp_1 i_ahb_U_arblite_hmastlock_reg ( .ip(n4855), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(ex_i_ahb_AHB_Slave_PID_hmastlock) );
  drp_1 i_apb_U_DW_apb_ahbsif_pipeline_reg ( .ip(n4854), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_pipeline_c) );
  drp_1 i_apb_U_DW_apb_ahbsif_state_reg_1_ ( .ip(
        i_apb_U_DW_apb_ahbsif_nextstate[1]), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_state[1]) );
  drp_1 i_apb_U_DW_apb_ahbsif_state_reg_2_ ( .ip(
        i_apb_U_DW_apb_ahbsif_nextstate[2]), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_state[2]) );
  drp_1 i_apb_U_DW_apb_ahbsif_piped_hwrite_reg ( .ip(n4853), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_piped_hwrite_c) );
  drp_1 i_apb_U_DW_apb_ahbsif_piped_haddr_reg_2_ ( .ip(n4852), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_piped_haddr_c[2]) );
  drp_1 i_apb_U_DW_apb_ahbsif_piped_haddr_reg_3_ ( .ip(n4851), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_piped_haddr_c[3]) );
  drp_1 i_apb_U_DW_apb_ahbsif_piped_haddr_reg_4_ ( .ip(n4850), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_piped_haddr_c[4]) );
  drp_1 i_apb_U_DW_apb_ahbsif_piped_haddr_reg_5_ ( .ip(n4849), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_piped_haddr_c[5]) );
  drp_1 i_apb_U_DW_apb_ahbsif_piped_haddr_reg_6_ ( .ip(n4848), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_piped_haddr_c[6]) );
  drp_1 i_apb_U_DW_apb_ahbsif_piped_haddr_reg_7_ ( .ip(n4847), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_piped_haddr_c[7]) );
  drp_1 i_apb_U_DW_apb_ahbsif_piped_haddr_reg_12_ ( .ip(n4846), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_piped_haddr_c[12]) );
  drp_1 i_apb_U_DW_apb_ahbsif_piped_haddr_reg_17_ ( .ip(n4841), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_piped_haddr_c[17]) );
  drp_1 i_apb_U_DW_apb_ahbsif_use_saved_reg ( .ip(n4826), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_use_saved_c) );
  drp_1 i_apb_U_DW_apb_ahbsif_use_saved_data_reg ( .ip(
        i_apb_U_DW_apb_ahbsif_N727), .ck(HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_use_saved_data) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_0_ ( .ip(n4822), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[0]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_1_ ( .ip(n4821), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[1]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_2_ ( .ip(n4820), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[2]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_3_ ( .ip(n4819), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[3]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_4_ ( .ip(n4818), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[4]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_5_ ( .ip(n4817), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[5]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_6_ ( .ip(n4816), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[6]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_7_ ( .ip(n4815), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[7]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_8_ ( .ip(n4814), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[8]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_9_ ( .ip(n4813), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[9]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_10_ ( .ip(n4812), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[10]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_11_ ( .ip(n4811), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[11]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_12_ ( .ip(n4810), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[12]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_13_ ( .ip(n4809), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[13]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_14_ ( .ip(n4808), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[14]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_15_ ( .ip(n4807), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[15]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_16_ ( .ip(n4806), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[16]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_17_ ( .ip(n4805), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[17]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_18_ ( .ip(n4804), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[18]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_19_ ( .ip(n4803), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[19]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_20_ ( .ip(n4802), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[20]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_21_ ( .ip(n4801), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[21]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_22_ ( .ip(n4800), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[22]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_23_ ( .ip(n4799), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[23]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_2_ ( .ip(n4759), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[2]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_3_ ( .ip(n4758), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[3]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_4_ ( .ip(n4757), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[4]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_5_ ( .ip(n4756), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[5]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_6_ ( .ip(n4755), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[6]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_7_ ( .ip(n4754), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[7]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_12_ ( .ip(n4753), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[12]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_13_ ( .ip(n4752), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[13]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_14_ ( .ip(n4751), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[14]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_15_ ( .ip(n4750), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[15]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_16_ ( .ip(n4749), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[16]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_17_ ( .ip(n4748), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[17]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_18_ ( .ip(n4747), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[18]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_19_ ( .ip(n4746), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[19]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_20_ ( .ip(n4745), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[20]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_21_ ( .ip(n4744), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[21]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_22_ ( .ip(n4743), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[22]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_23_ ( .ip(n4742), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[23]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_24_ ( .ip(n4741), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[24]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_25_ ( .ip(n4740), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[25]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_26_ ( .ip(n4739), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[26]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_27_ ( .ip(n4738), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[27]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_28_ ( .ip(n4737), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[28]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_29_ ( .ip(n4736), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[29]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_30_ ( .ip(n4735), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[30]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_31_ ( .ip(n4734), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[31]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_0_ ( .ip(n4791), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[0]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_1_ ( .ip(n4790), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[1]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_2_ ( .ip(n4789), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[2]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_3_ ( .ip(n4788), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[3]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_4_ ( .ip(n4787), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[4]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_5_ ( .ip(n4786), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[5]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_6_ ( .ip(n4785), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[6]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_7_ ( .ip(n4784), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[7]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_8_ ( .ip(n4783), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[8]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_9_ ( .ip(n4782), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[9]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_10_ ( .ip(n4781), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[10]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_11_ ( .ip(n4780), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[11]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_12_ ( .ip(n4779), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[12]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_13_ ( .ip(n4778), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[13]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_14_ ( .ip(n4777), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[14]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_15_ ( .ip(n4776), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[15]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_16_ ( .ip(n4775), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[16]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_17_ ( .ip(n4774), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[17]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_18_ ( .ip(n4773), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[18]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_19_ ( .ip(n4772), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[19]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_20_ ( .ip(n4771), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[20]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_21_ ( .ip(n4770), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[21]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_22_ ( .ip(n4769), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[22]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_23_ ( .ip(n4768), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[23]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwrite_reg ( .ip(n4825), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_pwrite) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_2_ ( .ip(n4733), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ssi_reg_addr[0]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_3_ ( .ip(n4732), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ssi_reg_addr[1]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_4_ ( .ip(n4731), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ssi_reg_addr[2]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_5_ ( .ip(n4730), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ssi_reg_addr[3]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_6_ ( .ip(n4729), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ssi_reg_addr[4]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_7_ ( .ip(n4728), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ssi_reg_addr[5]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_12_ ( .ip(n4727), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[12]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_13_ ( .ip(n4726), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[13]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_14_ ( .ip(n4725), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[14]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_15_ ( .ip(n4724), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[15]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_16_ ( .ip(n4723), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[16]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_17_ ( .ip(n4722), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[17]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_18_ ( .ip(n4721), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[18]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_19_ ( .ip(n4720), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[19]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_20_ ( .ip(n4719), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[20]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_21_ ( .ip(n4718), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[21]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_22_ ( .ip(n4717), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[22]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_23_ ( .ip(n4716), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[23]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_24_ ( .ip(n4715), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[24]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_25_ ( .ip(n4714), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[25]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_26_ ( .ip(n4713), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[26]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_27_ ( .ip(n4712), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[27]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_28_ ( .ip(n4711), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[28]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_29_ ( .ip(n4710), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[29]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_30_ ( .ip(n4709), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[30]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_31_ ( .ip(n4708), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[31]) );
  drp_1 i_ssi_U_biu_prdata_reg_16_ ( .ip(n4228), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[16]) );
  drp_1 i_ssi_U_biu_prdata_reg_17_ ( .ip(n4227), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[17]) );
  drp_1 i_ssi_U_biu_prdata_reg_18_ ( .ip(n4226), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[18]) );
  drp_1 i_ssi_U_biu_prdata_reg_19_ ( .ip(n4225), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[19]) );
  drp_1 i_ssi_U_biu_prdata_reg_20_ ( .ip(n4224), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[20]) );
  drp_1 i_ssi_U_biu_prdata_reg_21_ ( .ip(n4223), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[21]) );
  drp_1 i_ssi_U_biu_prdata_reg_22_ ( .ip(n4222), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[22]) );
  drp_1 i_ssi_U_biu_prdata_reg_23_ ( .ip(n4221), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[23]) );
  drp_1 i_ssi_U_biu_prdata_reg_24_ ( .ip(n4220), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[24]) );
  drp_1 i_ssi_U_biu_prdata_reg_25_ ( .ip(n4219), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[25]) );
  drp_1 i_ssi_U_biu_prdata_reg_26_ ( .ip(n4218), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[26]) );
  drp_1 i_ssi_U_biu_prdata_reg_27_ ( .ip(n4217), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[27]) );
  drp_1 i_ssi_U_biu_prdata_reg_28_ ( .ip(n4216), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[28]) );
  drp_1 i_ssi_U_biu_prdata_reg_29_ ( .ip(n4215), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[29]) );
  drp_1 i_ssi_U_biu_prdata_reg_30_ ( .ip(n4214), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[30]) );
  drp_1 i_ssi_U_biu_prdata_reg_31_ ( .ip(n4213), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[31]) );
  drp_1 i_ssi_U_regfile_ser_reg_0_ ( .ip(n4634), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_ser_0_) );
  drp_1 i_ssi_U_regfile_rxftlr_reg_0_ ( .ip(n4644), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_rxftlr[0]) );
  drp_1 i_ssi_U_regfile_rxftlr_reg_1_ ( .ip(n4643), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_rxftlr[1]) );
  drp_1 i_ssi_U_regfile_rxftlr_reg_2_ ( .ip(n4642), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_rxftlr[2]) );
  drp_1 i_ssi_U_regfile_txftlr_reg_0_ ( .ip(n4641), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_txftlr[0]) );
  drp_1 i_ssi_U_regfile_txftlr_reg_1_ ( .ip(n4640), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_txftlr[1]) );
  drp_1 i_ssi_U_regfile_txftlr_reg_2_ ( .ip(n4639), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_txftlr[2]) );
  drp_1 i_ssi_U_regfile_ssienr_reg ( .ip(n4638), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_ssi_en_int) );
  drp_1 i_ssi_U_regfile_mwcr_ir_reg_2_ ( .ip(n4635), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_mwcr[2]) );
  drp_1 i_ssi_U_regfile_baudr_reg_7_ ( .ip(n4627), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[7]) );
  drp_1 i_ssi_U_regfile_baudr_reg_8_ ( .ip(n4626), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[8]) );
  drp_1 i_ssi_U_regfile_baudr_reg_9_ ( .ip(n4625), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[9]) );
  drp_1 i_ssi_U_regfile_baudr_reg_11_ ( .ip(n4623), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[11]) );
  drp_1 i_ssi_U_regfile_baudr_reg_13_ ( .ip(n4621), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[13]) );
  drp_1 i_ssi_U_regfile_baudr_reg_15_ ( .ip(n4619), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[15]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_0_ ( .ip(n4610), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[0]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_2_ ( .ip(n4608), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[2]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_3_ ( .ip(n4607), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[3]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_4_ ( .ip(n4606), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[4]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_5_ ( .ip(n4605), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[5]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_6_ ( .ip(n4604), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[6]) );
  drp_1 i_ssi_U_biu_prdata_reg_7_ ( .ip(n4237), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[7]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_8_ ( .ip(n4618), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[8]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_9_ ( .ip(n4617), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[9]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_4_ ( .ip(n4592), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr0_ir_int[4]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_5_ ( .ip(n4593), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr0_ir_int[5]) );
  drp_1 i_ssi_U_regfile_sclk_active_reg ( .ip(n5242), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_sclk_active) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_8_ ( .ip(n4595), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_tmod[0]) );
  drp_1 i_ssi_U_biu_prdata_reg_8_ ( .ip(n4236), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[8]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_9_ ( .ip(n4596), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_tmod[1]) );
  drp_1 i_ssi_U_biu_prdata_reg_9_ ( .ip(n4235), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[9]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_10_ ( .ip(n4597), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_ctrlr0[10]) );
  drp_1 i_ssi_U_biu_prdata_reg_10_ ( .ip(n4234), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[10]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_11_ ( .ip(n4598), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_ctrlr0[11]) );
  drp_1 i_ssi_U_biu_prdata_reg_11_ ( .ip(n4233), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[11]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_12_ ( .ip(n4599), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_cfs[0]) );
  drp_1 i_ssi_U_biu_prdata_reg_12_ ( .ip(n4232), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[12]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_13_ ( .ip(n4600), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_cfs[1]) );
  drp_1 i_ssi_U_biu_prdata_reg_13_ ( .ip(n4231), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[13]) );
  drp_1 i_ssi_U_biu_prdata_reg_14_ ( .ip(n4230), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[14]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_15_ ( .ip(n4602), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_cfs[3]) );
  drp_1 i_ssi_U_biu_prdata_reg_15_ ( .ip(n4229), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[15]) );
  drp_1 i_ssi_U_sclkgen_sclk_fe_ir_reg ( .ip(i_ssi_U_sclkgen_N75), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_sclk_fe) );
  drp_1 i_ssi_U_fifo_tx_push_dly_reg ( .ip(n11780), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_fifo_tx_push_dly) );
  drp_1 i_ssi_U_fifo_rx_pop_dly_reg ( .ip(n11782), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_fifo_rx_pop_dly) );
  drp_1 i_ssi_U_mstfsm_U_ss_in_n_sync_sample_meta_reg_0_ ( .ip(i_ssi_ss_in_n), 
        .ck(i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_mstfsm_U_ss_in_n_sync_next_sample_syncm1_0_) );
  drp_1 i_ssi_U_mstfsm_U_ss_in_n_sync_sample_syncl_reg_0_ ( .ip(
        i_ssi_U_mstfsm_U_ss_in_n_sync_next_sample_syncm1_0_), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_ss_in_n_sync)
         );
  drp_1 i_ssi_U_mstfsm_c_state_reg_1_ ( .ip(i_ssi_U_mstfsm_N221), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_c_state[1]) );
  drp_1 i_ssi_U_mstfsm_c_state_reg_3_ ( .ip(i_ssi_U_mstfsm_N223), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_c_state[3]) );
  drp_1 i_ssi_U_mstfsm_c_done_ir_reg ( .ip(n4587), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_c_done_ir) );
  drp_1 i_ssi_U_mstfsm_last_frame_reg ( .ip(n4429), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_last_frame) );
  drp_1 i_ssi_U_mstfsm_abort_ir_reg ( .ip(n4428), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_abort_ir) );
  drp_1 i_ssi_U_fifo_tx_pop_edge_reg ( .ip(i_ssi_tx_pop), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_fifo_tx_pop_edge) );
  drp_1 i_ssi_U_fifo_tx_pop_sync_dly_reg ( .ip(i_ssi_tx_pop_sync), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_ssi_U_fifo_tx_pop_sync_dly) );
  drp_1 i_ssi_U_intctl_irisr_tx_empty_reg ( .ip(i_ssi_U_intctl_N2), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_ssi_risr[0]) );
  drp_1 i_ssi_U_intctl_irisr_tx_fifo_overflow_reg ( .ip(n4584), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_ssi_risr[1]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__0_ ( .ip(n4583), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[0]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__1_ ( .ip(n4582), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[1]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__2_ ( .ip(n4581), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[2]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__3_ ( .ip(n4580), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[3]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__4_ ( .ip(n4579), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[4]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__5_ ( .ip(n4578), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[5]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__6_ ( .ip(n4577), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[6]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__7_ ( .ip(n4576), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[7]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__8_ ( .ip(n4575), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[8]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__9_ ( .ip(n4574), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[9]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__10_ ( .ip(n4573), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[10]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__11_ ( .ip(n4572), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[11]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__12_ ( .ip(n4571), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[12]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__13_ ( .ip(n4570), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[13]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__14_ ( .ip(n4569), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[14]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__15_ ( .ip(n4568), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[15]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__0_ ( .ip(n4551), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[32]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__1_ ( .ip(n4550), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[33]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__2_ ( .ip(n4549), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[34]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__3_ ( .ip(n4548), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[35]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__4_ ( .ip(n4547), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[36]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__5_ ( .ip(n4546), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[37]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__6_ ( .ip(n4545), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[38]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__7_ ( .ip(n4544), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[39]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__8_ ( .ip(n4543), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[40]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__9_ ( .ip(n4542), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[41]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__10_ ( .ip(n4541), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[42]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__11_ ( .ip(n4540), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[43]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__12_ ( .ip(n4539), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[44]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__13_ ( .ip(n4538), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[45]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__14_ ( .ip(n4537), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[46]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__15_ ( .ip(n4536), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[47]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__0_ ( .ip(n4519), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[64]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__1_ ( .ip(n4518), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[65]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__2_ ( .ip(n4517), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[66]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__3_ ( .ip(n4516), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[67]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__4_ ( .ip(n4515), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[68]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__5_ ( .ip(n4514), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[69]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__6_ ( .ip(n4513), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[70]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__7_ ( .ip(n4512), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[71]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__8_ ( .ip(n4511), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[72]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__9_ ( .ip(n4510), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[73]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__10_ ( .ip(n4509), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[74]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__11_ ( .ip(n4508), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[75]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__12_ ( .ip(n4507), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[76]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__13_ ( .ip(n4506), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[77]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__14_ ( .ip(n4505), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[78]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__15_ ( .ip(n4504), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[79]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__0_ ( .ip(n4487), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[96]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__1_ ( .ip(n4486), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[97]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__2_ ( .ip(n4485), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[98]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__3_ ( .ip(n4484), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[99]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__4_ ( .ip(n4483), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[100]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__5_ ( .ip(n4482), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[101]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__6_ ( .ip(n4481), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[102]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__7_ ( .ip(n4480), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[103]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__8_ ( .ip(n4479), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[104]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__9_ ( .ip(n4478), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[105]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__10_ ( .ip(n4477), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[106]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__11_ ( .ip(n4476), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[107]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__12_ ( .ip(n4475), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[108]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__13_ ( .ip(n4474), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[109]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__14_ ( .ip(n4473), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[110]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__15_ ( .ip(n4472), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[111]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__0_ ( .ip(n4567), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[16]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__1_ ( .ip(n4566), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[17]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__2_ ( .ip(n4565), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[18]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__3_ ( .ip(n4564), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[19]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__4_ ( .ip(n4563), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[20]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__5_ ( .ip(n4562), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[21]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__6_ ( .ip(n4561), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[22]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__7_ ( .ip(n4560), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[23]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__8_ ( .ip(n4559), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[24]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__9_ ( .ip(n4558), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[25]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__10_ ( .ip(n4557), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[26]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__11_ ( .ip(n4556), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[27]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__12_ ( .ip(n4555), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[28]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__13_ ( .ip(n4554), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[29]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__14_ ( .ip(n4553), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[30]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__15_ ( .ip(n4552), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[31]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__0_ ( .ip(n4535), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[48]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__1_ ( .ip(n4534), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[49]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__2_ ( .ip(n4533), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[50]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__3_ ( .ip(n4532), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[51]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__4_ ( .ip(n4531), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[52]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__5_ ( .ip(n4530), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[53]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__6_ ( .ip(n4529), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[54]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__7_ ( .ip(n4528), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[55]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__8_ ( .ip(n4527), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[56]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__9_ ( .ip(n4526), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[57]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__10_ ( .ip(n4525), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[58]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__11_ ( .ip(n4524), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[59]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__12_ ( .ip(n4523), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[60]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__13_ ( .ip(n4522), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[61]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__14_ ( .ip(n4521), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[62]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__15_ ( .ip(n4520), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[63]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__0_ ( .ip(n4503), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[80]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__1_ ( .ip(n4502), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[81]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__2_ ( .ip(n4501), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[82]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__3_ ( .ip(n4500), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[83]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__4_ ( .ip(n4499), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[84]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__5_ ( .ip(n4498), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[85]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__6_ ( .ip(n4497), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[86]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__7_ ( .ip(n4496), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[87]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__8_ ( .ip(n4495), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[88]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__9_ ( .ip(n4494), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[89]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__10_ ( .ip(n4493), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[90]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__11_ ( .ip(n4492), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[91]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__12_ ( .ip(n4491), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[92]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__13_ ( .ip(n4490), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[93]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__14_ ( .ip(n4489), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[94]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__15_ ( .ip(n4488), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[95]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__0_ ( .ip(n4471), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[112]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__1_ ( .ip(n4470), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[113]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__2_ ( .ip(n4469), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[114]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__3_ ( .ip(n4468), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[115]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__4_ ( .ip(n4467), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[116]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__5_ ( .ip(n4466), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[117]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__6_ ( .ip(n4465), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[118]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__7_ ( .ip(n4464), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[119]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__8_ ( .ip(n4463), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[120]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__9_ ( .ip(n4462), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[121]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__10_ ( .ip(n4461), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[122]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__11_ ( .ip(n4460), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[123]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__12_ ( .ip(n4459), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[124]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__13_ ( .ip(n4458), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[125]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__14_ ( .ip(n4457), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[126]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__15_ ( .ip(n4456), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[127]) );
  drp_1 i_ssi_U_regfile_txflr_reg_0_ ( .ip(n4454), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_txflr[0]) );
  drp_1 i_ssi_U_regfile_txflr_reg_1_ ( .ip(n4453), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_txflr[1]) );
  drp_1 i_ssi_U_regfile_txflr_reg_2_ ( .ip(n4452), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_txflr[2]) );
  drp_1 i_ssi_U_regfile_txflr_reg_3_ ( .ip(n4455), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_txflr[3]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_load_start_bit_ir_reg ( .ip(
        i_ssi_load_start_bit), .ck(i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_load_start_bit_ir) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_0_ ( .ip(n4427), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[0]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_1_ ( .ip(n4426), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[1]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_2_ ( .ip(n4425), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[2]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_3_ ( .ip(n4424), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[3]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_4_ ( .ip(n4423), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[4]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_5_ ( .ip(n4422), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[5]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_6_ ( .ip(n4421), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[6]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_7_ ( .ip(n4420), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[7]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_8_ ( .ip(n4419), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[8]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_9_ ( .ip(n4418), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[9]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_10_ ( .ip(n4417), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[10]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_11_ ( .ip(n4416), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[11]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_12_ ( .ip(n4415), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[12]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_13_ ( .ip(n4414), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[13]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_14_ ( .ip(n4413), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[14]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_15_ ( .ip(n4412), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[15]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_1_ ( .ip(n4409), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[1]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_5_ ( .ip(n4405), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[5]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_8_ ( .ip(n4402), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[8]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_0_ ( .ip(n4394), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[0]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_1_ ( .ip(n4393), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[1]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_2_ ( .ip(n4392), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[2]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_3_ ( .ip(n4391), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[3]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_4_ ( .ip(n4390), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[4]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_5_ ( .ip(n4389), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[5]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_6_ ( .ip(n4388), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[6]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_7_ ( .ip(n4387), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[7]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_8_ ( .ip(n4386), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[8]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_9_ ( .ip(n4385), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[9]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_10_ ( .ip(n4384), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[10]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_11_ ( .ip(n4383), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[11]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_12_ ( .ip(n4382), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[12]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_13_ ( .ip(n4381), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[13]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_14_ ( .ip(n4380), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[14]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_15_ ( .ip(n4379), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[15]) );
  drp_1 i_ssi_U_fifo_rx_push_edge_reg ( .ip(i_ssi_rx_push), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_ssi_U_fifo_rx_push_edge) );
  drp_1 i_ssi_U_fifo_rx_push_sync_dly_reg ( .ip(n11760), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_fifo_rx_push_sync_dly) );
  drp_1 i_ssi_U_intctl_irisr_rx_full_reg ( .ip(i_ssi_U_intctl_N33), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_ssi_risr[4]) );
  drp_1 i_ssi_U_biu_prdata_reg_4_ ( .ip(n4240), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[4]) );
  drp_1 i_ssi_U_intctl_irisr_rx_fifo_overflow_reg ( .ip(n4450), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_ssi_risr[3]) );
  drp_1 i_ssi_U_intctl_irisr_rx_fifo_underflow_reg ( .ip(n4449), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(i_ssi_risr[2]) );
  drp_1 i_ssi_U_regfile_rxflr_reg_0_ ( .ip(n4447), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_rxflr[0]) );
  drp_1 i_ssi_U_regfile_rxflr_reg_1_ ( .ip(n4446), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_rxflr[1]) );
  drp_1 i_ssi_U_biu_prdata_reg_1_ ( .ip(n4243), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[1]) );
  drp_1 i_ssi_U_regfile_rxflr_reg_2_ ( .ip(n4445), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_rxflr[2]) );
  drp_1 i_ssi_U_regfile_rxflr_reg_3_ ( .ip(n4448), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_rxflr[3]) );
  drp_1 i_ssi_U_biu_prdata_reg_3_ ( .ip(n4241), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[3]) );
  drp_1 i_ssi_U_biu_prdata_reg_2_ ( .ip(n4242), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[2]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_1_ ( .ip(n4444), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[1]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__1_ ( .ip(n4369), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[1]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__1_ ( .ip(n4368), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[17]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__1_ ( .ip(n4367), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[33]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__1_ ( .ip(n4366), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[49]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__1_ ( .ip(n4365), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[65]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__1_ ( .ip(n4364), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[81]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__1_ ( .ip(n4363), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[97]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__1_ ( .ip(n4362), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[113]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_2_ ( .ip(n4443), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[2]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__2_ ( .ip(n4361), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[2]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__2_ ( .ip(n4360), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[18]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__2_ ( .ip(n4359), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[34]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__2_ ( .ip(n4358), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[50]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__2_ ( .ip(n4357), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[66]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__2_ ( .ip(n4356), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[82]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__2_ ( .ip(n4355), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[98]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__2_ ( .ip(n4354), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[114]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_3_ ( .ip(n4442), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[3]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__3_ ( .ip(n4353), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[3]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__3_ ( .ip(n4352), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[19]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__3_ ( .ip(n4351), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[35]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__3_ ( .ip(n4350), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[51]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__3_ ( .ip(n4349), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[67]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__3_ ( .ip(n4348), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[83]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__3_ ( .ip(n4347), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[99]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__3_ ( .ip(n4346), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[115]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_4_ ( .ip(n4441), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[4]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__4_ ( .ip(n4345), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[4]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__4_ ( .ip(n4344), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[20]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__4_ ( .ip(n4343), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[36]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__4_ ( .ip(n4342), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[52]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__4_ ( .ip(n4341), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[68]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__4_ ( .ip(n4340), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[84]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__4_ ( .ip(n4339), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[100]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__4_ ( .ip(n4338), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[116]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_5_ ( .ip(n4440), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[5]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__5_ ( .ip(n4337), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[5]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__5_ ( .ip(n4336), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[21]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__5_ ( .ip(n4335), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[37]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__5_ ( .ip(n4334), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[53]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__5_ ( .ip(n4333), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[69]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__5_ ( .ip(n4332), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[85]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__5_ ( .ip(n4331), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[101]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__5_ ( .ip(n4330), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[117]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_6_ ( .ip(n4439), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[6]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__6_ ( .ip(n4329), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[6]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__6_ ( .ip(n4328), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[22]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__6_ ( .ip(n4327), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[38]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__6_ ( .ip(n4326), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[54]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__6_ ( .ip(n4325), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[70]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__6_ ( .ip(n4324), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[86]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__6_ ( .ip(n4323), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[102]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__6_ ( .ip(n4322), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[118]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_7_ ( .ip(n4438), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[7]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__7_ ( .ip(n4321), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[7]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__7_ ( .ip(n4320), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[23]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__7_ ( .ip(n4319), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[39]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__7_ ( .ip(n4318), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[55]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__7_ ( .ip(n4317), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[71]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__7_ ( .ip(n4316), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[87]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__7_ ( .ip(n4315), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[103]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__7_ ( .ip(n4314), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[119]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_8_ ( .ip(n4437), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[8]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__8_ ( .ip(n4313), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[8]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__8_ ( .ip(n4312), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[24]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__8_ ( .ip(n4311), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[40]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__8_ ( .ip(n4310), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[56]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__8_ ( .ip(n4309), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[72]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__8_ ( .ip(n4308), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[88]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__8_ ( .ip(n4307), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[104]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__8_ ( .ip(n4306), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[120]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_9_ ( .ip(n4436), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[9]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__9_ ( .ip(n4305), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[9]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__9_ ( .ip(n4304), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[25]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__9_ ( .ip(n4303), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[41]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__9_ ( .ip(n4302), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[57]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__9_ ( .ip(n4301), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[73]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__9_ ( .ip(n4300), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[89]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__9_ ( .ip(n4299), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[105]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__9_ ( .ip(n4298), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[121]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_10_ ( .ip(n4435), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[10]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__10_ ( .ip(n4297), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[10]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__10_ ( .ip(n4296), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[26]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__10_ ( .ip(n4295), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[42]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__10_ ( .ip(n4294), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[58]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__10_ ( .ip(n4293), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[74]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__10_ ( .ip(n4292), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[90]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__10_ ( .ip(n4291), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[106]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__10_ ( .ip(n4290), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[122]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_11_ ( .ip(n4434), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[11]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__11_ ( .ip(n4289), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[11]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__11_ ( .ip(n4288), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[27]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__11_ ( .ip(n4287), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[43]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__11_ ( .ip(n4286), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[59]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__11_ ( .ip(n4285), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[75]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__11_ ( .ip(n4284), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[91]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__11_ ( .ip(n4283), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[107]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__11_ ( .ip(n4282), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[123]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_12_ ( .ip(n4433), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[12]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__12_ ( .ip(n4281), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[12]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__12_ ( .ip(n4280), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[28]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__12_ ( .ip(n4279), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[44]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__12_ ( .ip(n4278), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[60]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__12_ ( .ip(n4277), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[76]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__12_ ( .ip(n4276), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[92]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__12_ ( .ip(n4275), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[108]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__12_ ( .ip(n4274), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[124]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_13_ ( .ip(n4432), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[13]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__13_ ( .ip(n4273), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[13]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__13_ ( .ip(n4272), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[29]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__13_ ( .ip(n4271), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[45]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__13_ ( .ip(n4270), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[61]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__13_ ( .ip(n4269), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[77]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__13_ ( .ip(n4268), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[93]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__13_ ( .ip(n4267), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[109]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__13_ ( .ip(n4266), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[125]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_14_ ( .ip(n4431), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[14]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__14_ ( .ip(n4265), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[14]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__14_ ( .ip(n4264), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[30]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__14_ ( .ip(n4263), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[46]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__14_ ( .ip(n4262), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[62]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__14_ ( .ip(n4261), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[78]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__14_ ( .ip(n4260), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[94]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__14_ ( .ip(n4259), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[110]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__14_ ( .ip(n4258), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[126]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_15_ ( .ip(n4430), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[15]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__15_ ( .ip(n4257), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[15]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__15_ ( .ip(n4256), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[31]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__15_ ( .ip(n4255), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[47]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__15_ ( .ip(n4254), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[63]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__15_ ( .ip(n4253), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[79]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__15_ ( .ip(n4252), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[95]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__15_ ( .ip(n4251), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[111]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__15_ ( .ip(n4250), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[127]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_0_ ( .ip(n4378), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[0]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__0_ ( .ip(n4377), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[0]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__0_ ( .ip(n4376), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[16]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__0_ ( .ip(n4375), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[32]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__0_ ( .ip(n4374), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[48]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__0_ ( .ip(n4373), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[64]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__0_ ( .ip(n4372), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[80]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__0_ ( .ip(n4371), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[96]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__0_ ( .ip(n4370), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[112]) );
  drp_1 i_ssi_U_regfile_ssi_sleep_ir_reg ( .ip(i_ssi_U_regfile_N451), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_ssi_ssi_sleep) );
  drp_1 i_ssi_U_mstfsm_fsm_busy_reg ( .ip(n11778), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_fsm_busy) );
  drp_1 i_ssi_U_regfile_multi_mst_edge_reg ( .ip(i_ssi_fsm_multi_mst), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_ssi_U_regfile_multi_mst_edge)
         );
  drp_1 i_ssi_U_intctl_irisr_mst_collision_reg ( .ip(n4247), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_ssi_risr[5]) );
  drp_1 i_ssi_U_biu_prdata_reg_0_ ( .ip(n4244), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[0]) );
  drp_1 i_ssi_U_biu_prdata_reg_5_ ( .ip(n4239), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[5]) );
  drp_1 i_ssi_U_intctl_mst_contention_reg ( .ip(n4246), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_mst_contention) );
  drp_1 i_ssi_U_regfile_i_sr_reg ( .ip(n4245), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_sr_6_) );
  drp_1 i_ssi_U_biu_prdata_reg_6_ ( .ip(n4238), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_U_SYNC_sample_meta_reg_0_ ( 
        .ip(i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_U_SYNC_N2), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_U_SYNC_next_sample_syncm1_0_)
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_U_SYNC_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_U_SYNC_next_sample_syncm1_0_), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_data_d_int_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_U_SYNC_sample_meta_reg_0_ ( 
        .ip(i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_U_SYNC_N2), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_U_SYNC_next_sample_syncm1_0_)
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_U_SYNC_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_U_SYNC_next_sample_syncm1_0_), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_data_d_int_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_mst_arb_lost_reg ( .ip(n4939), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_mst_arb_lost) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_12_ ( 
        .ip(i_i2c_tx_abrt_source[12]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_12_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[12]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_12_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[12]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_mst_gen_ack_en_r_reg ( .ip(n11770), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_mst_gen_ack_en_r) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_ic_data_oe_early_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_N85), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_tx_shift_ic_data_oe_early) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_ic_data_oe_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_ic_data_oe_early), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_ic_data_oe) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_ic_rd_req_tog_reg ( .ip(n5037), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ic_rd_req_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_ic_rd_req_flg_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_ic_rd_req_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_ic_rd_req_flg_sync_next_sample_syncm1_0_)
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_ic_rd_req_flg_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_ic_rd_req_flg_sync_next_sample_syncm1_0_), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_ic_rd_req_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_rd_req_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_ic_rd_req_flg_sync), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_DW_apb_i2c_intctl_ic_rd_req_flg_sync_q)
         );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_mst_tx_flush_reg ( .ip(n4864), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_mst_tx_flush) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_sbyte_norstrt_tog_reg ( .ip(n4861), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_9_ ( 
        .ip(i_i2c_tx_abrt_source[9]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[9])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_9_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[9]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_9_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[9]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_9_ ( .ip(n4698), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_gen_call_sample_meta_reg_0_ ( .ip(
        i_i2c_ic_ack_general_call), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_U_DW_apb_i2c_sync_U_ic_gen_call_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_gen_call_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_gen_call_next_sample_syncm1_0_), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ic_ack_general_call_sync)
         );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_ic_sda_hold[0]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[0]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_1_ ( .ip(
        i_i2c_ic_sda_hold[1]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_2_ ( .ip(
        i_i2c_ic_sda_hold[2]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[2]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_3_ ( .ip(
        i_i2c_ic_sda_hold[3]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_3_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[3]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_4_ ( .ip(
        i_i2c_ic_sda_hold[4]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_4_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[4]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_5_ ( .ip(
        i_i2c_ic_sda_hold[5]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_5_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[5]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_6_ ( .ip(
        i_i2c_ic_sda_hold[6]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_6_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[6]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_7_ ( .ip(
        i_i2c_ic_sda_hold[7]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_7_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[7]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_8_ ( .ip(
        i_i2c_ic_sda_hold[8]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_8_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[8]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_9_ ( .ip(
        i_i2c_ic_sda_hold[9]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_9_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[9]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_10_ ( .ip(
        i_i2c_ic_sda_hold[10]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_10_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[10]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_11_ ( .ip(
        i_i2c_ic_sda_hold[11]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_11_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[11]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_12_ ( .ip(
        i_i2c_ic_sda_hold[12]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_12_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[12]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_13_ ( .ip(
        i_i2c_ic_sda_hold[13]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_13_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[13]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_14_ ( .ip(
        i_i2c_ic_sda_hold[14]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_14_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[14]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_15_ ( .ip(
        i_i2c_ic_sda_hold[15]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_15_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[15]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_16_ ( .ip(
        i_i2c_ic_sda_hold[16]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[16]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_16_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[16]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_rx_hold_sync[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_17_ ( .ip(
        i_i2c_ic_sda_hold[17]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[17]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_17_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[17]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_rx_hold_sync[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_18_ ( .ip(
        i_i2c_ic_sda_hold[18]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[18]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_18_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[18]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_rx_hold_sync[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_19_ ( .ip(
        i_i2c_ic_sda_hold[19]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[19]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_19_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[19]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_rx_hold_sync[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_20_ ( .ip(
        i_i2c_ic_sda_hold[20]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[20]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_20_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[20]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_rx_hold_sync[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_21_ ( .ip(
        i_i2c_ic_sda_hold[21]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[21]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_21_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[21]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_rx_hold_sync[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_22_ ( .ip(
        i_i2c_ic_sda_hold[22]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[22]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_22_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[22]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_rx_hold_sync[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_23_ ( .ip(
        i_i2c_ic_sda_hold[23]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[23]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_23_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[23]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_rx_hold_sync[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_rstrt_en_1_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_rstrt_en_1_sync_N2), .ck(i_i2c_ic_clk), 
        .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_rstrt_en_1_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_rstrt_en_1_sync_sample_syncl_reg_0_ ( 
        .ip(i_i2c_U_DW_apb_i2c_sync_U_ic_rstrt_en_1_sync_next_sample_syncm1_0_), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_ic_rstrt_en_sync_inv) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_push_dly_reg ( .ip(i_i2c_tx_push), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_push_dly) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_rx_pop_dly_reg ( .ip(i_i2c_rx_pop), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_rx_pop_dly) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_p_det_ifaddr_sample_meta_reg_0_ ( .ip(
        i_i2c_p_det_ifaddr), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_p_det_ifaddr_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_p_det_ifaddr_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_p_det_ifaddr_next_sample_syncm1_0_), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_p_det_ifaddr_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_slave_en_1_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_ic_slave_en), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_slave_en_1_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_slave_en_1_sync_sample_syncl_reg_0_ ( 
        .ip(i_i2c_U_DW_apb_i2c_sync_U_ic_slave_en_1_sync_next_sample_syncm1_0_), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ic_slave_en_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_slv_1_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_slv_1_sync_N2), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_slv_1_sync_next_sample_syncm1_0_)
         );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_slv_1_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_slv_1_sync_next_sample_syncm1_0_), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_ic_10bit_slv_sync_inv) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_mst_1_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_mst_1_sync_N2), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_mst_1_sync_next_sample_syncm1_0_)
         );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_mst_1_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_mst_1_sync_next_sample_syncm1_0_), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_ic_10bit_mst_sync_inv) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_master_1_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_master_1_sync_N2), .ck(i_i2c_ic_clk), 
        .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_master_1_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_master_1_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_master_1_sync_next_sample_syncm1_0_), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_master_dis_tog_reg ( .ip(n4862), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_11_ ( 
        .ip(i_i2c_tx_abrt_source[11]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_11_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[11]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_11_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[11]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_ss_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_ic_ss), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_ss_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_ss_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_ss_sync_next_sample_syncm1_0_), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ic_ss_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_fs_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_ic_fs), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_fs_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_fs_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_fs_sync_next_sample_syncm1_0_), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ic_fs_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_hs_sync_sample_meta_reg_0_ ( .ip(n11763), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_hs_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_hs_norstrt_tog_reg ( .ip(n4863), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_8_ ( 
        .ip(i_i2c_tx_abrt_source[8]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[8])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_8_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[8]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_8_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[8]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_enable_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_ic_enable[0]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_enable_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_enable_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_enable_sync_next_sample_syncm1_0_), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ic_enable_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_ic_bus_idle_reg ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N51), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ic_bus_idle) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_abort_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_ic_enable[1]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_abort_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_abort_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_abort_sync_next_sample_syncm1_0_), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ic_abort_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_sync_d_reg ( .ip(
        i_i2c_ic_abort_sync), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_sync_d) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_split_start_en_int_reg ( .ip(n5232), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_split_start_en) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_start_en_int_reg ( .ip(n5117), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_start_en) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_st_scl_s_hld_en_reg ( .ip(i_i2c_start_en), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_st_scl_s_hld_en) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cmplt_reg ( .ip(n5195), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_scl_s_hld_cmplt) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl_lcnt_en_reg ( .ip(n4962), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl_lcnt_en) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_lcnt_cmplt_reg ( .ip(n5200), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_scl_lcnt_cmplt) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_re_start_en_int_reg ( .ip(n5199), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_re_start_en) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_s_gen_reg ( .ip(
        i_i2c_U_DW_apb_i2c_toggle_N30), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_s_gen) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_byte_wait_scl_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_byte_wait_en), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_byte_wait_scl) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_rd_reg ( .ip(n11773), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_debug_rd) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_bit_count_reg_1_ ( .ip(n5115), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_mst_rx_bit_count[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_ack_int_reg ( .ip(n4959), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_mst_rx_ack_vld) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rxbyte_rdy_reg ( .ip(n4938), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_mst_rxbyte_rdy) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_byte_waiting_q_reg ( .ip(n5191), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_byte_waiting_q) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_mst_current_state_reg_3_ ( .ip(
        i_i2c_U_DW_apb_i2c_mstfsm_N75), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_mst_debug_cstate[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_mst_cstate_reg_3_ ( .ip(
        i_i2c_mst_debug_cstate[3]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_mst_cstate[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_mst_activity_reg ( .ip(
        i_i2c_U_DW_apb_i2c_mstfsm_N487), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_mst_activity) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_master_act_reg ( .ip(
        i_i2c_mst_activity), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_debug_master_act) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_mst_activity_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_mst_activity), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_mst_activity_sync_next_sample_syncm1_0_)
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_mst_activity_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_mst_activity_sync_next_sample_syncm1_0_), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_mst_activity_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_mst_current_state_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_mstfsm_N72), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_mst_debug_cstate[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_mst_cstate_reg_0_ ( .ip(
        i_i2c_mst_debug_cstate[0]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_mst_cstate[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_mst_current_state_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_mstfsm_N73), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_mst_debug_cstate[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_mst_cstate_reg_1_ ( .ip(
        i_i2c_mst_debug_cstate[1]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_mst_cstate[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_mst_current_state_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_mstfsm_N74), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_mst_debug_cstate[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_mst_cstate_reg_2_ ( .ip(
        i_i2c_mst_debug_cstate[2]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_mst_cstate[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_addr_2byte_sent_reg ( .ip(n5206), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_addr_2byte_sent) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_pop_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_tx_pop) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_pop_flg_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_tx_pop_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_pop_flg_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_pop_flg_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_pop_flg_sync_next_sample_syncm1_0_), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_pop_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_pop_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_tx_pop_flg_sync), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_DW_apb_i2c_fifo_tx_pop_flg_sync_q) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_pop_sync_dly_reg ( .ip(i_i2c_tx_pop_sync), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_pop_sync_dly) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_tx_empty_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_empty_n), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_tx_empty_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_tx_empty_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_tx_empty_sync_next_sample_syncm1_0_), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_tx_empty_int_inv) );
  drp_1 i_i2c_U_dff_tx_mem_reg_7__0_ ( .ip(n5035), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[0]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_7__1_ ( .ip(n5027), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[1]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_7__2_ ( .ip(n5019), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[2]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_7__3_ ( .ip(n5011), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[3]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_7__4_ ( .ip(n5003), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[4]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_7__5_ ( .ip(n4995), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[5]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_7__6_ ( .ip(n4987), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[6]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_7__7_ ( .ip(n4979), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[7]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_7__8_ ( .ip(n4971), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[8]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_5__0_ ( .ip(n5033), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[18]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_5__1_ ( .ip(n5025), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[19]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_5__2_ ( .ip(n5017), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[20]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_5__3_ ( .ip(n5009), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[21]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_5__4_ ( .ip(n5001), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[22]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_5__5_ ( .ip(n4993), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[23]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_5__6_ ( .ip(n4985), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[24]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_5__7_ ( .ip(n4977), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[25]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_5__8_ ( .ip(n4969), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[26]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_3__0_ ( .ip(n5031), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[36]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_3__1_ ( .ip(n5023), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[37]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_3__2_ ( .ip(n5015), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[38]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_3__3_ ( .ip(n5007), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[39]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_3__4_ ( .ip(n4999), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[40]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_3__5_ ( .ip(n4991), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[41]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_3__6_ ( .ip(n4983), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[42]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_3__7_ ( .ip(n4975), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[43]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_3__8_ ( .ip(n4967), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[44]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_1__0_ ( .ip(n5029), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[54]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_1__1_ ( .ip(n5021), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[55]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_1__2_ ( .ip(n5013), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[56]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_1__3_ ( .ip(n5005), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[57]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_1__4_ ( .ip(n4997), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[58]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_1__5_ ( .ip(n4989), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[59]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_1__6_ ( .ip(n4981), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[60]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_1__7_ ( .ip(n4973), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[61]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_1__8_ ( .ip(n4965), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[62]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_6__0_ ( .ip(n5034), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[9]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_6__1_ ( .ip(n5026), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[10]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_6__2_ ( .ip(n5018), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[11]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_6__3_ ( .ip(n5010), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[12]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_6__4_ ( .ip(n5002), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[13]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_6__5_ ( .ip(n4994), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[14]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_6__6_ ( .ip(n4986), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[15]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_6__7_ ( .ip(n4978), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[16]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_6__8_ ( .ip(n4970), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[17]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_4__0_ ( .ip(n5032), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[27]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_4__1_ ( .ip(n5024), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[28]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_4__2_ ( .ip(n5016), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[29]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_4__3_ ( .ip(n5008), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[30]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_4__4_ ( .ip(n5000), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[31]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_4__5_ ( .ip(n4992), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[32]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_4__6_ ( .ip(n4984), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[33]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_4__7_ ( .ip(n4976), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[34]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_4__8_ ( .ip(n4968), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[35]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_2__0_ ( .ip(n5030), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[45]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_2__1_ ( .ip(n5022), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[46]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_2__2_ ( .ip(n5014), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[47]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_2__3_ ( .ip(n5006), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[48]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_2__4_ ( .ip(n4998), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[49]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_2__5_ ( .ip(n4990), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[50]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_2__6_ ( .ip(n4982), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[51]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_2__7_ ( .ip(n4974), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[52]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_2__8_ ( .ip(n4966), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[53]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_0__0_ ( .ip(n5028), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[63]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_0__1_ ( .ip(n5020), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[64]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_0__2_ ( .ip(n5012), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[65]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_0__3_ ( .ip(n5004), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[66]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_0__4_ ( .ip(n4996), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[67]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_0__5_ ( .ip(n4988), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[68]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_0__6_ ( .ip(n4980), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[69]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_0__7_ ( .ip(n4972), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[70]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_0__8_ ( .ip(n4964), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[71]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_fifo_data_buf_reg_0_ ( .ip(n5229), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_fifo_data_buf[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_fifo_data_buf_reg_1_ ( .ip(n5228), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_fifo_data_buf[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_fifo_data_buf_reg_2_ ( .ip(n5227), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_fifo_data_buf[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_fifo_data_buf_reg_3_ ( .ip(n5226), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_fifo_data_buf[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_fifo_data_buf_reg_4_ ( .ip(n5225), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_fifo_data_buf[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_fifo_data_buf_reg_5_ ( .ip(n5224), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_fifo_data_buf[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_fifo_data_buf_reg_6_ ( .ip(n5223), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_fifo_data_buf[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_fifo_data_buf_reg_7_ ( .ip(n5222), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_fifo_data_buf[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_fifo_data_buf_reg_8_ ( .ip(n5221), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_fifo_data_buf[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_data_capture_reg ( .ip(n11772), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_debug_wr) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_scl_p_stp_int_reg ( .ip(n5068), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_scl_p_setup_en) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cmplt_reg ( .ip(n5051), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_scl_p_setup_cmplt) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_mst_current_state_reg_4_ ( .ip(
        i_i2c_U_DW_apb_i2c_mstfsm_N76), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_mst_debug_cstate[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_mst_cstate_reg_4_ ( .ip(
        i_i2c_mst_debug_cstate[4]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_mst_cstate[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_abrt_in_rcve_trns_reg ( .ip(n5190), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_abrt_in_rcve_trns) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_addr_1byte_sent_reg ( .ip(n5207), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_addr_1byte_sent) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_delay_stop_en_reg ( .ip(
        i_i2c_U_DW_apb_i2c_mstfsm_N421), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_mstfsm_delay_stop_en) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_p_gen_reg ( .ip(n11774), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_debug_p_gen) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_old_is_read_reg ( .ip(n5208), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_old_is_read) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_hs_mcode_en_r_reg ( .ip(i_i2c_hs_mcode_en), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_hs_mcode_en_r) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_hs_mcode_fed_dtctd_r_reg ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N50), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_hs_mcode_fed_dtctd_r)
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N82), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[0])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N83), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[1])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N84), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[2])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt_reg_3_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N85), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[3])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N123), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[0])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N124), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[1])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N125), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[2])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt_reg_3_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N126), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[3])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt_reg_4_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N127), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[4])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt_reg_5_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N128), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[5])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt_reg_6_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N129), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[6])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt_reg_7_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N130), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[7])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_p_det_reg ( .ip(n11775), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_p_det) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_sda_vld_int_reg ( .ip(n5234), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_sda_vld) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_s_det_reg ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_s_det_int), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_s_det) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_s_det_flg_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_s_det_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_s_det_flg_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_s_det_flg_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_s_det_flg_sync_next_sample_syncm1_0_), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_s_det_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_s_det_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_s_det_flg_sync), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_DW_apb_i2c_intctl_s_det_flg_sync_q) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N62), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N63), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N64), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_3_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N65), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_4_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N66), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_5_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N67), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_6_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N68), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_7_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N69), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_8_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N70), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_9_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N71), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_10_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N72), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_11_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N73), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_12_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N74), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_13_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N75), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_14_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N76), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_15_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N77), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt_reg_0_ ( .ip(n5103), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt_reg_1_ ( .ip(n5102), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt_reg_2_ ( .ip(n5101), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt_reg_3_ ( .ip(n5100), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt_reg_4_ ( .ip(n5099), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt_reg_5_ ( .ip(n5098), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt_reg_6_ ( .ip(n5097), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt_reg_7_ ( .ip(n5096), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_scl_edg_hl_q_reg ( .ip(n11769), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_scl_edg_hl_q) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_qq_reg ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_q), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_qq) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count_reg_3_ ( .ip(n5105), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_cmplt_reg ( .ip(n5112), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_tx_cmplt) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_current_state_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_slvfsm_N36), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_slv_debug_cstate[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_slv_cstate_reg_0_ ( .ip(
        i_i2c_slv_debug_cstate[0]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_slv_cstate[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly1_reg ( .ip(n5109), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly1) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ack_vld_reg ( .ip(n5111), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_tx_ack_vld) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_slv_ack_det_reg ( .ip(n5072), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_ack_det) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_rx_done_tog_reg ( .ip(n5071), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_done_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_rx_done_flg_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_rx_done_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_rx_done_flg_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_rx_done_flg_sync_sample_syncl_reg_0_ ( 
        .ip(i_i2c_U_DW_apb_i2c_intctl_U_rx_done_flg_sync_next_sample_syncm1_0_), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_rx_done_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_rx_done_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_rx_done_flg_sync), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_DW_apb_i2c_intctl_rx_done_flg_sync_q) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_tx_flush_reg ( .ip(n5230), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_slv_tx_flush) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_current_state_reg_3_ ( .ip(
        i_i2c_U_DW_apb_i2c_slvfsm_N39), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_slv_debug_cstate[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_slv_cstate_reg_3_ ( .ip(
        i_i2c_slv_debug_cstate[3]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_slv_cstate[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_current_state_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_slvfsm_N38), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_slv_debug_cstate[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_slv_cstate_reg_2_ ( .ip(
        i_i2c_slv_debug_cstate[2]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_slv_cstate[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_data_reg ( .ip(
        i_i2c_U_DW_apb_i2c_toggle_N31), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_data) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_reg_0_ ( .ip(n5084), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_reg_1_ ( .ip(n5083), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_reg_2_ ( .ip(n5082), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_reg_3_ ( .ip(n5081), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_3_) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg_reg_0_ ( .ip(n5080), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg_reg_2_ ( .ip(n5078), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg_reg_4_ ( .ip(n5076), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg_reg_6_ ( .ip(n5074), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg_reg_1_ ( .ip(n5079), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg_reg_3_ ( .ip(n5077), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg_reg_5_ ( .ip(n5075), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg_reg_7_ ( .ip(n5073), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_gen_call_reg ( .ip(n5091), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_gen_call) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_rx_gen_call_r_reg ( .ip(i_i2c_rx_gen_call), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_toggle_rx_gen_call_r) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_rx_gen_call_flg_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_rx_gen_call_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_rx_gen_call_flg_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_rx_gen_call_flg_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_rx_gen_call_flg_sync_next_sample_syncm1_0_), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync_q)
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_hs_mcode_reg ( .ip(n5090), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_hs_mcode) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_rx_hs_mcode_r_reg ( .ip(i_i2c_rx_hs_mcode), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_rx_hs_mcode_r) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_addr_10bit_reg ( .ip(n5093), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_addr_10bit) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_addr_10bit_reg ( .ip(
        i_i2c_rx_addr_10bit), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_debug_addr_10bit) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_slv_read_reg ( .ip(
        i_i2c_U_DW_apb_i2c_rx_shift_rx_slv_read_s), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_rx_slv_read) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_addr_match_reg ( .ip(n5092), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_addr_match) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_current_state_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_slvfsm_N37), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_slv_debug_cstate[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_slv_cstate_reg_1_ ( .ip(
        i_i2c_slv_debug_cstate[1]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_slv_cstate[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_rx_2addr_reg ( .ip(n5231), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_rx_2addr) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rxbyte_rdy_reg ( .ip(n5087), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_rxbyte_rdy) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_addr_reg ( .ip(
        i_i2c_U_DW_apb_i2c_toggle_N32), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_addr) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_activity_reg ( .ip(
        i_i2c_U_DW_apb_i2c_slvfsm_N284), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_activity) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_slave_act_reg ( .ip(i_i2c_slv_activity), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_debug_slave_act) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_slv_activity_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_slv_activity), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_slv_activity_sync_next_sample_syncm1_0_)
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_slv_activity_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_slv_activity_sync_next_sample_syncm1_0_), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_slv_activity_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_en_reg ( .ip(i_i2c_U_DW_apb_i2c_intctl_N4), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_en) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_empty_intr_reg ( .ip(
        i_i2c_ic_intr_stat[4]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_tx_empty_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_slvrd_intx_tog_reg ( .ip(n5118), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_15_ ( 
        .ip(i_i2c_tx_abrt_source[15]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_15_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[15]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_15_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[15]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_rx_aborted_reg ( .ip(n5210), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_rx_aborted) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_slv_rx_aborted_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_slv_rx_aborted), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_slv_rx_aborted_sync_next_sample_syncm1_0_)
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_slv_rx_aborted_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_slv_rx_aborted_sync_next_sample_syncm1_0_), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_slv_rx_aborted_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_push_reg ( .ip(
        i_i2c_U_DW_apb_i2c_rx_shift_N30), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_rx_push) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_push_flg_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_rx_push_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_push_flg_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_push_flg_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_push_flg_sync_next_sample_syncm1_0_), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_rx_push_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_rx_push_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_rx_push_flg_sync), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_DW_apb_i2c_fifo_rx_push_flg_sync_q) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_rx_push_sync_dly_reg ( .ip(i_i2c_rx_push_sync), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_rx_push_sync_dly) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_rx_full_intr_reg ( .ip(
        i_i2c_ic_intr_stat[2]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_rx_full_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_fifo_filled_and_flushed_reg ( .ip(n5086), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_slv_fifo_filled_and_flushed) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_slv_fifo_filled_and_flushed_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_slv_fifo_filled_and_flushed), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_slv_fifo_filled_and_flushed_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_slv_fifo_filled_and_flushed_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_slv_fifo_filled_and_flushed_sync_next_sample_syncm1_0_), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_slv_fifo_filled_and_flushed_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_addressed_reg ( .ip(n5085), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_addressed) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_p_det_intr_reg ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N241), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_p_det_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_p_det_flg_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_p_det_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_p_det_flg_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_p_det_flg_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_p_det_flg_sync_next_sample_syncm1_0_), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_p_det_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_p_det_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_p_det_flg_sync), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_DW_apb_i2c_intctl_p_det_flg_sync_q) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_ack_vld_reg ( .ip(n5089), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_rx_ack_vld) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_ic_enable_sync_vld_reg ( .ip(n5088), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_ic_enable_sync_vld) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count_reg_0_ ( .ip(n5218), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count_reg_1_ ( .ip(n5217), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count_reg_2_ ( .ip(n5216), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count_reg_3_ ( .ip(n5215), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count_reg_4_ ( .ip(n5214), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count_reg_5_ ( .ip(n5213), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count_reg_6_ ( .ip(n5212), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count_reg_7_ ( .ip(n5211), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_scl_hld_low_en_r_reg ( .ip(
        i_i2c_scl_hld_low_en), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_scl_hld_low_en_r) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_tx_abrt_tog_reg ( .ip(n5293), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_flg_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_tx_abrt_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_flg_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_flg_sync_sample_syncl_reg_0_ ( 
        .ip(i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_flg_sync_next_sample_syncm1_0_), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_flg_sync), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_flg_sync_q) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_slvflush_txfifo_tog_reg ( .ip(n5039), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[13])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_13_ ( 
        .ip(i_i2c_tx_abrt_source[13]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_13_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[13]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_13_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[13]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_slv_clr_leftover_tog_reg ( .ip(n5038), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_clr_leftover_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_slv_clr_leftover_flg_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_slv_clr_leftover_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_slv_clr_leftover_flg_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_slv_clr_leftover_flg_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_slv_clr_leftover_flg_sync_next_sample_syncm1_0_), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_slv_clr_leftover_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_slv_clr_leftover_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_slv_clr_leftover_flg_sync), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_slv_clr_leftover_flg_sync_q) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly2_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_N403), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly2) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_N402), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_slv_tx_ready_unconn) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count_reg_0_ ( .ip(n5108), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count_reg_1_ ( .ip(n5107), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count_reg_2_ ( .ip(n5106), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_hs_reg ( .ip(
        i_i2c_U_DW_apb_i2c_toggle_N33), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_hs) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_15_ ( .ip(n5135), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_0_ ( .ip(n5134), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_1_ ( .ip(n5133), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_2_ ( .ip(n5132), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_3_ ( .ip(n5131), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_4_ ( .ip(n5130), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_5_ ( .ip(n5129), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_6_ ( .ip(n5128), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_7_ ( .ip(n5127), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_8_ ( .ip(n5126), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_9_ ( .ip(n5125), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_10_ ( .ip(n5124), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_11_ ( .ip(n5123), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_12_ ( .ip(n5122), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_13_ ( .ip(n5121), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_14_ ( .ip(n5120), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cmplt_reg ( .ip(n5119), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_mstfsm_N382)
         );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_15_ ( .ip(n5067), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_0_ ( .ip(n5066), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_1_ ( .ip(n5065), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_2_ ( .ip(n5064), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_3_ ( .ip(n5063), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_4_ ( .ip(n5062), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_5_ ( .ip(n5061), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_6_ ( .ip(n5060), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_7_ ( .ip(n5059), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_8_ ( .ip(n5058), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_9_ ( .ip(n5057), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_10_ ( .ip(n5056), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_11_ ( .ip(n5055), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_12_ ( .ip(n5054), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_13_ ( .ip(n5053), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_14_ ( .ip(n5052), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_stop_scl_lcnt_en_reg ( .ip(n5048), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_stop_scl_lcnt_en) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_hs_ackdet_tog_reg ( .ip(n5189), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_6_ ( 
        .ip(i_i2c_tx_abrt_source[6]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[6])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_6_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[6]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_6_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[6]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_sbyte_ackdet_tog_reg ( .ip(n5187), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_7_ ( 
        .ip(i_i2c_tx_abrt_source[7]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[7])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_7_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[7]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_7_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[7]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_7b_addr_noack_tog_reg ( .ip(n5194), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_tx_abrt_source[0]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[0])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[0]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[0]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_txdata_noack_tog_reg ( .ip(n5193), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_3_ ( 
        .ip(i_i2c_tx_abrt_source[3]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[3])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_3_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[3]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_3_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[3]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_10addr1_noack_tog_reg ( .ip(n5192), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_1_ ( 
        .ip(i_i2c_tx_abrt_source[1]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[1])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_1_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[1]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[1]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_10addr2_noack_tog_reg ( .ip(n5188), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_2_ ( 
        .ip(i_i2c_tx_abrt_source[2]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[2])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_2_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[2]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[2]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_gcall_noack_tog_reg ( .ip(n5186), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_4_ ( 
        .ip(i_i2c_tx_abrt_source[4]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[4])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_4_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[4]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_4_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[4]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_10b_rd_norstrt_tog_reg ( .ip(n5209), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[10])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_10_ ( 
        .ip(i_i2c_tx_abrt_source[10]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_10_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[10]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_10_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[10]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_slv_arblost_tog_reg ( .ip(n5220), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_14_ ( 
        .ip(i_i2c_tx_abrt_source[14]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_14_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[14]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_14_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[14]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf_reg_0_ ( .ip(n5047), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf_reg_1_ ( .ip(n5046), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf_reg_2_ ( .ip(n5045), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf_reg_3_ ( .ip(n5044), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf_reg_4_ ( .ip(n5043), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf_reg_5_ ( .ip(n5042), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf_reg_6_ ( .ip(n5041), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf_reg_7_ ( .ip(n5040), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_tx_empty_hld_reg ( .ip(n5036), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_tx_empty_hld) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_user_abrt_tog_reg ( .ip(n5205), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[16]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_16_ ( 
        .ip(i_i2c_tx_abrt_source[16]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[16]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_16_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[16]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[16]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_16_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[16]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[16]) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_abrt_in_idle_reg ( .ip(n5204), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_abrt_in_idle) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_scl_lcnt_en_reg ( .ip(n5201), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_scl_lcnt_en) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_bit_count_reg_0_ ( .ip(n5116), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_mst_rx_bit_count[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_bit_count_reg_2_ ( .ip(n5114), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_mst_rx_bit_count[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_bit_count_reg_3_ ( .ip(n5113), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_mst_rx_bit_count[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_current_src_en_reg ( .ip(n5070), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_current_src_en) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_scl_hcnt_en_reg ( .ip(n5202), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_scl_hcnt_en) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_set_tx_empty_en_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_N74), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_set_tx_empty_en) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_set_tx_empty_en_flg_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_set_tx_empty_en_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_set_tx_empty_en_flg_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_set_tx_empty_en_flg_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_set_tx_empty_en_flg_sync_next_sample_syncm1_0_), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_set_tx_empty_en_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_set_tx_empty_en_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_set_tx_empty_en_flg_sync), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_set_tx_empty_en_flg_sync_q) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_current_src_en_reg ( .ip(n5069), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_current_src_en) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_ic_current_src_en_reg ( .ip(
        i_i2c_U_DW_apb_i2c_toggle_N29), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_ic_current_src_en) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en_reg_0_ ( 
        .ip(i_i2c_U_DW_apb_i2c_rx_filter_N207), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[0])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en_reg_1_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[0]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[1])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en_reg_2_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[1]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[2])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en_reg_3_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[2]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[3])
         );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_scl_s_stp_int_reg ( .ip(n5198), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_scl_s_setup_en) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cmplt_reg ( .ip(n5197), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_scl_s_setup_cmplt) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_0_ ( .ip(n5153), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_1_ ( .ip(n5152), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_2_ ( .ip(n5151), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_3_ ( .ip(n5150), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_4_ ( .ip(n5149), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_5_ ( .ip(n5148), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_6_ ( .ip(n5147), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_7_ ( .ip(n5146), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_8_ ( .ip(n5145), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_9_ ( .ip(n5144), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_10_ ( .ip(n5143), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_11_ ( .ip(n5142), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_13_ ( .ip(n5140), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_15_ ( .ip(n5138), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_re_scl_s_hld_en_reg ( .ip(n5196), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_re_scl_s_hld_en) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_gcall_read_tog_reg ( .ip(n4940), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_5_ ( 
        .ip(i_i2c_tx_abrt_source[5]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[5])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_5_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[5]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_5_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[5]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_0_ ( .ip(n5185), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_1_ ( .ip(n5184), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_2_ ( .ip(n5183), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_3_ ( .ip(n5182), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_4_ ( .ip(n5181), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_5_ ( .ip(n5180), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_6_ ( .ip(n5179), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_7_ ( .ip(n5178), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_8_ ( .ip(n5177), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_9_ ( .ip(n5176), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_10_ ( .ip(n5175), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_11_ ( .ip(n5174), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_12_ ( .ip(n5173), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_13_ ( .ip(n5172), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_14_ ( .ip(n5171), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_15_ ( .ip(n5170), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_0_ ( .ip(n5169), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_1_ ( .ip(n5168), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_2_ ( .ip(n5167), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_3_ ( .ip(n5166), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_4_ ( .ip(n5165), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_5_ ( .ip(n5164), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_6_ ( .ip(n5163), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_7_ ( .ip(n5162), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_8_ ( .ip(n5161), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_9_ ( .ip(n5160), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_10_ ( .ip(n5159), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_11_ ( .ip(n5158), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_12_ ( .ip(n5157), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_13_ ( .ip(n5156), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_14_ ( .ip(n5155), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_15_ ( .ip(n5154), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_ic_clk_oe_reg ( .ip(n4958), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ic_clk_oe) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_0_ ( .ip(n4957), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_1_ ( .ip(n4956), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_2_ ( .ip(n4955), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_3_ ( .ip(n4954), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_4_ ( .ip(n4953), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_5_ ( .ip(n4952), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_6_ ( .ip(n4951), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_7_ ( .ip(n4950), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_8_ ( .ip(n4949), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_9_ ( .ip(n4948), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_10_ ( .ip(n4947), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_11_ ( .ip(n4946), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_12_ ( .ip(n4945), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_start_sda_gate_r_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_N272), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_tx_shift_start_sda_gate_r) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_mst_slv_ack_ext_r_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_mst_slv_ack_ext), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_tx_shift_mst_slv_ack_ext_r) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_gen_call_reg ( .ip(n4660), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_gen_call_intr_reg ( .ip(
        i_i2c_ic_intr_stat[11]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_gen_call_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_activity_reg ( .ip(n4657), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_activity_intr_reg ( .ip(
        i_i2c_ic_intr_stat[8]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_activity_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_stop_det_reg ( .ip(n4659), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_stop_det_intr_reg ( .ip(
        i_i2c_ic_intr_stat[9]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_stop_det_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_start_det_reg ( .ip(n4658), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_start_det_intr_reg ( .ip(
        i_i2c_ic_intr_stat[10]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_start_det_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_rx_done_reg ( .ip(n4656), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_rx_done_intr_reg ( .ip(
        i_i2c_ic_intr_stat[7]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_rx_done_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_16_ ( .ip(n5219), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[16]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_0_ ( .ip(n4707), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_1_ ( .ip(n4706), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_2_ ( .ip(n4705), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_3_ ( .ip(n4704), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_4_ ( .ip(n4703), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_5_ ( .ip(n4702), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_6_ ( .ip(n4701), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_7_ ( .ip(n4700), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_8_ ( .ip(n4699), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_10_ ( .ip(n4697), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_11_ ( .ip(n4696), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_12_ ( .ip(n4695), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_13_ ( .ip(n4694), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_14_ ( .ip(n4693), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_15_ ( .ip(n4692), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_tx_abrt_reg ( .ip(n4655), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_intr_reg ( .ip(
        i_i2c_ic_intr_stat[6]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_tx_abrt_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_rd_req_reg ( .ip(n4654), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_rd_req_intr_reg ( .ip(
        i_i2c_ic_intr_stat[5]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_rd_req_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_rx_under_reg ( .ip(n4653), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_rx_under_intr_reg ( .ip(
        i_i2c_ic_intr_stat[0]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_rx_under_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_rx_over_reg ( .ip(n4652), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_rx_over_intr_reg ( .ip(
        i_i2c_ic_intr_stat[1]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_rx_over_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_tx_over_reg ( .ip(n4651), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_over_intr_reg ( .ip(
        i_i2c_ic_intr_stat[3]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_tx_over_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_0_ ( .ip(n4661), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_1_ ( .ip(n4662), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_2_ ( .ip(n4663), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_3_ ( .ip(n4664), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_4_ ( .ip(n4665), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_5_ ( .ip(n4666), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_6_ ( .ip(n4667), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_7_ ( .ip(n4668), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_8_ ( .ip(n4669), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_9_ ( .ip(n4670), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_10_ ( .ip(n4671), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_11_ ( .ip(n4672), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_12_ ( .ip(n4673), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_13_ ( .ip(n4674), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_14_ ( .ip(n4675), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_15_ ( .ip(n4676), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_16_ ( .ip(n4677), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[16]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_17_ ( .ip(n4678), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[17]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_18_ ( .ip(n4679), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[18]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_19_ ( .ip(n4680), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[19]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_20_ ( .ip(n4681), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[20]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_21_ ( .ip(n4682), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[21]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_22_ ( .ip(n4683), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[22]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_23_ ( .ip(n4684), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[23]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_24_ ( .ip(n4685), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[24]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_25_ ( .ip(n4686), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[25]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_26_ ( .ip(n4687), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[26]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_28_ ( .ip(n4689), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[28]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_29_ ( .ip(n4690), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[29]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_30_ ( .ip(n4691), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[30]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg_reg_0_ ( .ip(n4936), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[0]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_7__0_ ( .ip(n4928), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[0]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_6__0_ ( .ip(n4927), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[8]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_5__0_ ( .ip(n4926), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[16]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_4__0_ ( .ip(n4925), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[24]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_3__0_ ( .ip(n4924), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[32]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_2__0_ ( .ip(n4923), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[40]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_1__0_ ( .ip(n4922), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[48]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_0__0_ ( .ip(n4921), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[56]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg_reg_1_ ( .ip(n4935), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[1]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_7__1_ ( .ip(n4920), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[1]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_6__1_ ( .ip(n4919), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[9]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_5__1_ ( .ip(n4918), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[17]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_4__1_ ( .ip(n4917), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[25]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_3__1_ ( .ip(n4916), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[33]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_2__1_ ( .ip(n4915), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[41]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_1__1_ ( .ip(n4914), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[49]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_0__1_ ( .ip(n4913), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[57]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg_reg_2_ ( .ip(n4934), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[2]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_7__2_ ( .ip(n4912), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[2]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_6__2_ ( .ip(n4911), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[10]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_5__2_ ( .ip(n4910), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[18]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_4__2_ ( .ip(n4909), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[26]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_3__2_ ( .ip(n4908), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[34]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_2__2_ ( .ip(n4907), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[42]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_1__2_ ( .ip(n4906), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[50]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_0__2_ ( .ip(n4905), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[58]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg_reg_3_ ( .ip(n4933), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[3]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_7__3_ ( .ip(n4904), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[3]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_6__3_ ( .ip(n4903), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[11]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_5__3_ ( .ip(n4902), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[19]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_4__3_ ( .ip(n4901), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[27]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_3__3_ ( .ip(n4900), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[35]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_2__3_ ( .ip(n4899), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[43]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_1__3_ ( .ip(n4898), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[51]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_0__3_ ( .ip(n4897), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[59]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg_reg_4_ ( .ip(n4932), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[4]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_7__4_ ( .ip(n4896), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[4]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_6__4_ ( .ip(n4895), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[12]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_5__4_ ( .ip(n4894), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[20]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_4__4_ ( .ip(n4893), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[28]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_3__4_ ( .ip(n4892), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[36]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_2__4_ ( .ip(n4891), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[44]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_1__4_ ( .ip(n4890), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[52]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_0__4_ ( .ip(n4889), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[60]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg_reg_5_ ( .ip(n4931), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[5]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_7__5_ ( .ip(n4888), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[5]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_6__5_ ( .ip(n4887), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[13]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_5__5_ ( .ip(n4886), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[21]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_4__5_ ( .ip(n4885), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[29]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_3__5_ ( .ip(n4884), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[37]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_2__5_ ( .ip(n4883), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[45]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_1__5_ ( .ip(n4882), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[53]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_0__5_ ( .ip(n4881), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[61]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg_reg_6_ ( .ip(n4930), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[6]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_7__6_ ( .ip(n4880), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[6]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_6__6_ ( .ip(n4879), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[14]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_5__6_ ( .ip(n4878), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[22]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_4__6_ ( .ip(n4877), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[30]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_3__6_ ( .ip(n4876), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[38]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_2__6_ ( .ip(n4875), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[46]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_1__6_ ( .ip(n4874), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[54]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_0__6_ ( .ip(n4873), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[62]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg_reg_7_ ( .ip(n4929), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[7]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_7__7_ ( .ip(n4872), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[7]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_6__7_ ( .ip(n4871), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[15]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_5__7_ ( .ip(n4870), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[23]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_4__7_ ( .ip(n4869), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[31]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_3__7_ ( .ip(n4868), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[39]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_2__7_ ( .ip(n4867), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[47]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_1__7_ ( .ip(n4866), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[55]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_0__7_ ( .ip(n4865), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[63]) );
  drp_1 i_apb_U_DW_apb_ahbsif_psel_en_reg ( .ip(n4212), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_psel_en) );
  drp_1 i_apb_U_DW_apb_ahbsif_penable_reg ( .ip(n4211), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_penable) );
  drp_1 i_ssi_U_mstfsm_bit_cnt_reg_0_ ( .ip(n4210), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_bit_cnt[0]) );
  drp_1 i_ssi_U_mstfsm_bit_cnt_reg_1_ ( .ip(n4209), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_bit_cnt[1]) );
  drp_1 i_ssi_U_mstfsm_bit_cnt_reg_2_ ( .ip(n4208), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_bit_cnt[2]) );
  drp_1 i_ssi_U_mstfsm_bit_cnt_reg_3_ ( .ip(n4207), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_bit_cnt[3]) );
  drp_1 i_ssi_U_mstfsm_bit_cnt_reg_4_ ( .ip(n4206), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_bit_cnt[4]) );
  drp_1 i_ssi_U_mstfsm_ctrl_cnt_reg_0_ ( .ip(n4205), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_ctrl_cnt[0]) );
  drp_1 i_ssi_U_mstfsm_ctrl_cnt_reg_1_ ( .ip(n4204), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_ctrl_cnt[1]) );
  drp_1 i_ssi_U_mstfsm_ctrl_cnt_reg_2_ ( .ip(n4203), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_ctrl_cnt[2]) );
  drp_1 i_ssi_U_mstfsm_ctrl_cnt_reg_3_ ( .ip(n4202), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_ctrl_cnt[3]) );
  drp_1 i_ssi_U_mstfsm_spi1_control_reg ( .ip(n4201), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_spi1_control) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_14_ ( .ip(n4198), .ck(i_ssi_ssi_clk), 
        .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[14]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_13_ ( .ip(n4197), .ck(i_ssi_ssi_clk), 
        .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[13]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_11_ ( .ip(n4195), .ck(i_ssi_ssi_clk), 
        .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[11]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_9_ ( .ip(n4193), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[9]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_8_ ( .ip(n4192), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[8]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_7_ ( .ip(n4191), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[7]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_6_ ( .ip(n4190), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[6]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_5_ ( .ip(n4189), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[5]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_4_ ( .ip(n4188), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[4]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_3_ ( .ip(n4187), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[3]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_2_ ( .ip(n4186), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[2]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_0_ ( .ip(n4184), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[0]) );
  drp_1 i_ssi_U_mstfsm_spi0_control_reg ( .ip(n4183), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_spi0_control) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_arb_lost_tog_reg ( .ip(n4182), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_chk_win_reg ( .ip(n4181), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_chk_win) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_tx_pop_tog_reg ( .ip(n4180), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_pop_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_mst_tx_ack_int_reg ( .ip(n4179), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_mst_tx_ack_vld) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_s_det_tog_reg ( .ip(n4178), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_s_det_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_q_reg ( .ip(n4177), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_q) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr_reg_0_ ( .ip(n4176), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr_reg_1_ ( .ip(n4175), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr_reg_2_ ( .ip(n4174), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr_reg_3_ ( .ip(n4173), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_rx_gen_call_tog_reg ( .ip(n4172), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_gen_call_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_slv_arb_lost_reg ( .ip(n4171), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_slv_arb_lost) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_rx_push_tog_reg ( .ip(n4170), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_push_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_p_det_tog_reg ( .ip(n4169), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_p_det_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ack_det_reg ( .ip(n4168), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ack_det) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_bwen_reg ( .ip(n4167), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_mst_rx_bwen) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_hcnt_cmplt_int_reg ( .ip(n4166), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_hcnt_cmplt_int) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_0_ ( .ip(n4165), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_1_ ( .ip(n4164), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_2_ ( .ip(n4163), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_3_ ( .ip(n4162), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_4_ ( .ip(n4161), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_5_ ( .ip(n4160), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_7_ ( .ip(n4158), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_8_ ( .ip(n4157), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_9_ ( .ip(n4156), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_10_ ( .ip(n4155), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_11_ ( .ip(n4154), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_13_ ( .ip(n4152), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_scl_hcnt_en_int_reg ( .ip(n4149), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_scl_hcnt_en) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_data_scl_lcnt_en_reg ( .ip(n4148), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_data_scl_lcnt_en) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count_reg_0_ ( .ip(n4147), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count_reg_1_ ( .ip(n4146), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count_reg_2_ ( .ip(n4145), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count_reg_3_ ( .ip(n4144), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_set_tx_empty_en_tog_reg ( .ip(n4143), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_set_tx_empty_en_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr_reg_0_ ( .ip(n4142), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr_reg_1_ ( .ip(n4141), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr_reg_2_ ( .ip(n4140), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr_reg_3_ ( .ip(n4139), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr_reg_4_ ( .ip(n4138), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr_reg_5_ ( .ip(n4137), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr_reg_6_ ( .ip(n4136), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr_reg_7_ ( .ip(n4135), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_mst_tx_bwen_reg ( .ip(n4134), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_mst_tx_bwen) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_push_data_reg_0_ ( .ip(n4133), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_push_data[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_push_data_reg_1_ ( .ip(n4132), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_push_data[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_push_data_reg_2_ ( .ip(n4131), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_push_data[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_push_data_reg_3_ ( .ip(n4130), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_push_data[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_push_data_reg_4_ ( .ip(n4129), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_push_data[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_push_data_reg_5_ ( .ip(n4128), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_push_data[5]) );
  drp_2 i_ssi_U_sclkgen_ssi_cnt_reg_13_ ( .ip(i_ssi_U_sclkgen_N53), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[13])
         );
  drp_2 i_ssi_U_shift_U_tx_shifter_txd_reg ( .ip(n4395), .ck(i_ssi_ssi_clk), 
        .rb(i_ssi_ssi_rst_n), .q(i_ssi_txd) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_push_data_reg_6_ ( .ip(n4127), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_push_data[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_push_data_reg_7_ ( .ip(n4126), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_push_data[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[1]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_15_ ( .ip(n4942), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[15]) );
  drp_2 i_ssi_U_regfile_ctrlr1_reg_7_ ( .ip(n4603), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[7]) );
  drsp_1 i_apb_U_DW_apb_ahbsif_hready_resp_reg ( .ip(n4824), .ck(HCLK_hclk), 
        .rb(1'b1), .s(n11759), .q(i_apb_hready_resp) );
  drsp_1 i_ssi_U_regfile_imr_ir_reg_3_ ( .ip(n4647), .ck(PCLK_pclk), .rb(1'b1), 
        .s(n11766), .q(i_ssi_imr[3]) );
  drsp_1 i_ssi_U_regfile_imr_ir_reg_4_ ( .ip(n4646), .ck(PCLK_pclk), .rb(1'b1), 
        .s(n11766), .q(i_ssi_imr[4]) );
  drsp_1 i_ssi_U_regfile_imr_ir_reg_1_ ( .ip(n4649), .ck(PCLK_pclk), .rb(1'b1), 
        .s(n11766), .q(i_ssi_imr[1]) );
  drsp_1 i_ssi_U_regfile_imr_ir_reg_2_ ( .ip(n4648), .ck(PCLK_pclk), .rb(1'b1), 
        .s(n11766), .q(i_ssi_imr[2]) );
  drsp_1 i_ssi_U_regfile_imr_ir_reg_0_ ( .ip(n4650), .ck(PCLK_pclk), .rb(1'b1), 
        .s(n11766), .q(i_ssi_imr[0]) );
  drsp_1 i_ssi_U_regfile_imr_ir_reg_5_ ( .ip(n4645), .ck(PCLK_pclk), .rb(1'b1), 
        .s(n11766), .q(i_ssi_imr[5]) );
  drsp_1 i_ssi_U_regfile_ctrlr0_ir_reg_7_ ( .ip(n4594), .ck(PCLK_pclk), .rb(
        1'b1), .s(n11766), .q(i_ssi_U_regfile_ctrlr0_ir_int_7) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_rd_addr_int_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N44), .ck(PCLK_pclk), .q(
        i_i2c_tx_rd_addr[0]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_rd_addr_int_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N46), .ck(PCLK_pclk), .q(
        i_i2c_tx_rd_addr[2]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_rd_addr_int_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N45), .ck(PCLK_pclk), .q(
        i_i2c_tx_rd_addr[1]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_rd_addr_at_max_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N39), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_rd_addr_at_max) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_error_int_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N38), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_error_ir) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_wr_addr_int_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N41), .ck(PCLK_pclk), .q(
        i_i2c_tx_wr_addr[0]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_full_int_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N37), .ck(PCLK_pclk), .q(
        i_i2c_rx_full) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_word_count_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N47), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[0]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_rd_addr_int_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N45), .ck(PCLK_pclk), .q(
        i_i2c_rx_rd_addr[1]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_wr_addr_at_max_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N40), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_wr_addr_at_max) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_rd_addr_int_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N46), .ck(PCLK_pclk), .q(
        i_i2c_rx_rd_addr[2]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_wr_addr_int_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N42), .ck(PCLK_pclk), .q(
        i_i2c_rx_wr_addr[1]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_error_int_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N38), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_rx_error_ir) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_wr_addr_int_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N41), .ck(PCLK_pclk), .q(
        i_i2c_rx_wr_addr[0]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_rd_addr_int_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N44), .ck(PCLK_pclk), .q(
        i_i2c_rx_rd_addr[0]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_full_int_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N37), .ck(PCLK_pclk), .q(
        i_i2c_tx_full) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_wr_addr_int_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N42), .ck(PCLK_pclk), .q(
        i_i2c_tx_wr_addr[1]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_wr_addr_int_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N43), .ck(PCLK_pclk), .q(
        i_i2c_rx_wr_addr[2]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_word_count_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N48), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[1]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_wr_addr_at_max_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N40), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_wr_addr_at_max) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_rd_addr_at_max_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N39), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_rd_addr_at_max) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_word_count_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N47), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[0]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_word_count_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N48), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[1]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_wr_addr_int_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N43), .ck(PCLK_pclk), .q(
        i_i2c_tx_wr_addr[2]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_word_count_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N49), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[2]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_empty_n_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N33), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_empty_n) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_almost_empty_n_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N34), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_almost_empty_n) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_word_count_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N49), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[2]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_empty_n_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N33), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_empty_n) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_rd_addr_int_reg_1_ ( .ip(
        i_ssi_U_fifo_U_rx_fifo_N45), .ck(PCLK_pclk), .q(i_ssi_rx_rd_addr[1])
         );
  dp_1 i_ssi_U_fifo_U_rx_fifo_rd_addr_int_reg_2_ ( .ip(
        i_ssi_U_fifo_U_rx_fifo_N46), .ck(PCLK_pclk), .q(i_ssi_rx_rd_addr[2])
         );
  dp_1 i_ssi_U_fifo_U_rx_fifo_rd_addr_int_reg_0_ ( .ip(n11768), .ck(PCLK_pclk), 
        .q(i_ssi_rx_rd_addr[0]) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_rd_addr_at_max_reg ( .ip(
        i_ssi_U_fifo_U_rx_fifo_N39), .ck(PCLK_pclk), .q(
        i_ssi_U_fifo_U_rx_fifo_rd_addr_at_max) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_almost_full_int_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N36), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_i_rx_almost_full) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_error_int_reg ( .ip(i_ssi_U_fifo_U_tx_fifo_N38), 
        .ck(PCLK_pclk), .q(i_ssi_U_fifo_tx_error_ir) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_error_int_reg ( .ip(i_ssi_U_fifo_U_rx_fifo_N38), 
        .ck(PCLK_pclk), .q(i_ssi_U_fifo_rx_error_ir) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_rd_addr_int_reg_1_ ( .ip(
        i_ssi_U_fifo_U_tx_fifo_N45), .ck(PCLK_pclk), .q(i_ssi_tx_rd_addr[1])
         );
  dp_1 i_ssi_U_fifo_U_tx_fifo_rd_addr_int_reg_0_ ( .ip(n11767), .ck(PCLK_pclk), 
        .q(i_ssi_tx_rd_addr[0]) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_full_int_reg ( .ip(i_ssi_U_fifo_U_tx_fifo_N37), 
        .ck(PCLK_pclk), .q(i_ssi_tx_full) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_full_int_reg ( .ip(n11777), .ck(PCLK_pclk), .q(
        i_ssi_rx_full) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_wr_addr_int_reg_0_ ( .ip(
        i_ssi_U_fifo_U_tx_fifo_N41), .ck(PCLK_pclk), .q(i_ssi_tx_wr_addr[0])
         );
  dp_1 i_ssi_U_fifo_U_tx_fifo_rd_addr_at_max_reg ( .ip(
        i_ssi_U_fifo_U_tx_fifo_N39), .ck(PCLK_pclk), .q(
        i_ssi_U_fifo_U_tx_fifo_rd_addr_at_max) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_word_count_reg_0_ ( .ip(
        i_ssi_U_fifo_U_tx_fifo_N47), .ck(PCLK_pclk), .q(
        i_ssi_U_fifo_unconnected_tx_wrd_count[0]) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_wr_addr_int_reg_1_ ( .ip(
        i_ssi_U_fifo_U_tx_fifo_N42), .ck(PCLK_pclk), .q(i_ssi_tx_wr_addr[1])
         );
  dp_1 i_ssi_U_fifo_U_rx_fifo_word_count_reg_0_ ( .ip(
        i_ssi_U_fifo_U_rx_fifo_N47), .ck(PCLK_pclk), .q(
        i_ssi_U_fifo_unconnected_rx_wrd_count[0]) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_wr_addr_at_max_reg ( .ip(
        i_ssi_U_fifo_U_rx_fifo_N40), .ck(PCLK_pclk), .q(
        i_ssi_U_fifo_U_rx_fifo_wr_addr_at_max) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_wr_addr_at_max_reg ( .ip(
        i_ssi_U_fifo_U_tx_fifo_N40), .ck(PCLK_pclk), .q(
        i_ssi_U_fifo_U_tx_fifo_wr_addr_at_max) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_wr_addr_int_reg_2_ ( .ip(
        i_ssi_U_fifo_U_tx_fifo_N43), .ck(PCLK_pclk), .q(i_ssi_tx_wr_addr[2])
         );
  dp_1 i_ssi_U_fifo_U_tx_fifo_word_count_reg_2_ ( .ip(n11779), .ck(PCLK_pclk), 
        .q(i_ssi_U_fifo_unconnected_tx_wrd_count[2]) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_word_count_reg_1_ ( .ip(
        i_ssi_U_fifo_U_tx_fifo_N48), .ck(PCLK_pclk), .q(
        i_ssi_U_fifo_unconnected_tx_wrd_count[1]) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_word_count_reg_1_ ( .ip(
        i_ssi_U_fifo_U_rx_fifo_N48), .ck(PCLK_pclk), .q(
        i_ssi_U_fifo_unconnected_rx_wrd_count[1]) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_word_count_reg_2_ ( .ip(
        i_ssi_U_fifo_U_rx_fifo_N49), .ck(PCLK_pclk), .q(
        i_ssi_U_fifo_unconnected_rx_wrd_count[2]) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_empty_n_reg ( .ip(i_ssi_U_fifo_U_tx_fifo_N33), 
        .ck(PCLK_pclk), .q(i_ssi_U_fifo_U_tx_fifo_empty_n) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_almost_full_int_reg ( .ip(
        i_ssi_U_fifo_U_rx_fifo_N36), .ck(PCLK_pclk), .q(
        i_ssi_U_fifo_switch_almost_full) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_almost_empty_n_reg ( .ip(
        i_ssi_U_fifo_U_tx_fifo_N34), .ck(PCLK_pclk), .q(
        i_ssi_U_fifo_U_tx_fifo_almost_empty_n) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_empty_n_reg ( .ip(i_ssi_U_fifo_U_rx_fifo_N33), 
        .ck(PCLK_pclk), .q(i_ssi_U_fifo_U_rx_fifo_empty_n) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_rd_addr_int_reg_2_ ( .ip(
        i_ssi_U_fifo_U_tx_fifo_N46), .ck(PCLK_pclk), .q(i_ssi_tx_rd_addr[2])
         );
  drp_2 i_ssi_U_regfile_baudr_reg_4_ ( .ip(n4630), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[4]) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda_r_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda), .ck(i_i2c_ic_clk), .rb(1'b1), .s(n11747), .q(i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda_r) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_start_sda_reg ( .ip(n11771), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11747), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_start_sda) );
  drsp_1 i_i2c_U_DW_apb_i2c_clk_gen_count_en_reg ( .ip(n4125), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11747), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_count_en) );
  drsp_1 i_i2c_U_DW_apb_i2c_sync_tx_empty_sync_r_reg ( .ip(n5245), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11747), .q(
        i_i2c_U_DW_apb_i2c_sync_tx_empty_sync_r) );
  drsp_1 i_i2c_U_DW_apb_i2c_rx_filter_scl_int_q_reg ( .ip(n11776), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11726), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_scl_int_q) );
  drsp_1 i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt_reg_0_ ( .ip(n5094), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11726), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt[0]) );
  drsp_1 i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt_reg_1_ ( .ip(n5095), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11726), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt[1]) );
  drsp_1 i_i2c_U_DW_apb_i2c_rx_filter_scl_clk_int_reg ( .ip(n5137), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11747), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_scl_clk_int) );
  drsp_1 i_i2c_U_DW_apb_i2c_rx_filter_sda_data_int_reg ( .ip(n5136), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11726), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_sda_data_int) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_stop_scl_reg ( .ip(n5050), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11747), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_stop_scl) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_stop_sda_reg ( .ip(n5049), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11726), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_stop_sda) );
  drsp_1 i_i2c_U_DW_apb_i2c_rx_filter_sda_int_q_reg ( .ip(i_i2c_sda_int), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11726), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_sda_int_q) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl_reg ( .ip(n4961), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11747), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda_reg ( .ip(n4960), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11747), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_data_scl_reg ( .ip(n4124), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11747), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_data_scl) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_data_sda_reg ( .ip(n5110), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11747), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_data_sda) );
  drsp_1 i_i2c_U_DW_apb_i2c_rx_filter_sda_post_hold_done_reg ( .ip(n5104), 
        .ck(i_i2c_ic_clk), .rb(1'b1), .s(n11726), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_sda_post_hold_done) );
  drsp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_data_scl_reg ( .ip(n4937), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11726), .q(i_i2c_mst_rx_data_scl) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_data_sda_reg ( .ip(n4123), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11726), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_data_sda) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_stop_sda_gate_r_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_N281), .ck(i_i2c_ic_clk), .rb(1'b1), .s(
        n11747), .q(i_i2c_U_DW_apb_i2c_tx_shift_stop_sda_gate_r) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_data_sda_prev_r_reg ( .ip(n4941), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11726), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_data_sda_prev_r) );
  drp_2 i_ssi_U_sclkgen_ssi_cnt_reg_1_ ( .ip(i_ssi_U_sclkgen_N41), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[1])
         );
  drp_1 i_ssi_U_sclkgen_sclk_re_ir_reg ( .ip(i_ssi_U_sclkgen_N74), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_sclk_re) );
  drp_1 i_ssi_U_shift_rx_push_tgl_reg ( .ip(n4451), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_rx_push) );
  drp_2 i_ssi_U_regfile_ctrlr1_reg_11_ ( .ip(n4615), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[11]) );
  drsp_1 i_ssi_U_regfile_ctrlr0_ir_reg_1_ ( .ip(n4589), .ck(PCLK_pclk), .rb(
        1'b1), .s(n11766), .q(i_ssi_dfs[1]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_15_ ( .ip(n4611), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[15]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_1_ ( .ip(n4609), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[1]) );
  drp_1 i_ssi_U_regfile_mwcr_ir_reg_0_ ( .ip(n4637), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_mwcr[0]) );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_0_ ( .ip(n11781), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[0]) );
  drp_1 i_ssi_U_regfile_mwcr_ir_reg_1_ ( .ip(n4636), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_mwcr[1]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_3_ ( .ip(n4591), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_dfs[3]) );
  drp_1 i_apb_U_DW_apb_ahbsif_state_reg_0_ ( .ip(n5311), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_state[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_14_ ( .ip(n4943), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[14]) );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_14_ ( .ip(i_ssi_U_sclkgen_N54), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[14])
         );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_2_ ( .ip(i_ssi_U_sclkgen_N42), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[2])
         );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_11_ ( .ip(i_ssi_U_sclkgen_N51), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[11])
         );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_13_ ( .ip(n4944), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_12_ ( .ip(n5141), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_14_ ( .ip(n5139), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[14]) );
  drp_1 i_ssi_U_regfile_baudr_reg_14_ ( .ip(n4620), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[14]) );
  drp_1 i_ssi_U_regfile_baudr_reg_5_ ( .ip(n4629), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[5]) );
  drp_1 i_ssi_U_regfile_baudr_reg_6_ ( .ip(n4628), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_int_d_reg ( .ip(n11776), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_int_d) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_tx_abrt_r_reg ( .ip(
        i_i2c_U_DW_apb_i2c_toggle_tx_abrt), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_toggle_tx_abrt_r) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt_reg_7_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N89), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[7])
         );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_15_ ( .ip(n4150), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_6_ ( .ip(n4159), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[6]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_14_ ( .ip(n4601), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_cfs[2]) );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_4_ ( .ip(i_ssi_U_sclkgen_N44), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[4])
         );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_8_ ( .ip(i_ssi_U_sclkgen_N48), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[8])
         );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_9_ ( .ip(i_ssi_U_sclkgen_N49), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[9])
         );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_5_ ( .ip(i_ssi_U_sclkgen_N45), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[5])
         );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_10_ ( .ip(i_ssi_U_sclkgen_N50), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[10])
         );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_12_ ( .ip(i_ssi_U_sclkgen_N52), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[12])
         );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_3_ ( .ip(i_ssi_U_sclkgen_N43), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[3])
         );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_6_ ( .ip(i_ssi_U_sclkgen_N46), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[6])
         );
  drp_1 i_ssi_U_regfile_baudr_reg_2_ ( .ip(n4632), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[2]) );
  drp_1 i_ssi_U_mstfsm_fsm_multi_mst_reg ( .ip(n11761), .ck(i_ssi_ssi_clk), 
        .rb(i_ssi_ssi_rst_n), .q(i_ssi_fsm_multi_mst) );
  drp_1 i_ssi_U_regfile_baudr_reg_1_ ( .ip(n4633), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[1]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_12_ ( .ip(n4614), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[12]) );
  drsp_1 i_ssi_U_regfile_baudr_reg_12_ ( .ip(n4622), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .s(1'b0), .q(i_ssi_baudr[12]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_3_ ( .ip(n4407), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[3]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_6_ ( .ip(n4404), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[6]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_7_ ( .ip(n4403), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[7]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_4_ ( .ip(n4406), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[4]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_11_ ( .ip(n4399), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[11]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_13_ ( .ip(n4397), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[13]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_10_ ( .ip(n4400), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[10]) );
  drp_1 i_ssi_U_mstfsm_ssi_oe_n_reg ( .ip(n5677), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(n11748) );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_7_ ( .ip(i_ssi_U_sclkgen_N47), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[7])
         );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_2_ ( .ip(n4408), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[2]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_0_ ( .ip(n4410), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[0]) );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_15_ ( .ip(i_ssi_U_sclkgen_N55), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[15])
         );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_10_ ( .ip(n4194), .ck(i_ssi_ssi_clk), 
        .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[10]) );
  drp_1 i_ssi_U_mstfsm_c_state_reg_2_ ( .ip(i_ssi_U_mstfsm_N222), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_c_state[2]) );
  drp_1 i_ssi_U_mstfsm_c_state_reg_0_ ( .ip(i_ssi_U_mstfsm_N220), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_c_state[0]) );
  drp_1 i_ssi_U_mstfsm_fsm_sleep_reg ( .ip(n5233), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_fsm_sleep) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_15_ ( .ip(n4396), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[15]) );
  drp_1 i_ssi_U_shift_ss_n_reg_0_ ( .ip(n5679), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(n11724) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_16_ ( .ip(n4200), .ck(i_ssi_ssi_clk), 
        .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[16]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_12_ ( .ip(n4398), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[12]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_12_ ( .ip(n4196), .ck(i_ssi_ssi_clk), 
        .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[12]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_14_ ( .ip(n4411), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[14]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_1_ ( .ip(n4185), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_14_ ( .ip(n4151), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_12_ ( .ip(n4153), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[12]) );
  drp_1 i_ssi_U_regfile_baudr_reg_3_ ( .ip(n4631), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[3]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_14_ ( .ip(n4612), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[14]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_10_ ( .ip(n4616), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[10]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_9_ ( .ip(n4401), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[9]) );
  drp_2 i_i2c_U_DW_apb_i2c_sync_U_ic_hs_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_hs_sync_next_sample_syncm1_0_), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt_reg_5_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N87), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[5])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt_reg_6_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N88), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[6])
         );
  drp_1 i_ssi_U_shift_tx_pop_tgl_reg ( .ip(n4585), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_tx_pop) );
  drp_2 i_ssi_U_regfile_ctrlr1_reg_13_ ( .ip(n4613), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[13]) );
  drsp_2 i_ssi_U_regfile_ctrlr0_ir_reg_0_ ( .ip(n4588), .ck(PCLK_pclk), .rb(
        1'b1), .s(n11766), .q(i_ssi_dfs[0]) );
  drsp_2 i_ssi_U_regfile_ctrlr0_ir_reg_2_ ( .ip(n4590), .ck(PCLK_pclk), .rb(
        1'b1), .s(n11766), .q(i_ssi_dfs[2]) );
  drp_2 i_ssi_U_mstfsm_frame_cnt_reg_15_ ( .ip(n4199), .ck(i_ssi_ssi_clk), 
        .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[15]) );
  drp_1 i_ssi_U_regfile_baudr_reg_10_ ( .ip(n4624), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r_reg ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_hs), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt_reg_4_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N86), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[4])
         );
  drp_1 i_ssi_U_regfile_baud2_reg ( .ip(n5241), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baud2) );
  drp_1 i_ssi_U_regfile_start_xfer_reg ( .ip(i_ssi_U_regfile_N452), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_ssi_start_xfer) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_wr_addr_int_reg_1_ ( .ip(
        i_ssi_U_fifo_U_rx_fifo_N42), .ck(PCLK_pclk), .q(i_ssi_rx_wr_addr[1])
         );
  dp_1 i_ssi_U_fifo_U_rx_fifo_wr_addr_int_reg_0_ ( .ip(
        i_ssi_U_fifo_U_rx_fifo_N41), .ck(PCLK_pclk), .q(i_ssi_rx_wr_addr[0])
         );
  dp_1 i_ssi_U_fifo_U_rx_fifo_wr_addr_int_reg_2_ ( .ip(
        i_ssi_U_fifo_U_rx_fifo_N43), .ck(PCLK_pclk), .q(i_ssi_rx_wr_addr[2])
         );
  inv_1 U5566 ( .ip(n5322), .op(n9371) );
  inv_1 U5567 ( .ip(n5324), .op(n9370) );
  nand4_1 U5568 ( .ip1(n9666), .ip2(n9438), .ip3(n9437), .ip4(n9436), .op(
        n9439) );
  nand4_1 U5569 ( .ip1(n9666), .ip2(n9442), .ip3(n9441), .ip4(n9440), .op(
        n9443) );
  buf_2 U5570 ( .ip(n10116), .op(n5269) );
  nor3_2 U5571 ( .ip1(n11471), .ip2(n11470), .ip3(n11473), .op(n11507) );
  nand2_2 U5572 ( .ip1(n10041), .ip2(n10040), .op(n11461) );
  buf_2 U5573 ( .ip(n10042), .op(n5270) );
  inv_2 U5574 ( .ip(n10026), .op(n6596) );
  nor2_2 U5575 ( .ip1(n5377), .ip2(n5404), .op(n5380) );
  inv_2 U5576 ( .ip(n10371), .op(n5258) );
  nor2_2 U5577 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(n6551), .op(n9360) );
  inv_2 U5578 ( .ip(n8125), .op(n5273) );
  inv_2 U5579 ( .ip(n6720), .op(n6721) );
  nand2_4 U5580 ( .ip1(n5302), .ip2(n5535), .op(n10232) );
  nand2_2 U5581 ( .ip1(n5303), .ip2(n5534), .op(n5302) );
  xor2_2 U5582 ( .ip1(i_ssi_U_mstfsm_bit_cnt[1]), .ip2(i_ssi_dfs[1]), .op(
        n5663) );
  nand2_2 U5583 ( .ip1(n5613), .ip2(n5619), .op(n5803) );
  nand2_1 U5584 ( .ip1(n5795), .ip2(n5340), .op(n5404) );
  and3_2 U5585 ( .ip1(n5586), .ip2(n5585), .ip3(n5584), .op(n5587) );
  nand2_1 U5586 ( .ip1(n5674), .ip2(n5438), .op(n5328) );
  nor2_2 U5587 ( .ip1(n5805), .ip2(n9960), .op(n5794) );
  nand2_2 U5588 ( .ip1(n5327), .ip2(n5587), .op(n5329) );
  inv_2 U5589 ( .ip(n5761), .op(n5590) );
  nand2_2 U5590 ( .ip1(n5804), .ip2(n5589), .op(n5761) );
  nor2_2 U5591 ( .ip1(n5335), .ip2(n10350), .op(n6182) );
  nand3_4 U5592 ( .ip1(n6117), .ip2(n6116), .ip3(n6115), .op(n10350) );
  nand2_2 U5593 ( .ip1(n5796), .ip2(n5741), .op(n5842) );
  nand2_2 U5594 ( .ip1(n5852), .ip2(n5338), .op(n6077) );
  nand2_2 U5595 ( .ip1(n5808), .ip2(n5807), .op(n5852) );
  nor2_4 U5596 ( .ip1(n5887), .ip2(n5754), .op(n10355) );
  nand2_2 U5597 ( .ip1(n5433), .ip2(n5753), .op(n5754) );
  nand2_2 U5598 ( .ip1(n5845), .ip2(n5407), .op(n5846) );
  nor2_2 U5599 ( .ip1(n5847), .ip2(n5846), .op(n5881) );
  inv_2 U5600 ( .ip(n5839), .op(n5263) );
  buf_1 U5601 ( .ip(n5328), .op(n5252) );
  nor2_1 U5602 ( .ip1(n5608), .ip2(n5253), .op(n5672) );
  nor2_2 U5603 ( .ip1(n5601), .ip2(n5602), .op(n5253) );
  buf_2 U5604 ( .ip(i_ssi_start_xfer), .op(n10288) );
  or2_4 U5605 ( .ip1(n6085), .ip2(n6188), .op(n6168) );
  inv_4 U5606 ( .ip(n5300), .op(n5264) );
  nand2_2 U5607 ( .ip1(n5408), .ip2(n5618), .op(n5733) );
  inv_2 U5608 ( .ip(n5329), .op(n5804) );
  nand2_2 U5609 ( .ip1(n5852), .ip2(n5809), .op(n5354) );
  nand2_4 U5610 ( .ip1(n5354), .ip2(n6188), .op(n6143) );
  inv_2 U5611 ( .ip(n5571), .op(n5594) );
  nand3_2 U5612 ( .ip1(n5595), .ip2(n5423), .ip3(n5594), .op(n5597) );
  nand3_2 U5613 ( .ip1(n5624), .ip2(n5600), .ip3(n5599), .op(n5602) );
  nor2_2 U5614 ( .ip1(n5803), .ip2(n5802), .op(n5674) );
  nand2_2 U5615 ( .ip1(n5804), .ip2(n5435), .op(n5850) );
  nand2_2 U5616 ( .ip1(n5299), .ip2(n5481), .op(n5606) );
  nand2_2 U5617 ( .ip1(n5606), .ip2(n5539), .op(n5578) );
  inv_4 U5618 ( .ip(n6143), .op(n10349) );
  nand2_1 U5619 ( .ip1(n8181), .ip2(i_i2c_ic_fs_spklen[0]), .op(n8182) );
  nand2_1 U5620 ( .ip1(n8135), .ip2(n8034), .op(n8035) );
  mux2_2 U5621 ( .ip1(i_i2c_ic_fs_lcnt[0]), .ip2(i_i2c_ic_lcnt[0]), .s(n6717), 
        .op(n7943) );
  nor3_1 U5622 ( .ip1(n6446), .ip2(n6445), .ip3(n6444), .op(n6447) );
  nand4_1 U5623 ( .ip1(n6480), .ip2(n6479), .ip3(n6478), .ip4(n9414), .op(
        n6481) );
  nor4_1 U5624 ( .ip1(i_i2c_ic_sda_tx_hold_sync[9]), .ip2(
        i_i2c_ic_sda_tx_hold_sync[15]), .ip3(i_i2c_ic_sda_tx_hold_sync[14]), 
        .ip4(n7124), .op(n7200) );
  or2_2 U5625 ( .ip1(n6077), .ip2(n5261), .op(n6040) );
  nand4_1 U5626 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[3]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[2]), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[1]), .ip4(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[0]), .op(n10424) );
  nand4_1 U5627 ( .ip1(n6943), .ip2(n6942), .ip3(n9737), .ip4(n8333), .op(
        n6944) );
  inv_1 U5628 ( .ip(i_apb_U_DW_apb_ahbsif_nextstate[0]), .op(n10009) );
  nor4_1 U5629 ( .ip1(i_apb_paddr[31]), .ip2(i_apb_paddr[29]), .ip3(n5862), 
        .ip4(n5861), .op(n5863) );
  nand4_1 U5630 ( .ip1(i_i2c_ic_data_oe), .ip2(n8554), .ip3(n8551), .ip4(
        i_i2c_slv_rxbyte_rdy), .op(n8536) );
  inv_1 U5631 ( .ip(i_i2c_mst_debug_cstate[3]), .op(n6905) );
  nor2_1 U5632 ( .ip1(n6881), .ip2(n6913), .op(n6880) );
  inv_1 U5633 ( .ip(n9379), .op(n10108) );
  nor2_1 U5634 ( .ip1(n8390), .ip2(n5867), .op(n9356) );
  nand3_1 U5635 ( .ip1(n9988), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[6]), .ip3(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[7]), .op(n10058) );
  inv_1 U5636 ( .ip(i_apb_U_DW_apb_ahbsif_nextstate[1]), .op(n10017) );
  nand4_1 U5637 ( .ip1(n5866), .ip2(n5865), .ip3(n5864), .ip4(n5863), .op(
        n8390) );
  nor3_1 U5638 ( .ip1(n10422), .ip2(n10423), .ip3(n10421), .op(n11065) );
  nand2_1 U5639 ( .ip1(n10198), .ip2(n11543), .op(n11555) );
  nand4_1 U5640 ( .ip1(n5325), .ip2(n11222), .ip3(n5326), .ip4(n11226), .op(
        n5324) );
  nor3_1 U5641 ( .ip1(i_ssi_tx_wr_addr[2]), .ip2(i_ssi_tx_wr_addr[1]), .ip3(
        n11211), .op(n10031) );
  nor3_1 U5642 ( .ip1(n6599), .ip2(n6598), .ip3(n7778), .op(n11598) );
  buf_1 U5643 ( .ip(n9356), .op(n9335) );
  and2_2 U5644 ( .ip1(n11370), .ip2(n11369), .op(n11408) );
  nand2_1 U5645 ( .ip1(n11358), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_htrans[1]), 
        .op(n9379) );
  nor3_1 U5646 ( .ip1(i_ahb_U_mux_hsel_prev[3]), .ip2(i_ahb_U_mux_hsel_prev[4]), .ip3(n11356), .op(n9358) );
  nor4_1 U5647 ( .ip1(i_ahb_U_mux_hsel_prev[3]), .ip2(i_ahb_U_mux_hsel_prev[2]), .ip3(i_ahb_U_mux_hsel_prev[4]), .ip4(n9195), .op(n9359) );
  inv_1 U5648 ( .ip(n10047), .op(n11226) );
  inv_1 U5649 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[4]), .op(
        n10558) );
  nand4_1 U5650 ( .ip1(n6985), .ip2(n6984), .ip3(n6983), .ip4(n6982), .op(
        n10480) );
  nor3_1 U5651 ( .ip1(i_apb_paddr[12]), .ip2(n8390), .ip3(n7434), .op(n11762)
         );
  nor2_1 U5652 ( .ip1(n11082), .ip2(n11081), .op(n11083) );
  and2_1 U5653 ( .ip1(n10623), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[12]), .op(n10626) );
  nand4_1 U5654 ( .ip1(n9666), .ip2(n9446), .ip3(n9445), .ip4(n9444), .op(
        n9447) );
  nand4_1 U5655 ( .ip1(n9666), .ip2(n9452), .ip3(n9451), .ip4(n9450), .op(
        n9453) );
  nor2_2 U5656 ( .ip1(n10935), .ip2(n7964), .op(n10936) );
  nor2_1 U5657 ( .ip1(n10820), .ip2(n10838), .op(n10815) );
  nor4_1 U5658 ( .ip1(i_i2c_tx_wr_addr[2]), .ip2(i_i2c_tx_wr_addr[1]), .ip3(
        i_i2c_tx_wr_addr[0]), .ip4(n9783), .op(n9616) );
  nor4_1 U5659 ( .ip1(i_i2c_tx_wr_addr[2]), .ip2(i_i2c_tx_wr_addr[0]), .ip3(
        n11253), .ip4(n9783), .op(n9615) );
  inv_1 U5660 ( .ip(n6655), .op(n5266) );
  inv_2 U5661 ( .ip(n5739), .op(n10261) );
  and2_2 U5662 ( .ip1(n10165), .ip2(n11214), .op(n9696) );
  buf_1 U5663 ( .ip(i_ssi_baudr[11]), .op(n6224) );
  inv_1 U5664 ( .ip(n11369), .op(n11427) );
  nor3_1 U5665 ( .ip1(n7920), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[13]), 
        .ip3(n9070), .op(n11358) );
  inv_1 U5666 ( .ip(n11355), .op(n7920) );
  inv_1 U5667 ( .ip(n7920), .op(ex_i_ahb_AHB_Slave_PID_hready) );
  inv_4 U5668 ( .ip(i_ssi_baudr[9]), .op(n6238) );
  nor2_4 U5669 ( .ip1(n6248), .ip2(n6214), .op(n6228) );
  nand2_4 U5670 ( .ip1(n5267), .ip2(n9089), .op(n6248) );
  nor3_4 U5671 ( .ip1(i_ssi_baudr[11]), .ip2(i_ssi_baudr[12]), .ip3(n6232), 
        .op(n6226) );
  nand2_4 U5672 ( .ip1(n6225), .ip2(n6238), .op(n6232) );
  nand2_4 U5673 ( .ip1(n6213), .ip2(n6212), .op(n6253) );
  inv_2 U5674 ( .ip(i_ssi_baudr[1]), .op(n6213) );
  inv_2 U5675 ( .ip(i_ssi_baudr[2]), .op(n6212) );
  nor2_2 U5676 ( .ip1(i_ssi_baudr[4]), .ip2(i_ssi_baudr[3]), .op(n9089) );
  inv_2 U5677 ( .ip(i_ssi_baudr[7]), .op(n5254) );
  inv_1 U5678 ( .ip(n5254), .op(n5255) );
  inv_2 U5679 ( .ip(n5254), .op(n5256) );
  nand2_2 U5680 ( .ip1(n10373), .ip2(n5439), .op(n10374) );
  inv_2 U5681 ( .ip(i_ssi_baudr[10]), .op(n6225) );
  nor2_2 U5682 ( .ip1(n10361), .ip2(n10374), .op(n10408) );
  buf_1 U5683 ( .ip(i_ssi_baudr[10]), .op(n5257) );
  xnor2_2 U5684 ( .ip1(n10310), .ip2(n6253), .op(n6243) );
  inv_2 U5685 ( .ip(n6253), .op(n5267) );
  and2_2 U5686 ( .ip1(n10409), .ip2(n11569), .op(n5307) );
  nand2_2 U5687 ( .ip1(n10408), .ip2(n10407), .op(n10409) );
  xor2_2 U5688 ( .ip1(i_ssi_U_mstfsm_frame_cnt[13]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[13]), .op(n5510) );
  xor2_2 U5689 ( .ip1(i_ssi_U_mstfsm_frame_cnt[11]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[11]), .op(n5509) );
  xor2_2 U5690 ( .ip1(i_ssi_U_mstfsm_frame_cnt[7]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[7]), .op(n5499) );
  inv_2 U5691 ( .ip(n5258), .op(n5259) );
  nor3_4 U5692 ( .ip1(n10365), .ip2(n10372), .ip3(n5259), .op(n10373) );
  nor2_2 U5693 ( .ip1(n10812), .ip2(n10898), .op(n10810) );
  nand2_2 U5694 ( .ip1(n10811), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[10]), .op(n10812) );
  nor2_2 U5695 ( .ip1(n10816), .ip2(n10886), .op(n10811) );
  nand2_2 U5696 ( .ip1(n10815), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[8]), .op(n10816) );
  nor2_2 U5697 ( .ip1(n10824), .ip2(n10864), .op(n10819) );
  and2_1 U5698 ( .ip1(n5678), .ip2(n5677), .op(n5679) );
  nor2_1 U5699 ( .ip1(n5429), .ip2(n5683), .op(n5677) );
  nor2_1 U5700 ( .ip1(n10263), .ip2(n5676), .op(n5683) );
  inv_2 U5701 ( .ip(n10899), .op(n10792) );
  nand2_1 U5702 ( .ip1(n5767), .ip2(n9712), .op(n5345) );
  nor2_1 U5703 ( .ip1(n10263), .ip2(n5676), .op(n5372) );
  nand3_1 U5704 ( .ip1(n6144), .ip2(n6132), .ip3(n5373), .op(n6195) );
  nand2_1 U5705 ( .ip1(n10302), .ip2(n10304), .op(n5676) );
  nor2_2 U5706 ( .ip1(n10355), .ip2(n6176), .op(n9712) );
  nor2_2 U5707 ( .ip1(n6182), .ip2(n10355), .op(n6208) );
  and2_1 U5708 ( .ip1(n5429), .ip2(n10263), .op(n5233) );
  nor2_1 U5709 ( .ip1(n5252), .ip2(n5675), .op(n10302) );
  nor2_2 U5710 ( .ip1(n5766), .ip2(n5765), .op(n6176) );
  nand2_1 U5711 ( .ip1(n10306), .ip2(n9984), .op(n5675) );
  inv_1 U5712 ( .ip(n6168), .op(n6177) );
  nand2_2 U5713 ( .ip1(n6115), .ip2(n5409), .op(n5765) );
  buf_1 U5714 ( .ip(n10306), .op(n5362) );
  and2_1 U5715 ( .ip1(n5354), .ip2(n5265), .op(n6152) );
  nand2_2 U5716 ( .ip1(n5842), .ip2(n5265), .op(n5300) );
  nand2_2 U5717 ( .ip1(n5764), .ip2(n5763), .op(n6115) );
  inv_1 U5718 ( .ip(n5763), .op(n10306) );
  inv_4 U5719 ( .ip(n5265), .op(n5377) );
  nand2_1 U5720 ( .ip1(n6056), .ip2(n6117), .op(n5766) );
  or2_1 U5721 ( .ip1(n5662), .ip2(n5661), .op(n10263) );
  nand2_2 U5722 ( .ip1(n5591), .ip2(n5590), .op(n5763) );
  and2_4 U5723 ( .ip1(n5795), .ip2(n5339), .op(n5306) );
  nor2_1 U5724 ( .ip1(n10537), .ip2(n5278), .op(n10540) );
  or3_2 U5725 ( .ip1(n5323), .ip2(n11221), .ip3(i_ssi_rx_wr_addr[1]), .op(
        n10049) );
  inv_2 U5726 ( .ip(n5739), .op(n5279) );
  inv_2 U5727 ( .ip(n9694), .op(n11211) );
  and4_2 U5728 ( .ip1(n5326), .ip2(n11222), .ip3(i_ssi_rx_wr_addr[2]), .ip4(
        n11226), .op(n9369) );
  inv_2 U5729 ( .ip(n5265), .op(n5260) );
  inv_2 U5730 ( .ip(n6188), .op(n5261) );
  and2_1 U5731 ( .ip1(n5739), .ip2(n6072), .op(n5891) );
  nand2_1 U5732 ( .ip1(n5747), .ip2(n5746), .op(n5836) );
  or4_2 U5733 ( .ip1(n11222), .ip2(n5325), .ip3(n10047), .ip4(
        i_ssi_rx_wr_addr[0]), .op(n9697) );
  and2_4 U5734 ( .ip1(n5698), .ip2(n5697), .op(n5739) );
  nor2_1 U5735 ( .ip1(n10400), .ip2(n10399), .op(n10404) );
  nor2_1 U5736 ( .ip1(n5579), .ip2(n5580), .op(n5327) );
  xor2_1 U5737 ( .ip1(n10317), .ip2(n10369), .op(n6258) );
  nand3_2 U5738 ( .ip1(n5578), .ip2(n5577), .ip3(n5632), .op(n5579) );
  nand2_1 U5739 ( .ip1(n6227), .ip2(n6228), .op(n6231) );
  nand2_2 U5740 ( .ip1(n6228), .ip2(n5406), .op(n10366) );
  nor3_2 U5741 ( .ip1(i_apb_paddr[12]), .ip2(n8390), .ip3(n8389), .op(
        i_i2c_wr_en) );
  and2_1 U5742 ( .ip1(n5606), .ip2(n5607), .op(n5608) );
  inv_2 U5743 ( .ip(n10198), .op(n5851) );
  nor3_2 U5744 ( .ip1(i_ssi_tx_rd_addr[0]), .ip2(i_ssi_tx_rd_addr[2]), .ip3(
        n5699), .op(n5769) );
  nand2_1 U5745 ( .ip1(n5299), .ip2(n9058), .op(n5690) );
  mux2_1 U5746 ( .ip1(i_i2c_ic_hs_spklen[1]), .ip2(i_i2c_ic_fs_spklen[1]), .s(
        n7384), .op(n7156) );
  nor2_2 U5747 ( .ip1(n5664), .ip2(n5663), .op(n5670) );
  inv_2 U5748 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r), .op(n7384) );
  nor4_2 U5749 ( .ip1(i_apb_paddr[26]), .ip2(i_apb_paddr[25]), .ip3(
        i_apb_paddr[23]), .ip4(i_apb_paddr[22]), .op(n5866) );
  nor2_2 U5750 ( .ip1(i_apb_U_DW_apb_ahbsif_state[1]), .ip2(
        i_apb_U_DW_apb_ahbsif_state[0]), .op(n9374) );
  inv_2 U5751 ( .ip(i_ssi_sclk_fe), .op(n5481) );
  nand2_1 U5752 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[9]), .ip2(
        n11083), .op(n11088) );
  nand2_1 U5753 ( .ip1(n6542), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[8]), .op(n10216) );
  inv_1 U5754 ( .ip(n10058), .op(n6542) );
  inv_1 U5755 ( .ip(n9982), .op(n9988) );
  nand2_1 U5756 ( .ip1(n10649), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[5]), .op(n10654) );
  nand2_1 U5757 ( .ip1(n10643), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[3]), .op(n10648) );
  and2_1 U5758 ( .ip1(n8878), .ip2(n10997), .op(n11006) );
  nand3_1 U5759 ( .ip1(n9956), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[3]), .ip3(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[4]), .op(n9980) );
  inv_1 U5760 ( .ip(n9944), .op(n9956) );
  nand2_1 U5761 ( .ip1(n6651), .ip2(n5472), .op(n9944) );
  nor2_1 U5762 ( .ip1(n8090), .ip2(n8089), .op(n8092) );
  nor2_1 U5763 ( .ip1(n6097), .ip2(n6096), .op(n6098) );
  nor3_1 U5764 ( .ip1(n6429), .ip2(n6430), .ip3(n6431), .op(n6369) );
  xnor2_1 U5765 ( .ip1(n8138), .ip2(n8137), .op(n8922) );
  nor2_1 U5766 ( .ip1(n5313), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[9]), .op(n6431) );
  and2_1 U5767 ( .ip1(n10356), .ip2(n6144), .op(n10357) );
  nand2_1 U5768 ( .ip1(n5364), .ip2(n6144), .op(n6107) );
  and2_1 U5769 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[9]), .ip2(n6154), 
        .op(n6153) );
  and2_1 U5770 ( .ip1(n6172), .ip2(n6170), .op(n5341) );
  buf_2 U5771 ( .ip(n11407), .op(n5271) );
  nor2_1 U5772 ( .ip1(n5297), .ip2(n5298), .op(n6540) );
  and2_1 U5773 ( .ip1(n5427), .ip2(n6193), .op(n6194) );
  inv_1 U5774 ( .ip(n9022), .op(n5272) );
  nor2_1 U5775 ( .ip1(n10265), .ip2(n5605), .op(n10334) );
  and2_1 U5776 ( .ip1(n5621), .ip2(n10265), .op(n5429) );
  and2_1 U5777 ( .ip1(n6061), .ip2(n9714), .op(n5848) );
  nand2_1 U5778 ( .ip1(n5841), .ip2(n5840), .op(n5847) );
  inv_2 U5779 ( .ip(n6800), .op(n5262) );
  nand2_1 U5780 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_buffer[4]), .ip2(n6177), 
        .op(n6062) );
  buf_1 U5781 ( .ip(n5306), .op(n5363) );
  or2_1 U5782 ( .ip1(n10341), .ip2(n5300), .op(n5407) );
  nor2_1 U5783 ( .ip1(n10248), .ip2(n6143), .op(n5991) );
  and2_1 U5784 ( .ip1(n5306), .ip2(n5875), .op(n5876) );
  nor2_1 U5785 ( .ip1(n5874), .ip2(n5300), .op(n5877) );
  nor3_1 U5786 ( .ip1(n8336), .ip2(n6648), .ip3(n6928), .op(n6946) );
  nor2_1 U5787 ( .ip1(n5620), .ip2(n5388), .op(n5621) );
  mux2_1 U5788 ( .ip1(i_i2c_ic_fs_hcnt[15]), .ip2(i_i2c_ic_hcnt[15]), .s(n5277), .op(n8046) );
  mux2_1 U5789 ( .ip1(i_i2c_ic_fs_hcnt[9]), .ip2(i_i2c_ic_hcnt[9]), .s(n5277), 
        .op(n8079) );
  mux2_1 U5790 ( .ip1(i_i2c_ic_fs_hcnt[10]), .ip2(i_i2c_ic_hcnt[10]), .s(n5277), .op(n8100) );
  mux2_1 U5791 ( .ip1(i_i2c_ic_fs_lcnt[8]), .ip2(i_i2c_ic_lcnt[8]), .s(n5277), 
        .op(n7979) );
  mux2_1 U5792 ( .ip1(i_i2c_ic_fs_hcnt[12]), .ip2(i_i2c_ic_hcnt[12]), .s(n5277), .op(n8070) );
  mux2_1 U5793 ( .ip1(i_i2c_ic_fs_lcnt[9]), .ip2(i_i2c_ic_lcnt[9]), .s(n5277), 
        .op(n7938) );
  mux2_1 U5794 ( .ip1(i_i2c_ic_fs_lcnt[11]), .ip2(i_i2c_ic_lcnt[11]), .s(n5277), .op(n7969) );
  nor2_1 U5795 ( .ip1(n6086), .ip2(n6085), .op(n6087) );
  mux2_1 U5796 ( .ip1(i_i2c_ic_fs_lcnt[13]), .ip2(i_i2c_ic_lcnt[13]), .s(n5277), .op(n7925) );
  nor2_1 U5797 ( .ip1(n5377), .ip2(n5333), .op(n6131) );
  inv_2 U5798 ( .ip(n10355), .op(n6144) );
  and2_1 U5799 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[2]), .ip2(n5260), 
        .op(n5837) );
  nand3_4 U5800 ( .ip1(n10048), .ip2(n5325), .ip3(n11222), .op(n10050) );
  and2_1 U5801 ( .ip1(n5260), .ip2(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[14]), .op(n5875) );
  nor2_1 U5802 ( .ip1(n5887), .ip2(n5886), .op(n10281) );
  and2_1 U5803 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[1]), .ip2(n5377), 
        .op(n5797) );
  inv_1 U5804 ( .ip(n10265), .op(n10304) );
  nor3_1 U5805 ( .ip1(n5623), .ip2(n6137), .ip3(n5622), .op(n5662) );
  or2_1 U5806 ( .ip1(n5301), .ip2(n5553), .op(n10265) );
  nor2_1 U5807 ( .ip1(n5383), .ip2(n5382), .op(n5409) );
  nand2_1 U5808 ( .ip1(n5356), .ip2(n5308), .op(n5796) );
  nand2_1 U5809 ( .ip1(n6056), .ip2(n5337), .op(n5886) );
  nor2_1 U5810 ( .ip1(n10406), .ip2(n10405), .op(n10407) );
  nand2_1 U5811 ( .ip1(n5794), .ip2(n5328), .op(n5741) );
  nand2_1 U5812 ( .ip1(n9708), .ip2(n5758), .op(n6056) );
  inv_1 U5813 ( .ip(n10536), .op(n5278) );
  and2_1 U5814 ( .ip1(n10232), .ip2(n5370), .op(n5301) );
  nor2_1 U5815 ( .ip1(n5329), .ip2(n5806), .op(n5808) );
  nand2_1 U5816 ( .ip1(n5735), .ip2(i_ssi_cfs[1]), .op(n5738) );
  inv_2 U5817 ( .ip(n5836), .op(n5265) );
  and2_1 U5818 ( .ip1(n10232), .ip2(n5594), .op(n5622) );
  inv_1 U5819 ( .ip(n11776), .op(n10584) );
  nand2_1 U5820 ( .ip1(n5554), .ip2(n5561), .op(n5591) );
  xor2_2 U5821 ( .ip1(n6237), .ip2(n10378), .op(n6239) );
  xor2_1 U5822 ( .ip1(n10379), .ip2(n10378), .op(n10393) );
  inv_2 U5823 ( .ip(n10278), .op(n10346) );
  mux2_2 U5824 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_scl_clk_int), .ip2(n8437), 
        .s(n6463), .op(n11776) );
  nor2_1 U5825 ( .ip1(n6304), .ip2(n6303), .op(n10528) );
  nand2_1 U5826 ( .ip1(n5743), .ip2(n5742), .op(n5736) );
  nand2_1 U5827 ( .ip1(n6234), .ip2(n6233), .op(n10375) );
  xor2_2 U5828 ( .ip1(n10370), .ip2(n10369), .op(n10371) );
  and2_1 U5829 ( .ip1(n10340), .ip2(n5811), .op(n5337) );
  nor2_1 U5830 ( .ip1(n5560), .ip2(n5559), .op(n5755) );
  nor2_1 U5831 ( .ip1(n5508), .ip2(n5507), .op(n5303) );
  nand2_1 U5832 ( .ip1(n9832), .ip2(n11598), .op(n11165) );
  nor2_2 U5833 ( .ip1(n9379), .ip2(n9382), .op(n11359) );
  nand2_1 U5834 ( .ip1(n5733), .ip2(n5734), .op(n5742) );
  or2_1 U5835 ( .ip1(n10366), .ip2(i_ssi_baudr[13]), .op(n10369) );
  inv_1 U5836 ( .ip(n9660), .op(n9832) );
  nor3_1 U5837 ( .ip1(i_ssi_baudr[13]), .ip2(i_ssi_baudr[14]), .ip3(n10366), 
        .op(n10367) );
  xor2_1 U5838 ( .ip1(n5256), .ip2(n10380), .op(n6254) );
  nand2_1 U5839 ( .ip1(n5573), .ip2(n5572), .op(n5580) );
  nand2_1 U5840 ( .ip1(n5672), .ip2(n5673), .op(n5802) );
  nand2_1 U5841 ( .ip1(n10397), .ip2(n9088), .op(n10380) );
  and2_1 U5842 ( .ip1(n5555), .ip2(n5558), .op(n5534) );
  inv_1 U5843 ( .ip(n5733), .op(n5731) );
  and2_1 U5844 ( .ip1(n5636), .ip2(n5612), .op(n5613) );
  nand3_1 U5845 ( .ip1(n5670), .ip2(n5669), .ip3(n5668), .op(n5673) );
  and2_1 U5846 ( .ip1(n5733), .ip2(n5399), .op(n5619) );
  nand2_1 U5847 ( .ip1(n9335), .ip2(n7433), .op(n9660) );
  nand2_1 U5848 ( .ip1(n5575), .ip2(n5571), .op(n5572) );
  inv_1 U5849 ( .ip(n9740), .op(n9725) );
  nor2_1 U5850 ( .ip1(n5667), .ip2(n5666), .op(n5668) );
  inv_1 U5851 ( .ip(n6659), .op(n5764) );
  nor2_1 U5852 ( .ip1(n5494), .ip2(n5493), .op(n5557) );
  nor2_1 U5853 ( .ip1(i_ssi_baudr[4]), .ip2(n10382), .op(n10397) );
  nor2_1 U5854 ( .ip1(n5576), .ip2(n5410), .op(n5577) );
  and2_1 U5855 ( .ip1(n5575), .ip2(n5281), .op(n5554) );
  nand2_1 U5856 ( .ip1(n5492), .ip2(n5491), .op(n5493) );
  inv_1 U5857 ( .ip(n5606), .op(n5571) );
  nand2_1 U5858 ( .ip1(n5355), .ip2(n10231), .op(n5632) );
  and2_1 U5859 ( .ip1(n6226), .ip2(n6227), .op(n5406) );
  xor2_2 U5860 ( .ip1(n10321), .ip2(n6241), .op(n6242) );
  nor2_1 U5861 ( .ip1(n6905), .ip2(n10413), .op(n6469) );
  nor2_1 U5862 ( .ip1(n5287), .ip2(n5288), .op(n5286) );
  nor2_1 U5863 ( .ip1(n6335), .ip2(n7376), .op(n5285) );
  inv_1 U5864 ( .ip(n9093), .op(n6227) );
  nand2_1 U5865 ( .ip1(n6311), .ip2(n6867), .op(n6881) );
  nand2_1 U5866 ( .ip1(n7380), .ip2(n6334), .op(n7376) );
  nor2_2 U5867 ( .ip1(i_ssi_tx_rd_addr[0]), .ip2(n5705), .op(n5817) );
  nor2_2 U5868 ( .ip1(n6971), .ip2(n5705), .op(n5812) );
  mux2_1 U5869 ( .ip1(i_i2c_ic_fs_spklen[0]), .ip2(i_i2c_ic_hs_spklen[0]), .s(
        n7672), .op(n7154) );
  nand2_2 U5870 ( .ip1(i_i2c_mst_debug_cstate[0]), .ip2(n6632), .op(n10413) );
  nand2_1 U5871 ( .ip1(n6317), .ip2(n6316), .op(n7400) );
  nor2_1 U5872 ( .ip1(n10288), .ip2(n9850), .op(n5609) );
  nand2_1 U5873 ( .ip1(n7591), .ip2(n6211), .op(n9093) );
  nand2_1 U5874 ( .ip1(n5592), .ip2(i_ssi_sclk_re), .op(n5599) );
  nor2_2 U5875 ( .ip1(i_ssi_tx_rd_addr[0]), .ip2(n9953), .op(n5819) );
  nor2_2 U5876 ( .ip1(i_ssi_tx_rd_addr[2]), .ip2(n5706), .op(n5818) );
  inv_2 U5877 ( .ip(n5413), .op(n11760) );
  nand2_1 U5878 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[7]), 
        .ip2(n6507), .op(n7380) );
  and2_1 U5879 ( .ip1(n10507), .ip2(i_ssi_U_regfile_ctrlr1_int[3]), .op(n5502)
         );
  nand2_1 U5880 ( .ip1(i_i2c_ic_fs_spklen[5]), .ip2(n8251), .op(n6317) );
  inv_1 U5881 ( .ip(n10288), .op(n5400) );
  nand2_1 U5882 ( .ip1(i_i2c_ic_fs_spklen[4]), .ip2(n10558), .op(n6316) );
  xor2_1 U5883 ( .ip1(i_ssi_U_mstfsm_bit_cnt[3]), .ip2(i_ssi_dfs[3]), .op(
        n5665) );
  inv_1 U5884 ( .ip(n5255), .op(n7591) );
  inv_1 U5885 ( .ip(i_ssi_sclk_re), .op(n9058) );
  inv_2 U5886 ( .ip(i_ssi_baud2), .op(n5299) );
  inv_1 U5887 ( .ip(i_ssi_tmod[1]), .op(n5689) );
  inv_1 U5888 ( .ip(i_ssi_start_xfer), .op(n5592) );
  xor2_1 U5889 ( .ip1(i_i2c_ic_hs_spklen[0]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[0]), .op(n5288) );
  buf_1 U5890 ( .ip(i_ssi_U_regfile_ctrlr1_int[15]), .op(n5394) );
  inv_1 U5891 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[1]), .op(
        n7362) );
  inv_1 U5892 ( .ip(i_ssi_mwcr[1]), .op(n9850) );
  nor2_1 U5893 ( .ip1(n10955), .ip2(n8210), .op(n5135) );
  nor2_1 U5894 ( .ip1(n10677), .ip2(n8724), .op(n5067) );
  nor2_2 U5895 ( .ip1(n10680), .ip2(n10679), .op(n10678) );
  nand2_2 U5896 ( .ip1(n10673), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[13]), .op(n10680) );
  nand2_1 U5897 ( .ip1(n6545), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[11]), .op(n10242) );
  nor2_2 U5898 ( .ip1(n10672), .ip2(n10671), .op(n10673) );
  nor2_1 U5899 ( .ip1(n10630), .ip2(n8388), .op(n5170) );
  nor2_2 U5900 ( .ip1(n11035), .ip2(n11034), .op(n11036) );
  nand2_2 U5901 ( .ip1(n11030), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[11]), .op(n11035) );
  nand2_2 U5902 ( .ip1(n10667), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[11]), .op(n10672) );
  nor2_2 U5903 ( .ip1(n10666), .ip2(n10665), .op(n10667) );
  nor2_2 U5904 ( .ip1(n11029), .ip2(n11028), .op(n11030) );
  nand2_1 U5905 ( .ip1(n6543), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[9]), .op(n10228) );
  nand2_2 U5906 ( .ip1(n10661), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[9]), .op(n10666) );
  nand2_2 U5907 ( .ip1(n11024), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[9]), .op(n11029) );
  inv_1 U5908 ( .ip(n11088), .op(n11084) );
  inv_1 U5909 ( .ip(n10216), .op(n6543) );
  nor2_2 U5910 ( .ip1(n11023), .ip2(n11022), .op(n11024) );
  nor2_2 U5911 ( .ip1(n10660), .ip2(n10659), .op(n10661) );
  nand2_2 U5912 ( .ip1(n10655), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[7]), .op(n10660) );
  nand2_2 U5913 ( .ip1(n11018), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[7]), .op(n11023) );
  nor2_1 U5914 ( .ip1(n10425), .ip2(n7357), .op(n11056) );
  nor2_2 U5915 ( .ip1(n11017), .ip2(n11016), .op(n11018) );
  nor2_2 U5916 ( .ip1(n10654), .ip2(n10653), .op(n10655) );
  nand2_2 U5917 ( .ip1(n11012), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[5]), .op(n11017) );
  nor2_1 U5918 ( .ip1(n10974), .ip2(n10973), .op(n10975) );
  nor2_2 U5919 ( .ip1(n11011), .ip2(n11010), .op(n11012) );
  nor2_2 U5920 ( .ip1(n10648), .ip2(n10647), .op(n10649) );
  nand2_2 U5921 ( .ip1(n10926), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[3]), .op(n10930) );
  nand2_1 U5922 ( .ip1(n9052), .ip2(n9051), .op(n10958) );
  nand2_2 U5923 ( .ip1(n11006), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[3]), .op(n11011) );
  and2_1 U5924 ( .ip1(n8723), .ip2(n10634), .op(n10643) );
  inv_1 U5925 ( .ip(n9980), .op(n6459) );
  nand2_1 U5926 ( .ip1(n8722), .ip2(n8721), .op(n10634) );
  nand2_1 U5927 ( .ip1(n8877), .ip2(n8876), .op(n10997) );
  inv_1 U5928 ( .ip(n6969), .op(n6651) );
  nand2_1 U5929 ( .ip1(n9935), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[0]), .op(n6969) );
  and2_1 U5930 ( .ip1(n10590), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[1]), .op(n10593) );
  and2_1 U5931 ( .ip1(n8387), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[0]), 
        .op(n10590) );
  and2_1 U5932 ( .ip1(n9040), .ip2(n9039), .op(n9041) );
  nor2_1 U5933 ( .ip1(n6456), .ip2(n6457), .op(n9935) );
  nor2_1 U5934 ( .ip1(n8668), .ip2(n8667), .op(n8680) );
  nor2_1 U5935 ( .ip1(n8817), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[11]), .op(n8106) );
  and2_1 U5936 ( .ip1(n7848), .ip2(n7847), .op(n7849) );
  nor2_1 U5937 ( .ip1(n8895), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[10]), .op(n8668) );
  xnor2_1 U5938 ( .ip1(n8092), .ip2(n8091), .op(n8817) );
  xnor2_1 U5939 ( .ip1(n8052), .ip2(n8051), .op(n8881) );
  xnor2_1 U5940 ( .ip1(n8079), .ip2(n8081), .op(n8897) );
  xnor2_1 U5941 ( .ip1(n8072), .ip2(n8071), .op(n8888) );
  xnor2_1 U5942 ( .ip1(n8102), .ip2(n8101), .op(n8895) );
  xnor2_1 U5943 ( .ip1(n8064), .ip2(n8063), .op(n8887) );
  xnor2_1 U5944 ( .ip1(n8046), .ip2(n8045), .op(n8880) );
  nor2_1 U5945 ( .ip1(n8088), .ip2(n8087), .op(n8089) );
  nor2_1 U5946 ( .ip1(n8133), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[7]), .op(n8841) );
  nor2_1 U5947 ( .ip1(n8099), .ip2(n8098), .op(n8102) );
  nor2_1 U5948 ( .ip1(n6749), .ip2(n6748), .op(n6828) );
  nand2_1 U5949 ( .ip1(n6362), .ip2(n6439), .op(n6450) );
  xnor2_1 U5950 ( .ip1(n8150), .ip2(n8149), .op(n8928) );
  nor2_1 U5951 ( .ip1(n6382), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[11]), .op(n6383) );
  inv_1 U5952 ( .ip(n6378), .op(n6382) );
  nor2_1 U5953 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[13]), .ip2(
        n10711), .op(n10777) );
  nor3_1 U5954 ( .ip1(n6409), .ip2(n6408), .ip3(n6410), .op(n6395) );
  nand2_1 U5955 ( .ip1(n11242), .ip2(n11241), .op(n11243) );
  nand2_1 U5956 ( .ip1(n6441), .ip2(n6442), .op(n6362) );
  nand2_1 U5957 ( .ip1(n6443), .ip2(n6361), .op(n6439) );
  nand3_1 U5958 ( .ip1(n6095), .ip2(n6094), .ip3(n6093), .op(n6096) );
  inv_2 U5959 ( .ip(n10907), .op(n10711) );
  xor2_2 U5960 ( .ip1(i_i2c_tx_abrt_flg), .ip2(n5296), .op(n5293) );
  nor2_1 U5961 ( .ip1(n7880), .ip2(n11082), .op(n7881) );
  or2_1 U5962 ( .ip1(n11240), .ip2(n11239), .op(n11241) );
  nor2_1 U5963 ( .ip1(n8128), .ip2(n8127), .op(n8132) );
  nor2_1 U5964 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[7]), .ip2(n6424), .op(n6421) );
  xnor2_1 U5965 ( .ip1(n8094), .ip2(n6368), .op(n5313) );
  xor2_1 U5966 ( .ip1(n8003), .ip2(n6365), .op(n6366) );
  nand2_1 U5967 ( .ip1(n6071), .ip2(n6070), .op(n6095) );
  nor2_1 U5968 ( .ip1(i_i2c_U_DW_apb_i2c_toggle_tx_abrt_r), .ip2(n6540), .op(
        n5296) );
  inv_1 U5969 ( .ip(n6415), .op(n6424) );
  nand2_1 U5970 ( .ip1(n6376), .ip2(n6364), .op(n6365) );
  nor4_1 U5971 ( .ip1(n6401), .ip2(n6403), .ip3(n6400), .ip4(n6399), .op(n6406) );
  nand2_1 U5972 ( .ip1(n11238), .ip2(n11237), .op(n11240) );
  inv_1 U5973 ( .ip(n6195), .op(n5268) );
  nand4_1 U5974 ( .ip1(n6062), .ip2(n6064), .ip3(n6065), .ip4(n6063), .op(
        n6067) );
  inv_1 U5975 ( .ip(n7321), .op(n7248) );
  nor2_2 U5976 ( .ip1(n6349), .ip2(n6390), .op(n6376) );
  nor2_1 U5977 ( .ip1(n6363), .ip2(n8070), .op(n6364) );
  xnor2_1 U5978 ( .ip1(n8173), .ip2(n8172), .op(n8935) );
  inv_1 U5979 ( .ip(n5298), .op(n9182) );
  nor2_1 U5980 ( .ip1(n8059), .ip2(n8063), .op(n8041) );
  nand2_1 U5981 ( .ip1(n6347), .ip2(n6416), .op(n6349) );
  nor2_1 U5982 ( .ip1(n8040), .ip2(n8093), .op(n8090) );
  nand2_1 U5983 ( .ip1(n5295), .ip2(n5294), .op(n5298) );
  nand2_1 U5984 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_buffer[12]), .ip2(n6177), 
        .op(n6052) );
  nand2_1 U5985 ( .ip1(n6756), .ip2(n6722), .op(n6738) );
  nand2_1 U5986 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_buffer[7]), .ip2(n10349), 
        .op(n6064) );
  xnor2_1 U5987 ( .ip1(n8180), .ip2(n8182), .op(n8939) );
  nand2_1 U5988 ( .ip1(n6373), .ip2(n6350), .op(n6363) );
  nor2_1 U5989 ( .ip1(n7989), .ip2(n7969), .op(n6722) );
  inv_1 U5990 ( .ip(n8003), .op(n8063) );
  nor2_2 U5991 ( .ip1(n8039), .ip2(n8079), .op(n6373) );
  nor2_1 U5992 ( .ip1(n8021), .ip2(n8023), .op(n6347) );
  nand2_1 U5993 ( .ip1(n6946), .ip2(n6841), .op(n5295) );
  nor2_1 U5994 ( .ip1(n9153), .ip2(n6481), .op(n5294) );
  nand2_1 U5995 ( .ip1(n7200), .ip2(n7199), .op(n7201) );
  nand2_1 U5996 ( .ip1(n8178), .ip2(n8006), .op(n8171) );
  mux2_1 U5997 ( .ip1(i_i2c_ic_fs_hcnt[14]), .ip2(i_i2c_ic_hcnt[14]), .s(n6346), .op(n6356) );
  mux2_1 U5998 ( .ip1(i_i2c_ic_fs_hcnt[13]), .ip2(i_i2c_ic_hcnt[13]), .s(n6721), .op(n8003) );
  mux2_1 U5999 ( .ip1(i_i2c_ic_fs_hcnt[11]), .ip2(i_i2c_ic_hcnt[11]), .s(n6721), .op(n8065) );
  buf_4 U6000 ( .ip(n10064), .op(n5274) );
  or2_2 U6001 ( .ip1(n8021), .ip2(n8020), .op(n8129) );
  buf_4 U6002 ( .ip(n10065), .op(n5275) );
  mux2_1 U6003 ( .ip1(i_i2c_ic_fs_lcnt[15]), .ip2(i_i2c_ic_lcnt[15]), .s(n6346), .op(n7937) );
  mux2_1 U6004 ( .ip1(i_i2c_ic_fs_lcnt[10]), .ip2(i_i2c_ic_lcnt[10]), .s(n6721), .op(n7989) );
  mux2_1 U6005 ( .ip1(i_i2c_ic_fs_lcnt[12]), .ip2(i_i2c_ic_lcnt[12]), .s(n6721), .op(n7977) );
  mux2_1 U6006 ( .ip1(i_i2c_ic_fs_lcnt[14]), .ip2(i_i2c_ic_lcnt[14]), .s(n6721), .op(n7934) );
  and2_1 U6007 ( .ip1(n10355), .ip2(n10280), .op(n5859) );
  mux2_1 U6008 ( .ip1(i_i2c_ic_fs_hcnt[8]), .ip2(i_i2c_ic_hcnt[8]), .s(n6721), 
        .op(n8039) );
  mux2_2 U6009 ( .ip1(i_i2c_ic_hcnt[7]), .ip2(i_i2c_ic_fs_hcnt[7]), .s(n6720), 
        .op(n8021) );
  nand2_1 U6010 ( .ip1(n8012), .ip2(n8011), .op(n8169) );
  and2_1 U6011 ( .ip1(n5457), .ip2(n6277), .op(n6278) );
  nand2_1 U6012 ( .ip1(n5290), .ip2(n8266), .op(n6648) );
  nand2_1 U6013 ( .ip1(n11152), .ip2(n5291), .op(n5290) );
  inv_4 U6014 ( .ip(n10875), .op(n5276) );
  inv_4 U6015 ( .ip(n6720), .op(n5277) );
  and2_1 U6016 ( .ip1(n6276), .ip2(n6275), .op(n6277) );
  nand2_2 U6017 ( .ip1(i_ssi_rx_wr_addr[0]), .ip2(n11226), .op(n11221) );
  inv_1 U6018 ( .ip(n6616), .op(n8266) );
  nand2_1 U6019 ( .ip1(n5292), .ip2(n6465), .op(n11152) );
  xor2_1 U6020 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[12]), .ip2(n6229), .op(n6230) );
  inv_1 U6021 ( .ip(n10109), .op(n11473) );
  nand2_1 U6022 ( .ip1(n5478), .ip2(n5750), .op(n5753) );
  nor2_1 U6023 ( .ip1(n6662), .ip2(n6670), .op(n6664) );
  nand3_1 U6024 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_int_d), .ip2(n6464), 
        .ip3(n10584), .op(n5292) );
  inv_1 U6025 ( .ip(n10232), .op(n5750) );
  nand3_1 U6026 ( .ip1(n10394), .ip2(n10393), .ip3(n10392), .op(n10406) );
  nor2_2 U6027 ( .ip1(n11760), .ip2(n11124), .op(n10223) );
  nand2_2 U6028 ( .ip1(n11760), .ip2(n9368), .op(n10047) );
  nand2_1 U6029 ( .ip1(i_apb_U_DW_apb_ahbsif_nextstate[2]), .ip2(n10017), .op(
        n10105) );
  nand2_2 U6030 ( .ip1(n9690), .ip2(n11569), .op(n10051) );
  mux2_1 U6031 ( .ip1(i_apb_pwdata_int[7]), .ip2(i_ssi_U_regfile_ctrlr1_int[7]), .s(n9896), .op(n4603) );
  mux2_1 U6032 ( .ip1(n10005), .ip2(n11776), .s(
        i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv), .op(n11099) );
  nand2_1 U6033 ( .ip1(n11217), .ip2(i_ssi_tx_wr_addr[0]), .op(n9695) );
  nor3_1 U6034 ( .ip1(i_i2c_rx_push_sync), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[0]), .ip3(n11205), .op(n6670)
         );
  mux2_1 U6035 ( .ip1(n9072), .ip2(i_ssi_U_fifo_unconnected_tx_wrd_count[0]), 
        .s(i_ssi_U_fifo_unconnected_tx_wrd_count[1]), .op(n9073) );
  nand2_1 U6036 ( .ip1(n5674), .ip2(n5438), .op(n5807) );
  and2_1 U6037 ( .ip1(n10303), .ip2(n10288), .op(n10289) );
  inv_4 U6038 ( .ip(n10854), .op(n5280) );
  buf_1 U6039 ( .ip(n10366), .op(n5402) );
  inv_1 U6040 ( .ip(n11189), .op(n11205) );
  xnor2_1 U6041 ( .ip1(n10360), .ip2(n10375), .op(n10361) );
  nor2_1 U6042 ( .ip1(n6224), .ip2(n10375), .op(n10376) );
  xnor2_1 U6043 ( .ip1(n10364), .ip2(n10366), .op(n10365) );
  nand4_1 U6044 ( .ip1(n9314), .ip2(n9313), .ip3(n9312), .ip4(n9311), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[19]) );
  nand2_1 U6045 ( .ip1(n6314), .ip2(n5419), .op(n6345) );
  nand2_2 U6046 ( .ip1(n5448), .ip2(n6142), .op(n6655) );
  xor2_1 U6047 ( .ip1(n10368), .ip2(n10367), .op(n10372) );
  nand4_1 U6048 ( .ip1(n9299), .ip2(n9298), .ip3(n9297), .ip4(n9296), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[7]) );
  and2_1 U6049 ( .ip1(n6114), .ip2(n5752), .op(n5433) );
  inv_1 U6050 ( .ip(n9708), .op(n10278) );
  nand4_1 U6051 ( .ip1(n9209), .ip2(n9208), .ip3(n9207), .ip4(n9206), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[31]) );
  nand4_1 U6052 ( .ip1(n9269), .ip2(n9268), .ip3(n9267), .ip4(n9266), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[17]) );
  nand2_1 U6053 ( .ip1(n10499), .ip2(n10500), .op(n6303) );
  nand4_1 U6054 ( .ip1(n9214), .ip2(n9213), .ip3(n9212), .ip4(n9211), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[20]) );
  nand4_1 U6055 ( .ip1(n9204), .ip2(n9203), .ip3(n9202), .ip4(n9201), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[27]) );
  nand4_1 U6056 ( .ip1(n9274), .ip2(n9273), .ip3(n9272), .ip4(n9271), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[1]) );
  nor2_1 U6057 ( .ip1(n5247), .ip2(n11209), .op(n11189) );
  nand4_1 U6058 ( .ip1(n9284), .ip2(n9283), .ip3(n9282), .ip4(n9281), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[0]) );
  nand4_1 U6059 ( .ip1(n9340), .ip2(n9339), .ip3(n9338), .ip4(n9337), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[22]) );
  nand4_1 U6060 ( .ip1(n9229), .ip2(n9228), .ip3(n9227), .ip4(n9226), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[2]) );
  nand4_1 U6061 ( .ip1(n9264), .ip2(n9263), .ip3(n9262), .ip4(n9261), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[3]) );
  nand2_1 U6062 ( .ip1(n9897), .ip2(n6581), .op(
        i_apb_U_DW_apb_ahbsif_nextstate[1]) );
  nand4_1 U6063 ( .ip1(n9334), .ip2(n9333), .ip3(n9332), .ip4(n9331), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[26]) );
  nor2_1 U6064 ( .ip1(n5951), .ip2(n5950), .op(n10251) );
  nand4_1 U6065 ( .ip1(n9224), .ip2(n9223), .ip3(n9222), .ip4(n9221), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[16]) );
  nand2_1 U6066 ( .ip1(n5401), .ip2(n5557), .op(n5559) );
  nand4_1 U6067 ( .ip1(n9249), .ip2(n9248), .ip3(n9247), .ip4(n9246), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[10]) );
  nand4_1 U6068 ( .ip1(n9329), .ip2(n9328), .ip3(n9327), .ip4(n9326), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[23]) );
  nand4_1 U6069 ( .ip1(n9219), .ip2(n9218), .ip3(n9217), .ip4(n9216), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[13]) );
  nand4_1 U6070 ( .ip1(n9304), .ip2(n9303), .ip3(n9302), .ip4(n9301), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[18]) );
  and2_1 U6071 ( .ip1(n9608), .ip2(n9569), .op(n9570) );
  nand4_1 U6072 ( .ip1(n9345), .ip2(n9344), .ip3(n9343), .ip4(n9342), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[29]) );
  nand4_1 U6073 ( .ip1(n9364), .ip2(n9363), .ip3(n9362), .ip4(n9361), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[30]) );
  nand4_1 U6074 ( .ip1(n9350), .ip2(n9349), .ip3(n9348), .ip4(n9347), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[24]) );
  nand4_1 U6075 ( .ip1(n9289), .ip2(n9288), .ip3(n9287), .ip4(n9286), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[14]) );
  nand4_1 U6076 ( .ip1(n9239), .ip2(n9238), .ip3(n9237), .ip4(n9236), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[12]) );
  nand4_1 U6077 ( .ip1(n9259), .ip2(n9258), .ip3(n9257), .ip4(n9256), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[11]) );
  nand4_1 U6078 ( .ip1(n9324), .ip2(n9323), .ip3(n9322), .ip4(n9321), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[25]) );
  nand4_1 U6079 ( .ip1(n9254), .ip2(n9253), .ip3(n9252), .ip4(n9251), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[21]) );
  nand4_1 U6080 ( .ip1(n9319), .ip2(n9318), .ip3(n9317), .ip4(n9316), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[15]) );
  nor2_1 U6081 ( .ip1(n5790), .ip2(n5789), .op(n9707) );
  nand4_1 U6082 ( .ip1(n9309), .ip2(n9308), .ip3(n9307), .ip4(n9306), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[6]) );
  nand4_1 U6083 ( .ip1(n9244), .ip2(n9243), .ip3(n9242), .ip4(n9241), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[9]) );
  and2_1 U6084 ( .ip1(n5811), .ip2(n9717), .op(n6114) );
  inv_1 U6085 ( .ip(n10487), .op(n10499) );
  nand4_1 U6086 ( .ip1(n9279), .ip2(n9278), .ip3(n9277), .ip4(n9276), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[4]) );
  nor2_1 U6087 ( .ip1(n6015), .ip2(n6014), .op(n10254) );
  nand4_1 U6088 ( .ip1(n9355), .ip2(n9354), .ip3(n9353), .ip4(n9352), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[28]) );
  nand4_1 U6089 ( .ip1(n9294), .ip2(n9293), .ip3(n9292), .ip4(n9291), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[8]) );
  nand4_1 U6090 ( .ip1(n9234), .ip2(n9233), .ip3(n9232), .ip4(n9231), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[5]) );
  xor2_1 U6091 ( .ip1(n10401), .ip2(n10322), .op(n5457) );
  nand2_1 U6092 ( .ip1(n5646), .ip2(n5645), .op(n5732) );
  nor2_1 U6093 ( .ip1(n5533), .ip2(n5532), .op(n5401) );
  nand2_1 U6094 ( .ip1(n6296), .ip2(n6295), .op(n10487) );
  nor2_1 U6095 ( .ip1(n5521), .ip2(n5520), .op(n5555) );
  nor2_1 U6096 ( .ip1(n5289), .ip2(n5284), .op(n6336) );
  nor2_1 U6097 ( .ip1(n5505), .ip2(n5506), .op(n5556) );
  mux2_1 U6098 ( .ip1(i_i2c_prdata[9]), .ip2(i_ssi_prdata[9]), .s(n9356), .op(
        n9240) );
  mux2_1 U6099 ( .ip1(i_i2c_prdata[12]), .ip2(i_ssi_prdata[12]), .s(n9356), 
        .op(n9235) );
  mux2_1 U6100 ( .ip1(i_i2c_prdata[11]), .ip2(i_ssi_prdata[11]), .s(n9356), 
        .op(n9255) );
  mux2_1 U6101 ( .ip1(i_i2c_prdata[28]), .ip2(i_ssi_prdata[28]), .s(n9356), 
        .op(n9351) );
  nand2_1 U6102 ( .ip1(n5286), .ip2(n5285), .op(n5284) );
  mux2_1 U6103 ( .ip1(i_i2c_prdata[10]), .ip2(i_ssi_prdata[10]), .s(n9356), 
        .op(n9245) );
  nand2_1 U6104 ( .ip1(n5610), .ip2(n5609), .op(n5636) );
  mux2_1 U6105 ( .ip1(i_i2c_prdata[30]), .ip2(i_ssi_prdata[30]), .s(n9356), 
        .op(n9357) );
  nand2_1 U6106 ( .ip1(n7145), .ip2(n7144), .op(n7163) );
  nor2_2 U6107 ( .ip1(n7158), .ip2(n7157), .op(n7159) );
  and2_1 U6108 ( .ip1(i_ssi_mwcr[1]), .ip2(n5610), .op(n5539) );
  mux2_1 U6109 ( .ip1(i_i2c_prdata[21]), .ip2(i_ssi_prdata[21]), .s(n9356), 
        .op(n9250) );
  mux2_1 U6110 ( .ip1(i_i2c_prdata[23]), .ip2(i_ssi_prdata[23]), .s(n9356), 
        .op(n9325) );
  mux2_1 U6111 ( .ip1(i_i2c_prdata[24]), .ip2(i_ssi_prdata[24]), .s(n9356), 
        .op(n9346) );
  nand2_1 U6112 ( .ip1(n5531), .ip2(n5530), .op(n5532) );
  mux2_1 U6113 ( .ip1(i_i2c_prdata[25]), .ip2(i_ssi_prdata[25]), .s(n9356), 
        .op(n9320) );
  mux2_1 U6114 ( .ip1(i_i2c_prdata[8]), .ip2(i_ssi_prdata[8]), .s(n9356), .op(
        n9290) );
  mux2_1 U6115 ( .ip1(i_i2c_prdata[6]), .ip2(i_ssi_prdata[6]), .s(n9356), .op(
        n9305) );
  mux2_1 U6116 ( .ip1(i_i2c_prdata[5]), .ip2(i_ssi_prdata[5]), .s(n9356), .op(
        n9230) );
  mux2_1 U6117 ( .ip1(i_i2c_prdata[4]), .ip2(i_ssi_prdata[4]), .s(n9356), .op(
        n9275) );
  nand2_1 U6118 ( .ip1(n10489), .ip2(n5443), .op(n6304) );
  buf_1 U6119 ( .ip(n11762), .op(n7435) );
  mux2_1 U6120 ( .ip1(i_i2c_prdata[14]), .ip2(i_ssi_prdata[14]), .s(n9356), 
        .op(n9285) );
  mux2_1 U6121 ( .ip1(i_i2c_prdata[15]), .ip2(i_ssi_prdata[15]), .s(n9356), 
        .op(n9315) );
  mux2_1 U6122 ( .ip1(i_i2c_prdata[13]), .ip2(i_ssi_prdata[13]), .s(n9356), 
        .op(n9215) );
  mux2_1 U6123 ( .ip1(i_i2c_prdata[16]), .ip2(i_ssi_prdata[16]), .s(n9356), 
        .op(n9220) );
  mux2_1 U6124 ( .ip1(i_i2c_prdata[26]), .ip2(i_ssi_prdata[26]), .s(n9356), 
        .op(n9330) );
  mux2_1 U6125 ( .ip1(i_i2c_prdata[29]), .ip2(i_ssi_prdata[29]), .s(n9356), 
        .op(n9341) );
  mux2_1 U6126 ( .ip1(i_i2c_prdata[18]), .ip2(i_ssi_prdata[18]), .s(n9356), 
        .op(n9300) );
  nand2_1 U6127 ( .ip1(n5487), .ip2(n5486), .op(n5494) );
  nand2_1 U6128 ( .ip1(n5525), .ip2(n5524), .op(n5533) );
  and2_1 U6129 ( .ip1(n5376), .ip2(n9684), .op(n9685) );
  xnor2_1 U6130 ( .ip1(n5411), .ip2(n5267), .op(n10389) );
  inv_1 U6131 ( .ip(n7160), .op(n7144) );
  nor2_1 U6132 ( .ip1(n5482), .ip2(n5756), .op(n5757) );
  mux2_1 U6133 ( .ip1(i_ssi_U_mstfsm_bit_cnt[1]), .ip2(n6287), .s(n5398), .op(
        n10489) );
  nand4_2 U6134 ( .ip1(n6555), .ip2(n6554), .ip3(n6553), .ip4(n6552), .op(
        n11355) );
  nand4_1 U6135 ( .ip1(n9200), .ip2(n9199), .ip3(n9198), .ip4(n9197), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hresp[0]) );
  nand2_1 U6136 ( .ip1(n6319), .ip2(n6318), .op(n7396) );
  and3_1 U6137 ( .ip1(n10387), .ip2(i_ssi_U_sclkgen_ssi_cnt[0]), .ip3(n10386), 
        .op(n10388) );
  xnor2_1 U6138 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[3]), .ip2(n10310), .op(n5411)
         );
  nand2_1 U6139 ( .ip1(n7367), .ip2(i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r), 
        .op(n5287) );
  xnor2_1 U6140 ( .ip1(n5310), .ip2(n5523), .op(n5524) );
  nand2_1 U6141 ( .ip1(n7379), .ip2(n7365), .op(n5289) );
  mux2_1 U6142 ( .ip1(n9366), .ip2(n6293), .s(n5358), .op(n6294) );
  nor2_1 U6143 ( .ip1(i_i2c_ic_fs_spklen[5]), .ip2(n8251), .op(n7394) );
  mux2_1 U6144 ( .ip1(n7100), .ip2(n7099), .s(n7672), .op(n7180) );
  nand2_1 U6145 ( .ip1(n5616), .ip2(n5615), .op(n5618) );
  and2_1 U6146 ( .ip1(i_i2c_scl_lcnt_cmplt), .ip2(i_i2c_mst_rx_ack_vld), .op(
        n5291) );
  nand2_1 U6147 ( .ip1(n5640), .ip2(n5639), .op(n5734) );
  mux2_1 U6148 ( .ip1(n7118), .ip2(n7117), .s(n7672), .op(n7160) );
  and2_1 U6149 ( .ip1(n10535), .ip2(i_ssi_U_regfile_ctrlr1_int[12]), .op(n5511) );
  and2_1 U6150 ( .ip1(n10531), .ip2(i_ssi_U_regfile_ctrlr1_int[10]), .op(n5396) );
  and2_1 U6151 ( .ip1(n10539), .ip2(i_ssi_U_regfile_ctrlr1_int[13]), .op(n5310) );
  and2_1 U6152 ( .ip1(n10519), .ip2(i_ssi_U_regfile_ctrlr1_int[6]), .op(n5500)
         );
  nor2_1 U6153 ( .ip1(n5663), .ip2(n5665), .op(n5640) );
  and2_1 U6154 ( .ip1(n10527), .ip2(i_ssi_U_regfile_ctrlr1_int[9]), .op(n5527)
         );
  nor2_1 U6155 ( .ip1(i_ssi_U_mstfsm_bit_cnt[4]), .ip2(n5664), .op(n5639) );
  nor2_1 U6156 ( .ip1(n5722), .ip2(n5721), .op(n5723) );
  nand2_1 U6157 ( .ip1(n7362), .ip2(i_i2c_ic_hs_spklen[1]), .op(n7367) );
  nand2_1 U6158 ( .ip1(n6515), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[5]), .op(n7365) );
  nand2_1 U6159 ( .ip1(n8251), .ip2(i_i2c_ic_hs_spklen[5]), .op(n7379) );
  inv_1 U6160 ( .ip(n5315), .op(n5316) );
  nor2_1 U6161 ( .ip1(i_i2c_ic_hs_spklen[3]), .ip2(n10554), .op(n7370) );
  nor2_1 U6162 ( .ip1(i_i2c_ic_fs_spklen[2]), .ip2(n10552), .op(n7389) );
  inv_4 U6163 ( .ip(n11148), .op(n11569) );
  nor2_2 U6164 ( .ip1(n6867), .ip2(n6310), .op(n6632) );
  xor2_1 U6165 ( .ip1(i_ssi_baudr[4]), .ip2(n10441), .op(n10383) );
  inv_2 U6166 ( .ip(n7384), .op(n7672) );
  xnor2_1 U6167 ( .ip1(n10455), .ip2(n5257), .op(n6237) );
  buf_1 U6168 ( .ip(i_ssi_U_regfile_ctrlr1_int[1]), .op(n5395) );
  nor4_2 U6169 ( .ip1(i_apb_paddr[19]), .ip2(i_apb_paddr[21]), .ip3(
        i_apb_paddr[20]), .ip4(i_apb_paddr[18]), .op(n5865) );
  nor4_2 U6170 ( .ip1(i_apb_paddr[16]), .ip2(i_apb_paddr[15]), .ip3(
        i_apb_paddr[14]), .ip4(i_apb_paddr[13]), .op(n5864) );
  nor4_2 U6171 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[13]), .ip2(
        i_ssi_U_sclkgen_ssi_cnt[14]), .ip3(i_ssi_U_sclkgen_ssi_cnt[0]), .ip4(
        i_ssi_U_sclkgen_ssi_cnt[15]), .op(n10296) );
  xor2_1 U6172 ( .ip1(i_i2c_ic_fs_spklen[0]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[0]), .op(n6325) );
  inv_1 U6173 ( .ip(i_ssi_tx_rd_addr[0]), .op(n6971) );
  inv_1 U6174 ( .ip(i_ssi_rx_wr_addr[1]), .op(n11222) );
  inv_1 U6175 ( .ip(i_ssi_baudr[8]), .op(n6211) );
  or2_1 U6176 ( .ip1(i_i2c_mst_debug_cstate[2]), .ip2(
        i_i2c_mst_debug_cstate[4]), .op(n6310) );
  inv_1 U6177 ( .ip(i_ssi_rx_wr_addr[2]), .op(n5325) );
  xor2_1 U6178 ( .ip1(i_ssi_U_mstfsm_bit_cnt[2]), .ip2(i_ssi_dfs[2]), .op(
        n5667) );
  buf_1 U6179 ( .ip(i_ssi_U_regfile_ctrlr1_int[6]), .op(n5392) );
  inv_2 U6180 ( .ip(n5689), .op(n5281) );
  buf_1 U6181 ( .ip(i_ssi_U_regfile_ctrlr1_int[8]), .op(n5393) );
  inv_1 U6182 ( .ip(n6978), .op(n5282) );
  inv_1 U6183 ( .ip(i_i2c_ic_sda_tx_hold_sync[2]), .op(n7161) );
  nand3_1 U6184 ( .ip1(n9366), .ip2(n5283), .ip3(n6291), .op(n6292) );
  nand2_1 U6185 ( .ip1(i_ssi_U_mstfsm_bit_cnt[1]), .ip2(n10205), .op(n5283) );
  nor2_1 U6186 ( .ip1(n5990), .ip2(n5991), .op(n5992) );
  inv_2 U6187 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[5]), .op(
        n8251) );
  inv_1 U6188 ( .ip(n8282), .op(n5297) );
  nand2_1 U6189 ( .ip1(n5304), .ip2(n10337), .op(n10338) );
  nor2_1 U6190 ( .ip1(n10334), .ip2(n5305), .op(n5304) );
  nand2_1 U6191 ( .ip1(n10336), .ip2(n10335), .op(n5305) );
  nor2_1 U6192 ( .ip1(n10302), .ip2(n10301), .op(n10335) );
  nand3_1 U6193 ( .ip1(n5350), .ip2(n5745), .ip3(n5742), .op(n5746) );
  nand2_1 U6194 ( .ip1(n5733), .ip2(n5732), .op(n5350) );
  nor2_4 U6195 ( .ip1(n10275), .ip2(n6458), .op(n4162) );
  nor2_2 U6196 ( .ip1(n8029), .ip2(n8028), .op(n8151) );
  nand2_1 U6197 ( .ip1(n6459), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[5]), .op(n9982) );
  nand2_1 U6198 ( .ip1(n10684), .ip2(n10683), .op(n10748) );
  nand2_2 U6199 ( .ip1(n10819), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[6]), .op(n10820) );
  inv_4 U6200 ( .ip(i_i2c_ic_ss_sync), .op(n10719) );
  nor4_2 U6201 ( .ip1(n10799), .ip2(n10798), .ip3(n10914), .ip4(n10797), .op(
        n5450) );
  nor3_1 U6202 ( .ip1(n10732), .ip2(n10835), .ip3(n10731), .op(n10798) );
  xor2_1 U6203 ( .ip1(n10723), .ip2(n10724), .op(n10835) );
  xor2_2 U6204 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[15]), .ip2(
        n10273), .op(n6548) );
  nor2_1 U6205 ( .ip1(n10275), .ip2(n6548), .op(n4150) );
  xor2_2 U6206 ( .ip1(n11056), .ip2(n7358), .op(n5462) );
  nor2_1 U6207 ( .ip1(n11099), .ip2(n5462), .op(n4957) );
  nand2_1 U6208 ( .ip1(n5804), .ip2(n5432), .op(n5308) );
  nand2_1 U6209 ( .ip1(n5804), .ip2(n5432), .op(n5740) );
  inv_1 U6210 ( .ip(n5561), .op(n5309) );
  nand2_1 U6211 ( .ip1(n5519), .ip2(n5518), .op(n5520) );
  xor2_2 U6212 ( .ip1(n5517), .ip2(n5516), .op(n5518) );
  xor2_1 U6213 ( .ip1(n6231), .ip2(n6238), .op(n6260) );
  inv_1 U6214 ( .ip(n6231), .op(n10395) );
  xor2_1 U6215 ( .ip1(i_ssi_U_mstfsm_frame_cnt[14]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[14]), .op(n5523) );
  xor2_2 U6216 ( .ip1(n5489), .ip2(n5488), .op(n5492) );
  xor2_2 U6217 ( .ip1(n5485), .ip2(n5484), .op(n5486) );
  xor2_2 U6218 ( .ip1(n5515), .ip2(n5514), .op(n5519) );
  inv_4 U6219 ( .ip(i_apb_pclk_en), .op(n10106) );
  mux2_1 U6220 ( .ip1(n10106), .ip2(i_apb_pclk_en), .s(
        i_apb_U_DW_apb_ahbsif_piped_hwrite_c), .op(n6566) );
  nand2_1 U6221 ( .ip1(n6573), .ip2(n6572), .op(n5311) );
  not_ab_or_c_or_d U6222 ( .ip1(n6568), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite), .ip3(n6567), .ip4(n10020), .op(
        n5312) );
  nand2_1 U6223 ( .ip1(n5312), .ip2(n6572), .op(
        i_apb_U_DW_apb_ahbsif_nextstate[0]) );
  inv_4 U6224 ( .ip(n9397), .op(n9396) );
  inv_4 U6225 ( .ip(n9397), .op(n9398) );
  inv_4 U6226 ( .ip(n9395), .op(n9397) );
  nand2_1 U6227 ( .ip1(n8065), .ip2(n8070), .op(n8059) );
  nor2_1 U6228 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[13]), .ip2(
        n6447), .op(n6448) );
  nor2_4 U6229 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[13]), .ip2(
        n6366), .op(n6445) );
  inv_1 U6230 ( .ip(n7362), .op(n5314) );
  inv_1 U6231 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[6]), .op(
        n5315) );
  inv_1 U6232 ( .ip(n10558), .op(n5317) );
  inv_1 U6233 ( .ip(n5320), .op(n5318) );
  inv_1 U6234 ( .ip(n6529), .op(n5319) );
  inv_1 U6235 ( .ip(n8251), .op(n5320) );
  nand3_2 U6236 ( .ip1(n8437), .ip2(n6463), .ip3(n6465), .op(n6461) );
  nor2_1 U6237 ( .ip1(n6435), .ip2(n6389), .op(n6457) );
  inv_4 U6238 ( .ip(n6720), .op(n6346) );
  nand2_2 U6239 ( .ip1(n6339), .ip2(n6338), .op(n6463) );
  inv_4 U6240 ( .ip(n6717), .op(n6720) );
  nand2_1 U6241 ( .ip1(n10270), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[14]), .op(n10273) );
  nand2_2 U6242 ( .ip1(n6605), .ip2(n9071), .op(n10052) );
  nand2_2 U6243 ( .ip1(n6991), .ip2(n6604), .op(n6605) );
  inv_2 U6244 ( .ip(n9692), .op(n6972) );
  nand2_2 U6245 ( .ip1(n9074), .ip2(n6607), .op(n6608) );
  xnor2_2 U6246 ( .ip1(i_ssi_U_fifo_rx_push_edge), .ip2(i_ssi_rx_push), .op(
        n5413) );
  inv_1 U6247 ( .ip(i_ssi_rx_wr_addr[2]), .op(n5323) );
  xnor2_1 U6248 ( .ip1(n5321), .ip2(n6667), .op(n6989) );
  inv_1 U6249 ( .ip(i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[2]), .op(n5321) );
  inv_1 U6250 ( .ip(i_ssi_rx_wr_addr[0]), .op(n5326) );
  nand4_2 U6251 ( .ip1(n5323), .ip2(n5326), .ip3(i_ssi_rx_wr_addr[1]), .ip4(
        n11226), .op(n5322) );
  nand2_1 U6252 ( .ip1(n6718), .ip2(n6798), .op(n6766) );
  nor2_1 U6253 ( .ip1(n7949), .ip2(n7941), .op(n6718) );
  nand2_1 U6254 ( .ip1(n7254), .ip2(n7251), .op(n7243) );
  nand2_1 U6255 ( .ip1(n7272), .ip2(n7110), .op(n7252) );
  or2_1 U6256 ( .ip1(n7281), .ip2(n7271), .op(n7110) );
  nor2_1 U6257 ( .ip1(n7140), .ip2(n7139), .op(n7284) );
  nand2_1 U6258 ( .ip1(n7289), .ip2(n7121), .op(n7140) );
  or2_1 U6259 ( .ip1(n7297), .ip2(n7288), .op(n7121) );
  nor2_1 U6260 ( .ip1(n7105), .ip2(n7255), .op(n7114) );
  nand2_1 U6261 ( .ip1(n7870), .ip2(n7869), .op(n7902) );
  or2_1 U6262 ( .ip1(n7141), .ip2(n7284), .op(n7245) );
  nand2_1 U6263 ( .ip1(n7114), .ip2(n7265), .op(n7141) );
  nand2_1 U6264 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[3]), 
        .ip2(n6321), .op(n6318) );
  nand2_1 U6265 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[4]), 
        .ip2(n6487), .op(n6319) );
  nor2_1 U6266 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[6]), 
        .ip2(n7100), .op(n7404) );
  nand2_1 U6267 ( .ip1(n6380), .ip2(n6379), .op(n6428) );
  nand2_1 U6268 ( .ip1(n6384), .ip2(n6385), .op(n6380) );
  and2_1 U6269 ( .ip1(n6114), .ip2(n6113), .op(n6116) );
  nand2_1 U6270 ( .ip1(n9024), .ip2(n9023), .op(n9026) );
  inv_1 U6271 ( .ip(n8154), .op(n8144) );
  nand2_1 U6272 ( .ip1(n8031), .ip2(n8030), .op(n8147) );
  mux2_1 U6273 ( .ip1(i_i2c_ic_fs_lcnt[5]), .ip2(i_i2c_ic_lcnt[5]), .s(n6717), 
        .op(n7940) );
  nor2_1 U6274 ( .ip1(n7104), .ip2(n7103), .op(n7255) );
  mux2_1 U6275 ( .ip1(i_i2c_ic_fs_lcnt[7]), .ip2(i_i2c_ic_lcnt[7]), .s(n6717), 
        .op(n7939) );
  mux2_1 U6276 ( .ip1(i_i2c_ic_fs_lcnt[4]), .ip2(i_i2c_ic_lcnt[4]), .s(n6717), 
        .op(n7958) );
  xnor2_1 U6277 ( .ip1(n7938), .ip2(n6759), .op(n9013) );
  inv_1 U6278 ( .ip(n7255), .op(n7264) );
  nand2_1 U6279 ( .ip1(n8917), .ip2(n8901), .op(n8906) );
  xnor2_1 U6280 ( .ip1(n7934), .ip2(n6731), .op(n8967) );
  nand2_1 U6281 ( .ip1(n6764), .ip2(n6730), .op(n6731) );
  inv_1 U6282 ( .ip(n9018), .op(n8762) );
  xnor2_1 U6283 ( .ip1(n6356), .ip2(n6355), .op(n6441) );
  nor2_1 U6284 ( .ip1(n6395), .ip2(n5466), .op(n6411) );
  nand2_1 U6285 ( .ip1(n7930), .ip2(n7932), .op(n7975) );
  nand2_1 U6286 ( .ip1(n5263), .ip2(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[4]), .op(n5872) );
  xnor2_1 U6287 ( .ip1(n8065), .ip2(n6377), .op(n6378) );
  xnor2_1 U6288 ( .ip1(n8100), .ip2(n6372), .op(n6384) );
  xnor2_1 U6289 ( .ip1(n8046), .ip2(n6360), .op(n6443) );
  xnor2_1 U6290 ( .ip1(i_i2c_ic_sda_tx_hold_sync[15]), .ip2(n7143), .op(n7202)
         );
  nor2_1 U6291 ( .ip1(n7111), .ip2(n5471), .op(n7142) );
  and2_1 U6292 ( .ip1(n5700), .ip2(n6971), .op(n6029) );
  nand2_1 U6293 ( .ip1(n5548), .ip2(n10287), .op(n5570) );
  and2_1 U6294 ( .ip1(n5544), .ip2(n9058), .op(n5545) );
  and2_1 U6295 ( .ip1(n5568), .ip2(n5543), .op(n5544) );
  xnor2_1 U6296 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[14]), .ip2(i_ssi_baudr[14]), 
        .op(n10370) );
  nand3_1 U6297 ( .ip1(n10348), .ip2(n5828), .ip3(n5827), .op(n5829) );
  nand2_1 U6298 ( .ip1(n5739), .ip2(n5458), .op(n5828) );
  nor2_1 U6299 ( .ip1(n5756), .ip2(n9714), .op(n5752) );
  or2_1 U6300 ( .ip1(n6342), .ip2(n5431), .op(n6343) );
  nor2_1 U6301 ( .ip1(i_ssi_U_fifo_unconnected_rx_wrd_count[0]), .ip2(n10219), 
        .op(n10220) );
  nor2_1 U6302 ( .ip1(n5904), .ip2(n6040), .op(n5916) );
  nor2_1 U6303 ( .ip1(n10246), .ip2(n6040), .op(n5990) );
  nand2_1 U6304 ( .ip1(n5642), .ip2(n6979), .op(n6985) );
  inv_1 U6305 ( .ip(n6841), .op(n8294) );
  nor2_1 U6306 ( .ip1(n8266), .ip2(n10582), .op(n8339) );
  inv_1 U6307 ( .ip(n9969), .op(n11513) );
  inv_1 U6308 ( .ip(i_ssi_cfs[2]), .op(n9960) );
  nand2_1 U6309 ( .ip1(n9358), .ip2(i_apb_hready_resp), .op(n6554) );
  nor2_1 U6310 ( .ip1(n10341), .ip2(n10340), .op(n10345) );
  and2_1 U6311 ( .ip1(n5739), .ip2(n10343), .op(n10344) );
  nand2_1 U6312 ( .ip1(n6603), .ip2(n11569), .op(n11227) );
  nand2_1 U6313 ( .ip1(n6602), .ip2(n6601), .op(n6603) );
  inv_1 U6314 ( .ip(n8339), .op(n9699) );
  nor2_1 U6315 ( .ip1(n9725), .ip2(n9699), .op(n9153) );
  nand2_1 U6316 ( .ip1(n11283), .ip2(n9096), .op(n6841) );
  or2_1 U6317 ( .ip1(n8335), .ip2(n6631), .op(n6843) );
  nor2_1 U6318 ( .ip1(n6956), .ip2(n6955), .op(n6957) );
  nor2_1 U6319 ( .ip1(n7740), .ip2(n6954), .op(n6955) );
  nor3_1 U6320 ( .ip1(n11304), .ip2(n6952), .ip3(n7760), .op(n6953) );
  nor2_1 U6321 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_N487), .ip2(n6474), .op(n9727)
         );
  nand2_1 U6322 ( .ip1(n9921), .ip2(n9920), .op(n9922) );
  mux2_1 U6323 ( .ip1(n11522), .ip2(n9680), .s(n11529), .op(n9678) );
  nand2_1 U6324 ( .ip1(n9975), .ip2(n9974), .op(n11512) );
  nor2_1 U6325 ( .ip1(n10545), .ip2(n11581), .op(n9974) );
  inv_1 U6326 ( .ip(n9973), .op(n9975) );
  nand2_1 U6327 ( .ip1(n9946), .ip2(n7090), .op(n9970) );
  mux2_1 U6328 ( .ip1(n9969), .ip2(n9973), .s(n11581), .op(n7090) );
  nand2_1 U6329 ( .ip1(n9838), .ip2(n11598), .op(n7087) );
  or2_1 U6330 ( .ip1(n8994), .ip2(n8993), .op(n8995) );
  nor2_1 U6331 ( .ip1(n8992), .ip2(n8991), .op(n8993) );
  nor2_1 U6332 ( .ip1(n8987), .ip2(n10968), .op(n8994) );
  and2_1 U6333 ( .ip1(n8988), .ip2(n10964), .op(n8992) );
  nand2_1 U6334 ( .ip1(n8987), .ip2(n10968), .op(n8996) );
  nand2_1 U6335 ( .ip1(n8983), .ip2(n8982), .op(n9003) );
  mux2_1 U6336 ( .ip1(i_i2c_ic_fs_spklen[4]), .ip2(i_i2c_ic_hs_spklen[4]), .s(
        n7672), .op(n7164) );
  nor2_1 U6337 ( .ip1(n8040), .ip2(n8095), .op(n8058) );
  nand2_1 U6338 ( .ip1(n8079), .ip2(n8100), .op(n8040) );
  mux2_1 U6339 ( .ip1(n7318), .ip2(i_i2c_ic_sda_tx_hold_sync[1]), .s(n7321), 
        .op(n7324) );
  xnor2_1 U6340 ( .ip1(i_i2c_ic_sda_tx_hold_sync[2]), .ip2(n7122), .op(n7123)
         );
  mux2_1 U6341 ( .ip1(i_i2c_ic_fs_spklen[7]), .ip2(i_i2c_ic_hs_spklen[7]), .s(
        n7672), .op(n7182) );
  inv_1 U6342 ( .ip(n7182), .op(n7185) );
  nor2_1 U6343 ( .ip1(n9007), .ip2(n9006), .op(n9008) );
  nand2_1 U6344 ( .ip1(n8986), .ip2(n8985), .op(n9007) );
  and2_1 U6345 ( .ip1(n9005), .ip2(n9004), .op(n9006) );
  nor2_1 U6346 ( .ip1(n5464), .ip2(n8979), .op(n8986) );
  inv_1 U6347 ( .ip(n8065), .op(n8091) );
  mux2_1 U6348 ( .ip1(n7303), .ip2(i_i2c_ic_sda_tx_hold_sync[3]), .s(n7321), 
        .op(n7831) );
  nor2_1 U6349 ( .ip1(n7123), .ip2(n9773), .op(n7305) );
  nor2_1 U6350 ( .ip1(n7134), .ip2(n7133), .op(n7308) );
  inv_1 U6351 ( .ip(n7314), .op(n7134) );
  nor2_1 U6352 ( .ip1(n7313), .ip2(n7316), .op(n7133) );
  mux2_1 U6353 ( .ip1(i_i2c_ic_fs_lcnt[3]), .ip2(i_i2c_ic_lcnt[3]), .s(n6717), 
        .op(n7941) );
  mux2_1 U6354 ( .ip1(i_i2c_ic_fs_lcnt[2]), .ip2(i_i2c_ic_lcnt[2]), .s(n6717), 
        .op(n7949) );
  nor2_2 U6355 ( .ip1(n8010), .ip2(n8009), .op(n8162) );
  nor2_1 U6356 ( .ip1(n8135), .ip2(n8134), .op(n8138) );
  nor2_1 U6357 ( .ip1(n8144), .ip2(n5452), .op(n8134) );
  nand2_1 U6358 ( .ip1(n8080), .ip2(n8093), .op(n8081) );
  nand2_1 U6359 ( .ip1(n8097), .ip2(n8082), .op(n8080) );
  inv_1 U6360 ( .ip(n7274), .op(n7282) );
  xnor2_1 U6361 ( .ip1(i_i2c_ic_sda_tx_hold_sync[5]), .ip2(n7107), .op(n7113)
         );
  xnor2_1 U6362 ( .ip1(i_i2c_ic_sda_tx_hold_sync[6]), .ip2(n7106), .op(n7109)
         );
  or2_1 U6363 ( .ip1(i_i2c_ic_sda_tx_hold_sync[5]), .ip2(n7107), .op(n7108) );
  inv_1 U6364 ( .ip(n7263), .op(n7254) );
  nor2_1 U6365 ( .ip1(n7113), .ip2(n7112), .op(n7274) );
  nor2_1 U6366 ( .ip1(n7109), .ip2(n7108), .op(n7271) );
  nor2_1 U6367 ( .ip1(n8133), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[7]), 
        .op(n8142) );
  and2_1 U6368 ( .ip1(n10741), .ip2(n10742), .op(n10739) );
  nor2_1 U6369 ( .ip1(n8133), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[7]), .op(n8687) );
  nand2_1 U6370 ( .ip1(n6810), .ip2(n6809), .op(n6812) );
  or2_1 U6371 ( .ip1(n6808), .ip2(n6807), .op(n6809) );
  nand2_1 U6372 ( .ip1(n6794), .ip2(n6793), .op(n6817) );
  xnor2_1 U6373 ( .ip1(n7939), .ip2(n6768), .op(n9018) );
  nand2_1 U6374 ( .ip1(n7113), .ip2(n7112), .op(n7281) );
  inv_1 U6375 ( .ip(n7271), .op(n7273) );
  nand2_1 U6376 ( .ip1(n7109), .ip2(n7108), .op(n7272) );
  inv_1 U6377 ( .ip(n7105), .op(n7251) );
  nand2_1 U6378 ( .ip1(n7225), .ip2(n7243), .op(n7226) );
  nor2_1 U6379 ( .ip1(n7230), .ip2(n7224), .op(n7225) );
  xnor2_1 U6380 ( .ip1(i_i2c_ic_sda_tx_hold_sync[10]), .ip2(n7234), .op(n7235)
         );
  nor2_1 U6381 ( .ip1(n7232), .ip2(n5471), .op(n7233) );
  inv_1 U6382 ( .ip(n7250), .op(n7230) );
  nand2_1 U6383 ( .ip1(n8943), .ip2(n8942), .op(n8947) );
  nor2_1 U6384 ( .ip1(n8886), .ip2(n8885), .op(n8909) );
  nor2_1 U6385 ( .ip1(n8881), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[14]), .op(n8886) );
  nor2_1 U6386 ( .ip1(n8903), .ip2(n8896), .op(n8917) );
  nor2_1 U6387 ( .ip1(n7965), .ip2(n7939), .op(n6716) );
  nor2_1 U6388 ( .ip1(n7977), .ip2(n7925), .op(n6728) );
  nand2_1 U6389 ( .ip1(n7971), .ip2(n7970), .op(n7986) );
  nand2_1 U6390 ( .ip1(n8629), .ip2(n8628), .op(n8633) );
  or2_1 U6391 ( .ip1(n8627), .ip2(n8626), .op(n8628) );
  nand2_1 U6392 ( .ip1(n8619), .ip2(n8618), .op(n8620) );
  nor2_1 U6393 ( .ip1(n8616), .ip2(n8615), .op(n8638) );
  nand2_1 U6394 ( .ip1(n8780), .ip2(n8779), .op(n8785) );
  or2_1 U6395 ( .ip1(n8778), .ip2(n8777), .op(n8779) );
  nand2_1 U6396 ( .ip1(n8770), .ip2(n8769), .op(n8771) );
  nor2_1 U6397 ( .ip1(n8767), .ip2(n8766), .op(n8790) );
  nand2_1 U6398 ( .ip1(n6268), .ip2(n6267), .op(n6270) );
  nor2_1 U6399 ( .ip1(n6224), .ip2(i_ssi_baudr[12]), .op(n6268) );
  inv_1 U6400 ( .ip(n9088), .op(n6261) );
  nor2_1 U6401 ( .ip1(n5564), .ip2(n5563), .op(n5628) );
  nand2_1 U6402 ( .ip1(n6297), .ip2(n5562), .op(n5564) );
  nor2_1 U6403 ( .ip1(n5653), .ip2(n5652), .op(n5654) );
  nor2_1 U6404 ( .ip1(n9059), .ip2(n5594), .op(n5653) );
  inv_1 U6405 ( .ip(n5261), .op(n6081) );
  xnor2_1 U6406 ( .ip1(n8021), .ip2(n6414), .op(n6415) );
  xnor2_1 U6407 ( .ip1(n8023), .ip2(n6418), .op(n6422) );
  mux2_1 U6408 ( .ip1(n7270), .ip2(i_i2c_ic_sda_tx_hold_sync[7]), .s(n7321), 
        .op(n7343) );
  xnor2_1 U6409 ( .ip1(n7269), .ip2(n7268), .op(n7270) );
  nand2_1 U6410 ( .ip1(n7264), .ip2(n7263), .op(n7269) );
  mux2_1 U6411 ( .ip1(n7261), .ip2(i_i2c_ic_sda_tx_hold_sync[8]), .s(n7321), 
        .op(n7880) );
  xnor2_1 U6412 ( .ip1(n7260), .ip2(n7259), .op(n7261) );
  nand2_1 U6413 ( .ip1(n7251), .ip2(n7250), .op(n7260) );
  nand2_1 U6414 ( .ip1(n7258), .ip2(n7257), .op(n7259) );
  or4_1 U6415 ( .ip1(i_i2c_ic_sda_tx_hold_sync[13]), .ip2(
        i_i2c_ic_sda_tx_hold_sync[12]), .ip3(i_i2c_ic_sda_tx_hold_sync[11]), 
        .ip4(i_i2c_ic_sda_tx_hold_sync[10]), .op(n7124) );
  xnor2_1 U6416 ( .ip1(i_i2c_ic_sda_tx_hold_sync[9]), .ip2(n7247), .op(n7249)
         );
  nor2_1 U6417 ( .ip1(n7244), .ip2(n5471), .op(n7246) );
  nand2_1 U6418 ( .ip1(n7212), .ip2(n7243), .op(n7213) );
  nor2_1 U6419 ( .ip1(n7230), .ip2(n7211), .op(n7212) );
  nand2_1 U6420 ( .ip1(n7219), .ip2(n7243), .op(n7220) );
  nor2_1 U6421 ( .ip1(n7230), .ip2(n7218), .op(n7219) );
  inv_1 U6422 ( .ip(n7217), .op(n7218) );
  and2_1 U6423 ( .ip1(n10735), .ip2(n10736), .op(n10768) );
  nand2_1 U6424 ( .ip1(n10700), .ip2(n10699), .op(n10769) );
  nand4_1 U6425 ( .ip1(n6522), .ip2(n7668), .ip3(n7664), .ip4(n7654), .op(
        n6523) );
  nor2_1 U6426 ( .ip1(n8602), .ip2(n8601), .op(n8603) );
  nand2_1 U6427 ( .ip1(n8584), .ip2(n8583), .op(n8585) );
  nand2_1 U6428 ( .ip1(n6694), .ip2(n6631), .op(n6635) );
  nor2_1 U6429 ( .ip1(n6701), .ip2(n6700), .op(n6931) );
  mux2_1 U6430 ( .ip1(i_i2c_tx_fifo_data_buf[8]), .ip2(n9096), .s(
        i_i2c_U_DW_apb_i2c_mstfsm_old_is_read), .op(n6927) );
  and2_1 U6431 ( .ip1(n10772), .ip2(n10773), .op(n10709) );
  nand2_1 U6432 ( .ip1(n10708), .ip2(n10707), .op(n10710) );
  nor2_1 U6433 ( .ip1(i_ssi_U_mstfsm_bit_cnt[4]), .ip2(n5665), .op(n5669) );
  nand2_1 U6434 ( .ip1(n5610), .ip2(n9850), .op(n5596) );
  nor2_1 U6435 ( .ip1(n6215), .ip2(n6224), .op(n6218) );
  inv_1 U6436 ( .ip(n6267), .op(n6215) );
  inv_1 U6437 ( .ip(n6216), .op(n6217) );
  nor2_1 U6438 ( .ip1(n6253), .ip2(n10310), .op(n6241) );
  inv_1 U6439 ( .ip(n5449), .op(n6246) );
  xnor2_1 U6440 ( .ip1(n10433), .ip2(n6243), .op(n5449) );
  nor3_1 U6441 ( .ip1(n5635), .ip2(n5634), .ip3(n5633), .op(n5637) );
  nand2_1 U6442 ( .ip1(n6489), .ip2(n6488), .op(n7644) );
  nor2_1 U6443 ( .ip1(n9059), .ip2(i_ssi_U_mstfsm_c_state[1]), .op(n5607) );
  nor2_1 U6444 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[7]), 
        .ip2(n6507), .op(n6331) );
  nor2_1 U6445 ( .ip1(n7901), .ip2(n7900), .op(n7904) );
  nand2_1 U6446 ( .ip1(n7891), .ip2(n7890), .op(n7901) );
  nor2_1 U6447 ( .ip1(n7902), .ip2(n7875), .op(n7906) );
  xnor2_1 U6448 ( .ip1(i_i2c_ic_sda_tx_hold_sync[14]), .ip2(n7209), .op(n7210)
         );
  nor2_1 U6449 ( .ip1(n7207), .ip2(n5471), .op(n7208) );
  nor2_1 U6450 ( .ip1(n7887), .ip2(n11094), .op(n7888) );
  nor2_1 U6451 ( .ip1(n7931), .ip2(n7975), .op(n8001) );
  nand2_1 U6452 ( .ip1(n7034), .ip2(n7033), .op(n7039) );
  nand2_1 U6453 ( .ip1(n10894), .ip2(n10774), .op(n10787) );
  nor3_1 U6454 ( .ip1(n10765), .ip2(n10870), .ip3(n10763), .op(n10767) );
  inv_1 U6455 ( .ip(n7031), .op(n7044) );
  or4_1 U6456 ( .ip1(n6708), .ip2(n6707), .ip3(n6706), .ip4(n6705), .op(n6709)
         );
  nor3_1 U6457 ( .ip1(n6699), .ip2(n9666), .ip3(n10582), .op(n6706) );
  nor2_1 U6458 ( .ip1(n6616), .ip2(n6470), .op(n6708) );
  nor2_1 U6459 ( .ip1(n11578), .ip2(n11579), .op(n11580) );
  mux2_1 U6460 ( .ip1(n11577), .ip2(i_ssi_fsm_busy), .s(n11576), .op(n11578)
         );
  or2_1 U6461 ( .ip1(n11581), .ip2(n11580), .op(n11582) );
  inv_1 U6462 ( .ip(n6114), .op(n5382) );
  nand2_1 U6463 ( .ip1(n11217), .ip2(n9698), .op(n10166) );
  inv_1 U6464 ( .ip(n6231), .op(n6234) );
  xor2_1 U6465 ( .ip1(n10461), .ip2(i_ssi_baudr[12]), .op(n6216) );
  inv_1 U6466 ( .ip(n11235), .op(n11236) );
  nand2_1 U6467 ( .ip1(n11239), .ip2(n11235), .op(n11233) );
  nor2_1 U6468 ( .ip1(n6610), .ip2(n10223), .op(n10219) );
  nor2_1 U6469 ( .ip1(n6678), .ip2(n6674), .op(n6662) );
  nor2_1 U6470 ( .ip1(n6850), .ip2(n6965), .op(n6860) );
  xor2_1 U6471 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[4]), 
        .ip2(i_i2c_ic_hs_spklen[4]), .op(n6335) );
  nand2_1 U6472 ( .ip1(n7388), .ip2(n7393), .op(n6320) );
  xor2_1 U6473 ( .ip1(i_i2c_ic_fs_spklen[7]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[7]), .op(n6324) );
  nor2_1 U6474 ( .ip1(n6323), .ip2(n6322), .op(n7398) );
  nor2_1 U6475 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[3]), 
        .ip2(n6321), .op(n6322) );
  nor2_1 U6476 ( .ip1(i_i2c_ic_hs_spklen[1]), .ip2(n7362), .op(n6329) );
  nor2_1 U6477 ( .ip1(n10250), .ip2(n6040), .op(n6041) );
  mux2_1 U6478 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_buffer[3]), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[15]), .s(n6143), .op(n6070) );
  nand2_1 U6479 ( .ip1(n6090), .ip2(n6089), .op(n6091) );
  nor2_1 U6480 ( .ip1(n6088), .ip2(n6087), .op(n6090) );
  nand2_1 U6481 ( .ip1(n10490), .ip2(n10489), .op(n10502) );
  mux2_1 U6482 ( .ip1(n11547), .ip2(n9366), .s(n6290), .op(n10490) );
  nor2_1 U6483 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[15]), .ip2(
        n7203), .op(n10423) );
  nor2_1 U6484 ( .ip1(n7354), .ip2(n11102), .op(n10427) );
  nor2_1 U6485 ( .ip1(n7863), .ip2(n7862), .op(n10425) );
  inv_1 U6486 ( .ip(n8535), .op(n8551) );
  nor2_1 U6487 ( .ip1(n7422), .ip2(n8286), .op(n8296) );
  nand2_1 U6488 ( .ip1(n8527), .ip2(n11302), .op(n8535) );
  nand2_1 U6489 ( .ip1(n7422), .ip2(n7921), .op(n8525) );
  mux2_1 U6490 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_data_d_int_0_), 
        .ip2(n6534), .s(n6533), .op(n7048) );
  nand2_1 U6491 ( .ip1(n6532), .ip2(n9404), .op(n6533) );
  nand2_1 U6492 ( .ip1(n6528), .ip2(n6527), .op(n6532) );
  inv_1 U6493 ( .ip(n6694), .op(n8335) );
  nand3_1 U6494 ( .ip1(n9662), .ip2(n9664), .ip3(n8334), .op(n6643) );
  nand2_1 U6495 ( .ip1(n10413), .ip2(n8335), .op(n6845) );
  or4_1 U6496 ( .ip1(n6639), .ip2(n6638), .ip3(n8332), .ip4(n6637), .op(n6640)
         );
  nor3_1 U6497 ( .ip1(n9429), .ip2(n6933), .ip3(n6932), .op(n6943) );
  nand4_1 U6498 ( .ip1(n6894), .ip2(n6893), .ip3(n6892), .ip4(n6891), .op(
        n6895) );
  inv_1 U6499 ( .ip(n8217), .op(n6900) );
  nand2_1 U6500 ( .ip1(n9449), .ip2(n6922), .op(n6945) );
  nor2_1 U6501 ( .ip1(n6920), .ip2(n6919), .op(n6951) );
  nand4_1 U6502 ( .ip1(n9402), .ip2(n6918), .ip3(n6917), .ip4(n6916), .op(
        n6919) );
  nand2_1 U6503 ( .ip1(n6622), .ip2(n6621), .op(n6715) );
  nand3_1 U6504 ( .ip1(n6912), .ip2(n6908), .ip3(n6620), .op(n6622) );
  nor2_1 U6505 ( .ip1(n5749), .ip2(n5696), .op(n5697) );
  nor2_1 U6506 ( .ip1(n5695), .ip2(n5751), .op(n5696) );
  nand2_1 U6507 ( .ip1(n7626), .ip2(n5647), .op(n5537) );
  nor2_1 U6508 ( .ip1(n5542), .ip2(n5601), .op(n5550) );
  inv_1 U6509 ( .ip(n6140), .op(n5549) );
  inv_1 U6510 ( .ip(i_ssi_baudr[14]), .op(n7583) );
  nor2_1 U6511 ( .ip1(n9908), .ip2(n9786), .op(n11692) );
  nor2_1 U6512 ( .ip1(n9908), .ip2(n7802), .op(n11693) );
  inv_1 U6513 ( .ip(n9899), .op(n7500) );
  mux2_1 U6514 ( .ip1(ex_i_ahb_AHB_Slave_RAM_hready_resp), .ip2(n6549), .s(
        n9195), .op(n6550) );
  nor4_1 U6515 ( .ip1(n10322), .ip2(n10321), .ip3(n10320), .ip4(n10319), .op(
        n10327) );
  mux2_1 U6516 ( .ip1(i_i2c_prdata[0]), .ip2(i_ssi_prdata[0]), .s(n9335), .op(
        n9280) );
  mux2_1 U6517 ( .ip1(i_i2c_prdata[1]), .ip2(i_ssi_prdata[1]), .s(n9335), .op(
        n9270) );
  mux2_1 U6518 ( .ip1(i_i2c_prdata[2]), .ip2(i_ssi_prdata[2]), .s(n9335), .op(
        n9225) );
  mux2_1 U6519 ( .ip1(i_i2c_prdata[3]), .ip2(i_ssi_prdata[3]), .s(n9335), .op(
        n9260) );
  mux2_1 U6520 ( .ip1(i_i2c_prdata[7]), .ip2(i_ssi_prdata[7]), .s(n9335), .op(
        n9295) );
  mux2_1 U6521 ( .ip1(i_i2c_prdata[17]), .ip2(i_ssi_prdata[17]), .s(n9335), 
        .op(n9265) );
  mux2_1 U6522 ( .ip1(i_i2c_prdata[19]), .ip2(i_ssi_prdata[19]), .s(n9335), 
        .op(n9310) );
  mux2_1 U6523 ( .ip1(i_i2c_prdata[20]), .ip2(i_ssi_prdata[20]), .s(n9335), 
        .op(n9210) );
  mux2_1 U6524 ( .ip1(i_i2c_prdata[22]), .ip2(i_ssi_prdata[22]), .s(n9335), 
        .op(n9336) );
  nor2_1 U6525 ( .ip1(n10244), .ip2(n6547), .op(n10270) );
  inv_1 U6526 ( .ip(n6250), .op(n6251) );
  nand2_1 U6527 ( .ip1(n10352), .ip2(n10351), .op(n10356) );
  nand2_1 U6528 ( .ip1(n5833), .ip2(n5359), .op(n5834) );
  nand2_1 U6529 ( .ip1(n5848), .ip2(n5389), .op(n5856) );
  nand2_1 U6530 ( .ip1(n5854), .ip2(n5853), .op(n5855) );
  nand2_1 U6531 ( .ip1(n10188), .ip2(n10187), .op(n10189) );
  mux2_1 U6532 ( .ip1(i_ssi_U_fifo_unconnected_rx_wrd_count[2]), .ip2(n6614), 
        .s(n6613), .op(n11244) );
  nand2_1 U6533 ( .ip1(i_i2c_fifo_rst_n), .ip2(n11192), .op(n11198) );
  nand2_1 U6534 ( .ip1(i_i2c_fifo_rst_n), .ip2(n11184), .op(n11201) );
  nand2_1 U6535 ( .ip1(n10240), .ip2(n8375), .op(n5680) );
  inv_1 U6536 ( .ip(n5233), .op(n5682) );
  nand2_1 U6537 ( .ip1(n6651), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[1]), .op(n9942) );
  nand2_1 U6538 ( .ip1(n6455), .ip2(n6454), .op(n6456) );
  nor2_1 U6539 ( .ip1(n6388), .ip2(n6387), .op(n6389) );
  nor2_1 U6540 ( .ip1(n7068), .ip2(n11167), .op(n8569) );
  nand2_1 U6541 ( .ip1(n10528), .ip2(i_ssi_U_mstfsm_frame_cnt[10]), .op(n10532) );
  nor2_2 U6542 ( .ip1(n10532), .ip2(n10533), .op(n10536) );
  nor2_1 U6543 ( .ip1(n7916), .ip2(n11099), .op(n7913) );
  nand2_1 U6544 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[0]), .ip2(
        n11056), .op(n11057) );
  nor2_1 U6545 ( .ip1(n9096), .ip2(n6947), .op(n9661) );
  inv_1 U6546 ( .ip(n6901), .op(n9735) );
  nor2_1 U6547 ( .ip1(i_i2c_mst_debug_cstate[1]), .ip2(n6926), .op(n9448) );
  inv_1 U6548 ( .ip(n9410), .op(n9667) );
  nand2_1 U6549 ( .ip1(n6694), .ip2(n8336), .op(n9737) );
  nand2_1 U6550 ( .ip1(n10951), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[13]), .op(n10957) );
  inv_1 U6551 ( .ip(n11284), .op(n6482) );
  nor2_1 U6552 ( .ip1(n7921), .ip2(n7634), .op(n8259) );
  nor2_1 U6553 ( .ip1(n11146), .ip2(n11147), .op(n11145) );
  nor3_1 U6554 ( .ip1(n7046), .ip2(n7045), .ip3(n9752), .op(n7047) );
  nor3_1 U6555 ( .ip1(n7043), .ip2(n9757), .ip3(n9753), .op(n7045) );
  inv_1 U6556 ( .ip(n11133), .op(n7505) );
  nand2_1 U6557 ( .ip1(n8339), .ip2(n8338), .op(n8342) );
  or3_1 U6558 ( .ip1(n8337), .ip2(n11051), .ip3(n9409), .op(n8338) );
  inv_1 U6559 ( .ip(n11047), .op(n7760) );
  mux2_1 U6560 ( .ip1(n11047), .ip2(n11045), .s(n11044), .op(n11304) );
  nor2_1 U6561 ( .ip1(n6715), .ip2(n6952), .op(n11305) );
  nand2_1 U6562 ( .ip1(n10722), .ip2(n10721), .op(n10726) );
  and2_1 U6563 ( .ip1(n10724), .ip2(n10723), .op(n10725) );
  inv_1 U6564 ( .ip(n10835), .op(n10910) );
  inv_1 U6565 ( .ip(n6899), .op(n6479) );
  inv_1 U6566 ( .ip(i_i2c_U_DW_apb_i2c_mstfsm_N487), .op(n11053) );
  nor3_1 U6567 ( .ip1(n11613), .ip2(n11612), .ip3(n11611), .op(n11622) );
  nor2_1 U6568 ( .ip1(i_ssi_ssi_txo_intr_n), .ip2(n11562), .op(n11613) );
  nand4_1 U6569 ( .ip1(n11604), .ip2(n11603), .ip3(n11602), .ip4(n11601), .op(
        n11612) );
  xnor2_1 U6570 ( .ip1(n8376), .ip2(n8375), .op(n9920) );
  nand3_1 U6571 ( .ip1(n5475), .ip2(n6141), .ip3(n6140), .op(n6142) );
  nor2_1 U6572 ( .ip1(n11531), .ip2(n11529), .op(n9676) );
  nand2_1 U6573 ( .ip1(n9670), .ip2(n9669), .op(n9671) );
  nand2_1 U6574 ( .ip1(n9685), .ip2(n5594), .op(n9689) );
  inv_1 U6575 ( .ip(n11702), .op(n5726) );
  nand2_1 U6576 ( .ip1(n5725), .ip2(n10486), .op(n5727) );
  or2_1 U6577 ( .ip1(n5689), .ip2(n5723), .op(n5725) );
  nor2_1 U6578 ( .ip1(n5720), .ip2(n5719), .op(n9708) );
  nor2_1 U6579 ( .ip1(n6980), .ip2(n5756), .op(n5720) );
  nand2_1 U6580 ( .ip1(n5718), .ip2(n5749), .op(n5719) );
  nand2_1 U6581 ( .ip1(n5717), .ip2(n5716), .op(n5718) );
  nor2_1 U6582 ( .ip1(n5779), .ip2(n5778), .op(n6101) );
  nand4_1 U6583 ( .ip1(n5949), .ip2(n5948), .ip3(n5947), .ip4(n5946), .op(
        n5950) );
  nor2_1 U6584 ( .ip1(n5979), .ip2(n5978), .op(n10248) );
  or2_1 U6585 ( .ip1(n11515), .ip2(n11514), .op(n11516) );
  nor3_1 U6586 ( .ip1(n9972), .ip2(n9971), .ip3(n9970), .op(n11519) );
  nor2_1 U6587 ( .ip1(n10545), .ip2(n9969), .op(n9972) );
  nand2_1 U6588 ( .ip1(n11513), .ip2(n7089), .op(n9976) );
  nand2_1 U6589 ( .ip1(n7084), .ip2(n7083), .op(n9973) );
  nand2_1 U6590 ( .ip1(n5482), .ip2(i_ssi_U_mstfsm_last_frame), .op(n5535) );
  nand2_1 U6591 ( .ip1(n5441), .ip2(n9963), .op(n9964) );
  xnor2_1 U6592 ( .ip1(n9960), .ip2(n11706), .op(n5441) );
  nor2_1 U6593 ( .ip1(n9962), .ip2(n9961), .op(n9963) );
  mux2_1 U6594 ( .ip1(i_ssi_U_mstfsm_ctrl_cnt[1]), .ip2(n11704), .s(
        i_ssi_cfs[1]), .op(n9965) );
  inv_1 U6595 ( .ip(n7628), .op(n9984) );
  nand2_1 U6596 ( .ip1(n10404), .ip2(n10403), .op(n10405) );
  nand2_1 U6597 ( .ip1(n7520), .ip2(n7519), .op(n11624) );
  and3_1 U6598 ( .ip1(n10107), .ip2(n6584), .ip3(n10008), .op(n6585) );
  nand2_1 U6599 ( .ip1(n5421), .ip2(n5474), .op(n9383) );
  nand2_1 U6600 ( .ip1(n9376), .ip2(n9375), .op(n9391) );
  nand3_1 U6601 ( .ip1(n10300), .ip2(n11569), .ip3(n10299), .op(n10301) );
  inv_1 U6602 ( .ip(n10579), .op(i_i2c_sda_int) );
  nand2_1 U6603 ( .ip1(n6993), .ip2(n6992), .op(n6994) );
  mux2_1 U6604 ( .ip1(i_ssi_imr[5]), .ip2(i_apb_pwdata_int[5]), .s(n9917), 
        .op(n4645) );
  mux2_1 U6605 ( .ip1(i_apb_hready_resp), .ip2(n10030), .s(n10029), .op(n4824)
         );
  nor2_1 U6606 ( .ip1(n6960), .ip2(n6959), .op(n5117) );
  nor2_1 U6607 ( .ip1(n6958), .ip2(n6957), .op(n6959) );
  nor2_1 U6608 ( .ip1(n5232), .ip2(n8442), .op(n6958) );
  nand2_1 U6609 ( .ip1(n6578), .ip2(n9377), .op(n6579) );
  nand2_1 U6610 ( .ip1(n10018), .ip2(n9377), .op(n6580) );
  nor2_1 U6611 ( .ip1(n8990), .ip2(n8989), .op(n8991) );
  nand2_1 U6612 ( .ip1(n7944), .ip2(n10959), .op(n8989) );
  nor2_1 U6613 ( .ip1(n8988), .ip2(n10964), .op(n8990) );
  mux2_1 U6614 ( .ip1(i_i2c_ic_fs_spklen[3]), .ip2(i_i2c_ic_hs_spklen[3]), .s(
        n7672), .op(n7145) );
  mux2_1 U6615 ( .ip1(i_i2c_ic_fs_spklen[5]), .ip2(i_i2c_ic_hs_spklen[5]), .s(
        n7672), .op(n7147) );
  nor2_1 U6616 ( .ip1(n9003), .ip2(n9002), .op(n9004) );
  nand2_1 U6617 ( .ip1(n9000), .ip2(n8999), .op(n9005) );
  nand2_1 U6618 ( .ip1(n8998), .ip2(n8997), .op(n8999) );
  nand2_1 U6619 ( .ip1(n8996), .ip2(n8995), .op(n8998) );
  nor2_1 U6620 ( .ip1(n9022), .ip2(n9021), .op(n9019) );
  nand2_1 U6621 ( .ip1(n7323), .ip2(n7358), .op(n7326) );
  mux2_1 U6622 ( .ip1(n7322), .ip2(i_i2c_ic_sda_tx_hold_sync[0]), .s(n7321), 
        .op(n7323) );
  nand2_1 U6623 ( .ip1(n7131), .ip2(i_i2c_ic_sda_tx_hold_sync[1]), .op(n7314)
         );
  inv_1 U6624 ( .ip(n7147), .op(n7150) );
  nor2_1 U6625 ( .ip1(n7171), .ip2(n7170), .op(n7172) );
  inv_1 U6626 ( .ip(n7169), .op(n7171) );
  xnor2_1 U6627 ( .ip1(i_i2c_ic_fs_spklen[1]), .ip2(i_i2c_ic_fs_spklen[2]), 
        .op(n8011) );
  mux2_1 U6628 ( .ip1(n7311), .ip2(i_i2c_ic_sda_tx_hold_sync[2]), .s(n7321), 
        .op(n7832) );
  xnor2_1 U6629 ( .ip1(i_i2c_ic_sda_tx_hold_sync[4]), .ip2(n7115), .op(n7120)
         );
  xnor2_1 U6630 ( .ip1(i_i2c_ic_sda_tx_hold_sync[3]), .ip2(n7116), .op(n7137)
         );
  nor2_1 U6631 ( .ip1(n7137), .ip2(n7136), .op(n7291) );
  nand2_1 U6632 ( .ip1(n7185), .ip2(n7184), .op(n7189) );
  nor2_1 U6633 ( .ip1(n7177), .ip2(n7176), .op(n7178) );
  inv_1 U6634 ( .ip(n7180), .op(n7176) );
  nand3_1 U6635 ( .ip1(n9028), .ip2(n5459), .ip3(n9027), .op(n9034) );
  nand2_1 U6636 ( .ip1(n9026), .ip2(n9025), .op(n9027) );
  nor2_1 U6637 ( .ip1(n7942), .ip2(n7943), .op(n6798) );
  nand2_1 U6638 ( .ip1(n10686), .ip2(n10685), .op(n10747) );
  nand2_1 U6639 ( .ip1(i_i2c_ic_fs_lcnt[1]), .ip2(n10719), .op(n10686) );
  nand2_1 U6640 ( .ip1(i_i2c_ic_lcnt[1]), .ip2(n10720), .op(n10685) );
  nor2_1 U6641 ( .ip1(n6806), .ip2(n6805), .op(n6807) );
  nor2_1 U6642 ( .ip1(n6804), .ip2(n6803), .op(n6805) );
  xnor2_1 U6643 ( .ip1(n7943), .ip2(n7942), .op(n8988) );
  xnor2_1 U6644 ( .ip1(n7949), .ip2(n6801), .op(n8987) );
  xnor2_1 U6645 ( .ip1(n7940), .ip2(n6786), .op(n8980) );
  xnor2_1 U6646 ( .ip1(n7965), .ip2(n6783), .op(n8977) );
  nor2_1 U6647 ( .ip1(n8146), .ip2(n8145), .op(n8150) );
  nor2_1 U6648 ( .ip1(n8062), .ip2(n8061), .op(n8064) );
  nor2_1 U6649 ( .ip1(n8050), .ip2(n8049), .op(n8052) );
  nor2_1 U6650 ( .ip1(n8039), .ip2(n8038), .op(n8095) );
  inv_1 U6651 ( .ip(n8136), .op(n8024) );
  inv_1 U6652 ( .ip(n8130), .op(n8026) );
  inv_1 U6653 ( .ip(n8033), .op(n8034) );
  nand2_1 U6654 ( .ip1(n8032), .ip2(n8147), .op(n8135) );
  nand2_1 U6655 ( .ip1(n8014), .ip2(n5447), .op(n8154) );
  nand2_1 U6656 ( .ip1(n8171), .ip2(n8008), .op(n8014) );
  nor2_1 U6657 ( .ip1(n8069), .ip2(n8068), .op(n8072) );
  inv_1 U6658 ( .ip(n5596), .op(n5581) );
  and2_1 U6659 ( .ip1(i_ssi_U_mstfsm_c_state[2]), .ip2(n9057), .op(n5583) );
  and2_1 U6660 ( .ip1(n9057), .ip2(n6281), .op(n5582) );
  nor2_1 U6661 ( .ip1(n8005), .ip2(n8181), .op(n6396) );
  inv_1 U6662 ( .ip(n6396), .op(n6398) );
  xnor2_1 U6663 ( .ip1(i_i2c_ic_sda_tx_hold_sync[7]), .ip2(n7098), .op(n7104)
         );
  mux2_1 U6664 ( .ip1(n7295), .ip2(i_i2c_ic_sda_tx_hold_sync[4]), .s(n7321), 
        .op(n7837) );
  xnor2_1 U6665 ( .ip1(n7294), .ip2(n7293), .op(n7295) );
  nand2_1 U6666 ( .ip1(n7290), .ip2(n7289), .op(n7294) );
  nand2_1 U6667 ( .ip1(n7297), .ip2(n7292), .op(n7293) );
  nand2_1 U6668 ( .ip1(n7231), .ip2(n7243), .op(n7232) );
  nand2_1 U6669 ( .ip1(n7094), .ip2(n7093), .op(n7224) );
  nand2_1 U6670 ( .ip1(n7120), .ip2(n7119), .op(n7289) );
  nor2_1 U6671 ( .ip1(n7120), .ip2(n7119), .op(n7288) );
  nand2_1 U6672 ( .ip1(n7137), .ip2(n7136), .op(n7297) );
  nand2_1 U6673 ( .ip1(n7306), .ip2(n7135), .op(n7299) );
  nor2_1 U6674 ( .ip1(n7291), .ip2(n7288), .op(n7138) );
  or2_1 U6675 ( .ip1(n5470), .ip2(n8941), .op(n8942) );
  nor2_1 U6676 ( .ip1(n8880), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[15]), .op(n8885) );
  nor2_1 U6677 ( .ip1(n8887), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[13]), .op(n8907) );
  nor2_1 U6678 ( .ip1(n7958), .ip2(n7940), .op(n6782) );
  nor4_1 U6679 ( .ip1(n7948), .ip2(n7950), .ip3(n7947), .ip4(n7946), .op(n7953) );
  nor2_1 U6680 ( .ip1(n8880), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[15]), .op(n8056) );
  nor2_1 U6681 ( .ip1(n8887), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[13]), .op(n8110) );
  nand2_1 U6682 ( .ip1(i_i2c_ic_lcnt[0]), .ip2(n10720), .op(n10683) );
  nand2_1 U6683 ( .ip1(i_i2c_ic_fs_lcnt[0]), .ip2(n10719), .op(n10684) );
  and2_1 U6684 ( .ip1(n10748), .ip2(n10747), .op(n10745) );
  nand2_1 U6685 ( .ip1(n10688), .ip2(n10687), .op(n10746) );
  and2_1 U6686 ( .ip1(n10745), .ip2(n10746), .op(n10743) );
  nand2_1 U6687 ( .ip1(n10690), .ip2(n10689), .op(n10744) );
  nand2_1 U6688 ( .ip1(n10694), .ip2(n10693), .op(n10740) );
  nor2_1 U6689 ( .ip1(n8880), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[15]), .op(n8652) );
  nor2_1 U6690 ( .ip1(n8817), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[11]), .op(n8667) );
  nor2_1 U6691 ( .ip1(n8887), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[13]), .op(n8660) );
  xnor2_1 U6692 ( .ip1(n7989), .ip2(n6757), .op(n9011) );
  xnor2_1 U6693 ( .ip1(n7925), .ip2(n6733), .op(n8969) );
  nand2_1 U6694 ( .ip1(n6764), .ip2(n6732), .op(n6733) );
  inv_1 U6695 ( .ip(n8987), .op(n8781) );
  xnor2_1 U6696 ( .ip1(n7977), .ip2(n6740), .op(n8970) );
  nand2_1 U6697 ( .ip1(n6764), .ip2(n6739), .op(n6740) );
  nor2_1 U6698 ( .ip1(n8880), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[15]), .op(n8805) );
  nor2_1 U6699 ( .ip1(n8817), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[11]), .op(n8821) );
  nor2_1 U6700 ( .ip1(n8887), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[13]), .op(n8813) );
  and2_1 U6701 ( .ip1(i_ssi_U_mstfsm_ss_in_n_sync), .ip2(i_ssi_sclk_re), .op(
        n5649) );
  and3_1 U6702 ( .ip1(n5575), .ip2(n5574), .ip3(n5689), .op(n5410) );
  inv_1 U6703 ( .ip(n6393), .op(n6394) );
  xnor2_1 U6704 ( .ip1(n8031), .ip2(n6392), .op(n6393) );
  xnor2_1 U6705 ( .ip1(n6397), .ip2(n8010), .op(n5430) );
  nor2_1 U6706 ( .ip1(n6398), .ip2(n8012), .op(n6397) );
  and2_1 U6707 ( .ip1(n6402), .ip2(n6404), .op(n6401) );
  nor2_1 U6708 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[3]), .ip2(n5430), .op(n6403) );
  xnor2_1 U6709 ( .ip1(n8012), .ip2(n6398), .op(n6402) );
  inv_1 U6710 ( .ip(n7252), .op(n7267) );
  nand2_1 U6711 ( .ip1(n7104), .ip2(n7103), .op(n7263) );
  mux2_1 U6712 ( .ip1(n7286), .ip2(i_i2c_ic_sda_tx_hold_sync[5]), .s(n7321), 
        .op(n7830) );
  inv_1 U6713 ( .ip(n7285), .op(n7286) );
  xnor2_1 U6714 ( .ip1(n7284), .ip2(n7283), .op(n7285) );
  nand2_1 U6715 ( .ip1(n7282), .ip2(n7281), .op(n7283) );
  nor2_1 U6716 ( .ip1(n7846), .ip2(n7845), .op(n7847) );
  and2_1 U6717 ( .ip1(n7844), .ip2(n7843), .op(n7845) );
  nor2_1 U6718 ( .ip1(n7840), .ip2(n7839), .op(n7846) );
  nand2_1 U6719 ( .ip1(n7265), .ip2(n7264), .op(n7256) );
  nor2_1 U6720 ( .ip1(n7254), .ip2(n7253), .op(n7258) );
  nor2_1 U6721 ( .ip1(n7255), .ip2(n7267), .op(n7253) );
  nand2_1 U6722 ( .ip1(n7250), .ip2(n7243), .op(n7244) );
  nand2_1 U6723 ( .ip1(n7217), .ip2(n7095), .op(n7211) );
  inv_1 U6724 ( .ip(i_i2c_ic_sda_tx_hold_sync[12]), .op(n7095) );
  nor2_1 U6725 ( .ip1(n7224), .ip2(i_i2c_ic_sda_tx_hold_sync[11]), .op(n7217)
         );
  nor2_1 U6726 ( .ip1(n7274), .ip2(n7271), .op(n7265) );
  nor2_1 U6727 ( .ip1(n8897), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[9]), .op(n8915) );
  nor2_1 U6728 ( .ip1(n8143), .ip2(n8142), .op(n8196) );
  nand2_1 U6729 ( .ip1(n8086), .ip2(n8085), .op(n8104) );
  nor2_1 U6730 ( .ip1(n8057), .ip2(n8056), .op(n8112) );
  nor2_1 U6731 ( .ip1(n8881), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[14]), .op(n8057) );
  nor2_1 U6732 ( .ip1(n8106), .ip2(n8103), .op(n8120) );
  nor2_1 U6733 ( .ip1(n8895), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[10]), .op(n8103) );
  nor2_1 U6734 ( .ip1(n8897), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[9]), 
        .op(n8118) );
  and2_1 U6735 ( .ip1(n10768), .ip2(n10769), .op(n10733) );
  nand2_1 U6736 ( .ip1(n10702), .ip2(n10701), .op(n10734) );
  and2_1 U6737 ( .ip1(n10743), .ip2(n10744), .op(n10741) );
  nand2_1 U6738 ( .ip1(n10692), .ip2(n10691), .op(n10742) );
  and2_1 U6739 ( .ip1(n10739), .ip2(n10740), .op(n10737) );
  nand2_1 U6740 ( .ip1(n10696), .ip2(n10695), .op(n10738) );
  and2_1 U6741 ( .ip1(n10737), .ip2(n10738), .op(n10735) );
  nand2_1 U6742 ( .ip1(n10698), .ip2(n10697), .op(n10736) );
  nand2_1 U6743 ( .ip1(n8599), .ip2(n8598), .op(n8600) );
  nor2_1 U6744 ( .ip1(n8688), .ip2(n8687), .op(n8710) );
  nor2_1 U6745 ( .ip1(n8653), .ip2(n8652), .op(n8662) );
  nor2_1 U6746 ( .ip1(n8881), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[14]), .op(n8653) );
  nor2_1 U6747 ( .ip1(n8897), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[9]), .op(n8678) );
  xnor2_1 U6748 ( .ip1(n7969), .ip2(n6743), .op(n9030) );
  nand2_1 U6749 ( .ip1(n6764), .ip2(n6742), .op(n6743) );
  inv_1 U6750 ( .ip(n9011), .op(n6760) );
  nor2_1 U6751 ( .ip1(n6817), .ip2(n6816), .op(n6818) );
  nand2_1 U6752 ( .ip1(n6814), .ip2(n6813), .op(n6819) );
  nand2_1 U6753 ( .ip1(n6812), .ip2(n6811), .op(n6813) );
  nand2_1 U6754 ( .ip1(n8749), .ip2(n8748), .op(n8750) );
  inv_1 U6755 ( .ip(n8969), .op(n8730) );
  inv_1 U6756 ( .ip(n8970), .op(n6744) );
  nor2_1 U6757 ( .ip1(n8842), .ip2(n8841), .op(n8864) );
  nor2_1 U6758 ( .ip1(n8806), .ip2(n8805), .op(n8815) );
  nor2_1 U6759 ( .ip1(n8881), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[14]), .op(n8806) );
  nor2_1 U6760 ( .ip1(n8822), .ip2(n8821), .op(n8834) );
  nor2_1 U6761 ( .ip1(n8895), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[10]), .op(n8822) );
  nor2_1 U6762 ( .ip1(n8897), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[9]), .op(n8832) );
  nor2_1 U6763 ( .ip1(n5641), .ip2(i_ssi_mwcr[0]), .op(n5644) );
  nand2_1 U6764 ( .ip1(n5569), .ip2(n5642), .op(n5589) );
  nor2_1 U6765 ( .ip1(n5282), .ip2(n5566), .op(n5567) );
  inv_1 U6766 ( .ip(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[5]), .op(n5397) );
  inv_1 U6767 ( .ip(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[10]), .op(n5843)
         );
  inv_1 U6768 ( .ip(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[6]), .op(n5838) );
  inv_1 U6769 ( .ip(n6356), .op(n8051) );
  xnor2_1 U6770 ( .ip1(n5565), .ip2(i_ssi_dfs[2]), .op(n5566) );
  mux2_1 U6771 ( .ip1(n7279), .ip2(i_i2c_ic_sda_tx_hold_sync[6]), .s(n7321), 
        .op(n7828) );
  xnor2_1 U6772 ( .ip1(n7278), .ip2(n7277), .op(n7279) );
  nand2_1 U6773 ( .ip1(n7273), .ip2(n7272), .op(n7278) );
  nand2_1 U6774 ( .ip1(n7897), .ip2(n7896), .op(n7899) );
  nand2_1 U6775 ( .ip1(n7206), .ip2(n7243), .op(n7207) );
  nor2_1 U6776 ( .ip1(n7230), .ip2(n7205), .op(n7206) );
  xnor2_1 U6777 ( .ip1(i_i2c_ic_sda_tx_hold_sync[11]), .ip2(n7228), .op(n7229)
         );
  nor2_1 U6778 ( .ip1(n7226), .ip2(n5471), .op(n7227) );
  nand2_1 U6779 ( .ip1(n7102), .ip2(n7243), .op(n7111) );
  nor2_1 U6780 ( .ip1(n7230), .ip2(n7097), .op(n7102) );
  nand2_1 U6781 ( .ip1(n7204), .ip2(n7096), .op(n7097) );
  nor2_1 U6782 ( .ip1(n8949), .ip2(n8948), .op(n8955) );
  nand2_1 U6783 ( .ip1(n8938), .ip2(n8937), .op(n8949) );
  nand2_1 U6784 ( .ip1(n8912), .ip2(n8911), .op(n8913) );
  inv_1 U6785 ( .ip(n8919), .op(n8911) );
  nand2_1 U6786 ( .ip1(n8906), .ip2(n5456), .op(n8912) );
  xnor2_1 U6787 ( .ip1(n7937), .ip2(n6726), .op(n8966) );
  nand2_1 U6788 ( .ip1(n6764), .ip2(n6725), .op(n6726) );
  nor2_1 U6789 ( .ip1(n7987), .ip2(n7986), .op(n7992) );
  nand2_1 U6790 ( .ip1(n8115), .ip2(n8114), .op(n8116) );
  inv_1 U6791 ( .ip(n8122), .op(n8114) );
  nand2_1 U6792 ( .ip1(n8109), .ip2(n5445), .op(n8115) );
  nand2_1 U6793 ( .ip1(n8104), .ip2(n8120), .op(n8109) );
  inv_1 U6794 ( .ip(n7001), .op(n7005) );
  inv_1 U6795 ( .ip(n7011), .op(n7002) );
  nor4_1 U6796 ( .ip1(i_i2c_ic_sda_rx_hold_sync[3]), .ip2(
        i_i2c_ic_sda_rx_hold_sync[2]), .ip3(i_i2c_ic_sda_rx_hold_sync[1]), 
        .ip4(i_i2c_ic_sda_rx_hold_sync[0]), .op(n7011) );
  and2_1 U6797 ( .ip1(n10733), .ip2(n10734), .op(n10770) );
  nand2_1 U6798 ( .ip1(n10704), .ip2(n10703), .op(n10771) );
  inv_1 U6799 ( .ip(n10865), .op(n10762) );
  nor2_1 U6800 ( .ip1(n8635), .ip2(n8634), .op(n8641) );
  nand2_1 U6801 ( .ip1(n8625), .ip2(n8624), .op(n8635) );
  and2_1 U6802 ( .ip1(n8633), .ip2(n8632), .op(n8634) );
  nor2_1 U6803 ( .ip1(n8622), .ip2(n8621), .op(n8643) );
  nand2_1 U6804 ( .ip1(n8614), .ip2(n8613), .op(n8622) );
  and2_1 U6805 ( .ip1(n8638), .ip2(n8620), .op(n8621) );
  nand2_1 U6806 ( .ip1(n6908), .ip2(n6910), .op(n6888) );
  nor2_1 U6807 ( .ip1(n6928), .ip2(n6625), .op(n6890) );
  inv_1 U6808 ( .ip(n9030), .op(n8741) );
  nor2_1 U6809 ( .ip1(n6821), .ip2(n6820), .op(n6822) );
  nand2_1 U6810 ( .ip1(n6797), .ip2(n6796), .op(n6821) );
  and2_1 U6811 ( .ip1(n6819), .ip2(n6818), .op(n6820) );
  nor2_1 U6812 ( .ip1(n6789), .ip2(n6788), .op(n6797) );
  nor2_1 U6813 ( .ip1(n8787), .ip2(n8786), .op(n8793) );
  nand2_1 U6814 ( .ip1(n8776), .ip2(n8775), .op(n8787) );
  and2_1 U6815 ( .ip1(n8785), .ip2(n8784), .op(n8786) );
  nor2_1 U6816 ( .ip1(n8773), .ip2(n8772), .op(n8795) );
  nand2_1 U6817 ( .ip1(n8765), .ip2(n8764), .op(n8773) );
  and2_1 U6818 ( .ip1(n8790), .ip2(n8771), .op(n8772) );
  nand4_1 U6819 ( .ip1(n6931), .ip2(n6894), .ip3(n6936), .ip4(n6704), .op(
        n6705) );
  and2_1 U6820 ( .ip1(n10770), .ip2(n10771), .op(n10772) );
  nand2_1 U6821 ( .ip1(n10706), .ip2(n10705), .op(n10773) );
  and2_1 U6822 ( .ip1(n10521), .ip2(i_ssi_U_regfile_ctrlr1_int[7]), .op(n5348)
         );
  nor2_1 U6823 ( .ip1(n5496), .ip2(n5434), .op(n5497) );
  xnor2_1 U6824 ( .ip1(i_ssi_U_mstfsm_frame_cnt[0]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[0]), .op(n5434) );
  xnor2_1 U6825 ( .ip1(n5405), .ip2(n5490), .op(n5491) );
  xor2_1 U6826 ( .ip1(i_ssi_U_mstfsm_frame_cnt[12]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[12]), .op(n5490) );
  or2_1 U6827 ( .ip1(i_ssi_baudr[5]), .ip2(i_ssi_baudr[6]), .op(n6214) );
  nand2_1 U6828 ( .ip1(n6271), .ip2(n10395), .op(n6272) );
  nor2_1 U6829 ( .ip1(n6270), .ip2(n6269), .op(n6271) );
  nand2_1 U6830 ( .ip1(n7583), .ip2(n6223), .op(n6269) );
  xnor2_1 U6831 ( .ip1(i_ssi_baudr[8]), .ip2(n6264), .op(n6265) );
  nand2_1 U6832 ( .ip1(n6263), .ip2(n6262), .op(n6264) );
  nor2_1 U6833 ( .ip1(n6261), .ip2(n5256), .op(n6262) );
  nand2_1 U6834 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[1]), 
        .ip2(n8004), .op(n7388) );
  nand2_1 U6835 ( .ip1(n5306), .ip2(n5797), .op(n5799) );
  nand2_1 U6836 ( .ip1(n5306), .ip2(n5837), .op(n5841) );
  nand2_1 U6837 ( .ip1(n6084), .ip2(n6083), .op(n6088) );
  nand2_1 U6838 ( .ip1(n6082), .ip2(n6081), .op(n6083) );
  nor2_1 U6839 ( .ip1(n6080), .ip2(n6079), .op(n6082) );
  inv_1 U6840 ( .ip(i_ssi_U_shift_U_tx_shifter_tx_buffer[5]), .op(n6059) );
  inv_2 U6841 ( .ip(n6040), .op(n6061) );
  xnor2_1 U6842 ( .ip1(n8070), .ip2(n6352), .op(n6444) );
  nand2_1 U6843 ( .ip1(n6434), .ip2(n6433), .op(n6436) );
  nor2_1 U6844 ( .ip1(n6431), .ip2(n6432), .op(n6433) );
  inv_1 U6845 ( .ip(n6428), .op(n6434) );
  nand2_1 U6846 ( .ip1(n6420), .ip2(n6419), .op(n6427) );
  nor2_1 U6847 ( .ip1(n6421), .ip2(n5468), .op(n6419) );
  nand2_1 U6848 ( .ip1(n6411), .ip2(n5418), .op(n6420) );
  or4_1 U6849 ( .ip1(i_apb_paddr[30]), .ip2(i_apb_paddr[28]), .ip3(
        i_apb_paddr[27]), .ip4(i_apb_paddr[24]), .op(n5861) );
  nor2_1 U6850 ( .ip1(n7343), .ip2(n11080), .op(n7857) );
  nor2_1 U6851 ( .ip1(n7876), .ip2(n7906), .op(n7886) );
  nand2_1 U6852 ( .ip1(n7884), .ip2(n7883), .op(n7885) );
  nor4_1 U6853 ( .ip1(i_i2c_ic_sda_tx_hold_sync[3]), .ip2(
        i_i2c_ic_sda_tx_hold_sync[4]), .ip3(n7127), .ip4(n7126), .op(n7128) );
  nand2_1 U6854 ( .ip1(n7161), .ip2(n7125), .op(n7126) );
  or4_1 U6855 ( .ip1(i_i2c_ic_sda_tx_hold_sync[7]), .ip2(
        i_i2c_ic_sda_tx_hold_sync[8]), .ip3(i_i2c_ic_sda_tx_hold_sync[6]), 
        .ip4(i_i2c_ic_sda_tx_hold_sync[5]), .op(n7127) );
  xnor2_1 U6856 ( .ip1(i_i2c_ic_sda_tx_hold_sync[13]), .ip2(n7215), .op(n7216)
         );
  nor2_1 U6857 ( .ip1(n7213), .ip2(n5471), .op(n7214) );
  xnor2_1 U6858 ( .ip1(i_i2c_ic_sda_tx_hold_sync[12]), .ip2(n7222), .op(n7223)
         );
  nor2_1 U6859 ( .ip1(n7220), .ip2(n5471), .op(n7221) );
  inv_1 U6860 ( .ip(n8962), .op(n8963) );
  nor2_1 U6861 ( .ip1(n9096), .ip2(n6910), .op(n6699) );
  nor4_1 U6862 ( .ip1(n9584), .ip2(n9583), .ip3(
        i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_slv_1_sync_N2), .ip4(n9607), .op(
        n9587) );
  nor3_1 U6863 ( .ip1(n9634), .ip2(n9602), .ip3(n9608), .op(n9589) );
  nor3_1 U6864 ( .ip1(n9620), .ip2(n9617), .ip3(n9594), .op(n9598) );
  nor3_1 U6865 ( .ip1(n10782), .ip2(n10781), .ip3(n10881), .op(n10784) );
  nand2_1 U6866 ( .ip1(n10917), .ip2(n10727), .op(n10730) );
  nand4_1 U6867 ( .ip1(n7655), .ip2(n6526), .ip3(n6525), .ip4(n7661), .op(
        n6527) );
  nor4_1 U6868 ( .ip1(n7671), .ip2(n7666), .ip3(n7659), .ip4(n6523), .op(n6526) );
  nand4_1 U6869 ( .ip1(n7644), .ip2(n6505), .ip3(n7643), .ip4(n7642), .op(
        n6528) );
  nand4_1 U6870 ( .ip1(n6502), .ip2(n7653), .ip3(n7636), .ip4(n7638), .op(
        n6503) );
  nor2_1 U6871 ( .ip1(n8587), .ip2(n8586), .op(n8605) );
  nand2_1 U6872 ( .ip1(n6629), .ip2(n6628), .op(n6638) );
  nand4_1 U6873 ( .ip1(n6636), .ip2(n6635), .ip3(n6634), .ip4(n6633), .op(
        n6637) );
  nand2_1 U6874 ( .ip1(n6890), .ip2(n6627), .op(n6894) );
  inv_1 U6875 ( .ip(n6929), .op(n6627) );
  nand2_1 U6876 ( .ip1(n9727), .ip2(n6887), .op(n6892) );
  nor2_1 U6877 ( .ip1(n6910), .ip2(n6909), .op(n6911) );
  and2_1 U6878 ( .ip1(n6626), .ip2(n6703), .op(n6908) );
  nor2_1 U6879 ( .ip1(n6727), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[15]), .op(n6830) );
  nor2_1 U6880 ( .ip1(n8736), .ip2(n8735), .op(n8755) );
  and2_1 U6881 ( .ip1(n10709), .ip2(n10710), .op(n10718) );
  nand2_1 U6882 ( .ip1(n10682), .ip2(n10681), .op(n10717) );
  nor2_1 U6883 ( .ip1(n9908), .ip2(n9829), .op(n11579) );
  nand2_1 U6884 ( .ip1(n6980), .ip2(n5694), .op(n6111) );
  nand2_1 U6885 ( .ip1(n6139), .ip2(n5717), .op(n5751) );
  nor2_1 U6886 ( .ip1(n5716), .ip2(n6111), .op(n5695) );
  nor2_1 U6887 ( .ip1(n5482), .ip2(n5751), .op(n5692) );
  nand2_1 U6888 ( .ip1(n5513), .ip2(n5512), .op(n5521) );
  xnor2_1 U6889 ( .ip1(n5511), .ip2(n5510), .op(n5512) );
  nand2_1 U6890 ( .ip1(n10397), .ip2(n6259), .op(n10401) );
  nand2_1 U6891 ( .ip1(n9820), .ip2(n6199), .op(n9908) );
  nand3_1 U6892 ( .ip1(n6582), .ip2(n6584), .ip3(n10008), .op(n6589) );
  nand2_1 U6893 ( .ip1(n9384), .ip2(n6586), .op(n6582) );
  nor3_1 U6894 ( .ip1(n10325), .ip2(n10324), .ip3(n10323), .op(n10326) );
  xnor2_1 U6895 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[4]), .ip2(i_ssi_baudr[5]), .op(
        n10312) );
  xnor2_1 U6896 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[6]), .ip2(n5256), .op(n10313)
         );
  xnor2_1 U6897 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[2]), .ip2(n10310), .op(n10311)
         );
  nor4_1 U6898 ( .ip1(n10318), .ip2(n10317), .ip3(n10316), .ip4(n10315), .op(
        n10328) );
  and2_1 U6899 ( .ip1(n5597), .ip2(n5596), .op(n5438) );
  nor4_1 U6900 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[23]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[22]), .ip3(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[25]), .ip4(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[18]), .op(n6556) );
  nand2_1 U6901 ( .ip1(n6152), .ip2(n6144), .op(n6154) );
  inv_1 U6902 ( .ip(i_ssi_baudr[3]), .op(n6240) );
  xnor2_1 U6903 ( .ip1(i_ssi_baudr[13]), .ip2(n5402), .op(n6229) );
  xnor2_1 U6904 ( .ip1(n6224), .ip2(n10375), .op(n6235) );
  nand2_1 U6905 ( .ip1(n10395), .ip2(n5451), .op(n6221) );
  or2_1 U6906 ( .ip1(n6218), .ip2(n6217), .op(n6219) );
  nor2_1 U6907 ( .ip1(n6242), .ip2(n6247), .op(n6252) );
  nand4_1 U6908 ( .ip1(n6246), .ip2(n10323), .ip3(n6245), .ip4(n6244), .op(
        n6247) );
  nand2_1 U6909 ( .ip1(n5739), .ip2(n6189), .op(n6192) );
  nand2_1 U6910 ( .ip1(n5625), .ip2(n5481), .op(n5626) );
  nand2_1 U6911 ( .ip1(n5659), .ip2(n5658), .op(n5660) );
  nor2_1 U6912 ( .ip1(n5657), .ip2(n5656), .op(n5658) );
  nor2_1 U6913 ( .ip1(n5344), .ip2(n5343), .op(n5375) );
  inv_1 U6914 ( .ip(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[3]), .op(n5810) );
  nand2_1 U6915 ( .ip1(n5444), .ip2(n5363), .op(n5849) );
  nand2_1 U6916 ( .ip1(n5739), .ip2(n6164), .op(n6167) );
  nor2_1 U6917 ( .ip1(n6860), .ip2(n6859), .op(n6863) );
  nor2_1 U6918 ( .ip1(n7419), .ip2(n11156), .op(n7429) );
  nand2_1 U6919 ( .ip1(n6386), .ip2(n5417), .op(n6387) );
  nand2_1 U6920 ( .ip1(n6382), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[11]), .op(n6386) );
  nor2_1 U6921 ( .ip1(n6453), .ip2(n6452), .op(n6454) );
  nand2_1 U6922 ( .ip1(n5416), .ip2(n5463), .op(n6453) );
  nor2_1 U6923 ( .ip1(n6451), .ip2(n6450), .op(n6452) );
  nand2_1 U6924 ( .ip1(n6438), .ip2(n6437), .op(n6455) );
  nand2_1 U6925 ( .ip1(n6427), .ip2(n6426), .op(n6438) );
  nor2_1 U6926 ( .ip1(n6436), .ip2(n6435), .op(n6437) );
  nor2_1 U6927 ( .ip1(n6425), .ip2(n5469), .op(n6426) );
  nor2_1 U6928 ( .ip1(n11156), .ip2(n11160), .op(n7746) );
  nor2_1 U6929 ( .ip1(n6288), .ip2(n10514), .op(n6289) );
  nor2_1 U6930 ( .ip1(n10483), .ip2(n6302), .op(n10500) );
  nand2_1 U6931 ( .ip1(n6301), .ip2(n6300), .op(n6302) );
  nor2_1 U6932 ( .ip1(n6299), .ip2(n6298), .op(n6300) );
  inv_1 U6933 ( .ip(n10484), .op(n6301) );
  nand2_1 U6934 ( .ip1(n10993), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[13]), .op(n10267) );
  nor2_1 U6935 ( .ip1(n9010), .ip2(n9012), .op(n10985) );
  inv_1 U6936 ( .ip(n9666), .op(n9429) );
  nand2_1 U6937 ( .ip1(n9429), .ip2(n6699), .op(n8334) );
  nand2_1 U6938 ( .ip1(n8208), .ip2(n8207), .op(n10918) );
  nor4_1 U6939 ( .ip1(n8001), .ip2(n8000), .ip3(n7999), .ip4(n7998), .op(n8002) );
  mux2_1 U6940 ( .ip1(n11769), .ip2(n7718), .s(n7717), .op(n11174) );
  nor2_1 U6941 ( .ip1(n8243), .ip2(n8242), .op(n8269) );
  nand4_1 U6942 ( .ip1(n9588), .ip2(n9587), .ip3(n9586), .ip4(n9585), .op(
        n9606) );
  nor4_1 U6943 ( .ip1(n9582), .ip2(n9581), .ip3(n9580), .ip4(n9579), .op(n9588) );
  nand4_1 U6944 ( .ip1(n9589), .ip2(n9620), .ip3(n9575), .ip4(n9574), .op(
        n9647) );
  nand4_1 U6945 ( .ip1(n9598), .ip2(n9597), .ip3(n9596), .ip4(n9595), .op(
        n9623) );
  nand4_1 U6946 ( .ip1(n11346), .ip2(n11339), .ip3(n11342), .ip4(n11352), .op(
        n9571) );
  nand2_1 U6947 ( .ip1(n11284), .ip2(n7924), .op(n9095) );
  nand2_1 U6948 ( .ip1(n11316), .ip2(n8295), .op(n8531) );
  nor2_1 U6949 ( .ip1(n8220), .ip2(n8219), .op(n11292) );
  nand2_1 U6950 ( .ip1(n7036), .ip2(n7035), .op(n9751) );
  nand2_1 U6951 ( .ip1(n7041), .ip2(n7040), .op(n7042) );
  and2_1 U6952 ( .ip1(n10881), .ip2(n10782), .op(n10775) );
  nor3_1 U6953 ( .ip1(n10779), .ip2(n10777), .ip3(n10837), .op(n10712) );
  inv_1 U6954 ( .ip(n7072), .op(n6915) );
  nand2_1 U6955 ( .ip1(i_i2c_tx_push), .ip2(n7489), .op(n9783) );
  nand2_1 U6956 ( .ip1(n6941), .ip2(n7073), .op(n6877) );
  nor3_1 U6957 ( .ip1(n6905), .ip2(n6881), .ip3(n6877), .op(n8332) );
  inv_1 U6958 ( .ip(n6928), .op(n6912) );
  inv_1 U6959 ( .ip(n6341), .op(n6464) );
  nor2_1 U6960 ( .ip1(n7420), .ip2(n6996), .op(n9612) );
  nand2_1 U6961 ( .ip1(n7689), .ip2(n10569), .op(n6996) );
  nand3_1 U6962 ( .ip1(n6714), .ip2(n6713), .ip3(n6712), .op(n6952) );
  and2_1 U6963 ( .ip1(n10718), .ip2(n10717), .op(n10724) );
  nand2_1 U6964 ( .ip1(n10716), .ip2(n10715), .op(n10723) );
  nand2_1 U6965 ( .ip1(n10414), .ip2(n6470), .op(n6471) );
  nor2_1 U6966 ( .ip1(n9658), .ip2(n9154), .op(n8344) );
  nand2_1 U6967 ( .ip1(n11583), .ip2(n11582), .op(n11586) );
  or2_1 U6968 ( .ip1(n11579), .ip2(n11580), .op(n11583) );
  nor2_1 U6969 ( .ip1(i_ssi_rx_wr_addr[2]), .ip2(n11223), .op(n10064) );
  nand2_1 U6970 ( .ip1(i_ssi_rx_full), .ip2(n11165), .op(n9368) );
  nor2_1 U6971 ( .ip1(n5323), .ip2(n11223), .op(n10065) );
  nand2_1 U6972 ( .ip1(n6134), .ip2(n5281), .op(n6135) );
  nand2_1 U6973 ( .ip1(n5690), .ip2(n10231), .op(n6140) );
  mux2_1 U6974 ( .ip1(n9851), .ip2(n9850), .s(n11568), .op(n9853) );
  nor2_1 U6975 ( .ip1(n5691), .ip2(n7629), .op(n5756) );
  nor2_1 U6976 ( .ip1(n5281), .ip2(n5574), .op(n5716) );
  inv_1 U6977 ( .ip(n5756), .op(n5717) );
  nand4_1 U6978 ( .ip1(n6037), .ip2(n6036), .ip3(n6035), .ip4(n6034), .op(
        n6038) );
  nand4_1 U6979 ( .ip1(n6025), .ip2(n6024), .ip3(n6023), .ip4(n6022), .op(
        n6026) );
  nand4_1 U6980 ( .ip1(n5912), .ip2(n5911), .ip3(n5910), .ip4(n5909), .op(
        n5913) );
  nand4_1 U6981 ( .ip1(n5964), .ip2(n5963), .ip3(n5962), .ip4(n5961), .op(
        n5965) );
  nor3_1 U6982 ( .ip1(i_ssi_tx_wr_addr[2]), .ip2(i_ssi_tx_wr_addr[1]), .ip3(
        n10166), .op(n10170) );
  nor3_1 U6983 ( .ip1(i_ssi_tx_wr_addr[2]), .ip2(n11212), .ip3(n10166), .op(
        n10167) );
  nor3_1 U6984 ( .ip1(i_ssi_tx_wr_addr[1]), .ip2(n10165), .ip3(n10166), .op(
        n10169) );
  nor3_1 U6985 ( .ip1(n10165), .ip2(n11212), .ip3(n10166), .op(n10168) );
  inv_1 U6986 ( .ip(n5557), .op(n5508) );
  inv_1 U6987 ( .ip(i_ssi_U_mstfsm_c_state[3]), .op(n6281) );
  xnor2_1 U6988 ( .ip1(n10363), .ip2(n10362), .op(n5439) );
  nor2_1 U6989 ( .ip1(n5371), .ip2(n10391), .op(n10392) );
  nor3_1 U6990 ( .ip1(n7531), .ip2(n11126), .ip3(n11123), .op(n11675) );
  inv_1 U6991 ( .ip(n11691), .op(n9900) );
  nor2_1 U6992 ( .ip1(n7783), .ip2(n7802), .op(n11568) );
  nor2_1 U6993 ( .ip1(n7783), .ip2(n9786), .op(n11567) );
  nor2_1 U6994 ( .ip1(n11616), .ip2(n9786), .op(n9852) );
  nor2_1 U6995 ( .ip1(n11616), .ip2(n7802), .op(n11573) );
  nand2_1 U6996 ( .ip1(n6600), .ip2(n7607), .op(n9786) );
  nand2_1 U6997 ( .ip1(n10112), .ip2(n10111), .op(n10116) );
  nor2_1 U6998 ( .ip1(n10024), .ip2(n6574), .op(n11471) );
  nor2_1 U6999 ( .ip1(n11368), .ip2(n11370), .op(n11407) );
  nand2_1 U7000 ( .ip1(n10024), .ip2(n9374), .op(n10008) );
  inv_1 U7001 ( .ip(n6586), .op(n10107) );
  nor2_1 U7002 ( .ip1(n9378), .ip2(n9381), .op(n9380) );
  inv_1 U7003 ( .ip(n10019), .op(n9382) );
  nor4_1 U7004 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[1]), .ip2(
        i_ssi_U_sclkgen_ssi_cnt[2]), .ip3(i_ssi_U_sclkgen_ssi_cnt[3]), .ip4(
        i_ssi_U_sclkgen_ssi_cnt[4]), .op(n10295) );
  nor4_1 U7005 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[9]), .ip2(
        i_ssi_U_sclkgen_ssi_cnt[10]), .ip3(i_ssi_U_sclkgen_ssi_cnt[11]), .ip4(
        i_ssi_U_sclkgen_ssi_cnt[12]), .op(n10297) );
  nor2_1 U7006 ( .ip1(n8386), .ip2(n8385), .op(n11607) );
  nand4_1 U7007 ( .ip1(n6559), .ip2(n6558), .ip3(n6557), .ip4(n6556), .op(
        n7051) );
  nor2_1 U7008 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[24]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[19]), .op(n6559) );
  nor4_1 U7009 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[31]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[29]), .ip3(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[28]), .ip4(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[30]), .op(n6557) );
  nor4_1 U7010 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[27]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[26]), .ip3(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[21]), .ip4(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[20]), .op(n6558) );
  nand2_1 U7011 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[17]), .ip2(n6560), 
        .op(n9070) );
  nor4_1 U7012 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[14]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[16]), .ip3(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[15]), .ip4(n7051), .op(n6560) );
  nand2_1 U7013 ( .ip1(n5739), .ip2(n6156), .op(n6159) );
  nor2_1 U7014 ( .ip1(n7761), .ip2(n9837), .op(n9844) );
  inv_1 U7015 ( .ip(n6240), .op(n10310) );
  nand2_1 U7016 ( .ip1(n10537), .ip2(n9084), .op(n9083) );
  nor4_1 U7017 ( .ip1(n9753), .ip2(n9752), .ip3(n9751), .ip4(n9750), .op(n9762) );
  inv_1 U7018 ( .ip(n7048), .op(n9765) );
  nand2_1 U7019 ( .ip1(n11175), .ip2(n11174), .op(n7750) );
  or2_1 U7020 ( .ip1(n7420), .ip2(n7428), .op(n11157) );
  nor2_1 U7021 ( .ip1(i_i2c_scl_lcnt_cmplt), .ip2(n8306), .op(n7741) );
  or2_1 U7022 ( .ip1(n7413), .ip2(n7412), .op(n8439) );
  nor2_1 U7023 ( .ip1(n7385), .ip2(n7384), .op(n7413) );
  nand2_1 U7024 ( .ip1(n5739), .ip2(n5714), .op(n5730) );
  nand2_1 U7025 ( .ip1(n5739), .ip2(n6146), .op(n6149) );
  inv_1 U7026 ( .ip(n11220), .op(n11223) );
  nand2_1 U7027 ( .ip1(n10222), .ip2(n10221), .op(n11235) );
  nor2_1 U7028 ( .ip1(n11222), .ip2(n11221), .op(n11220) );
  and2_1 U7029 ( .ip1(n9693), .ip2(n11780), .op(n11217) );
  and2_1 U7030 ( .ip1(n9692), .ip2(n11780), .op(n6991) );
  inv_1 U7031 ( .ip(n11124), .op(n11164) );
  nand2_1 U7032 ( .ip1(n11782), .ip2(i_ssi_U_fifo_U_rx_fifo_empty_n), .op(
        n11124) );
  nand2_1 U7033 ( .ip1(n6666), .ip2(n6665), .op(n6667) );
  or2_1 U7034 ( .ip1(n6669), .ip2(n6664), .op(n6665) );
  mux2_1 U7035 ( .ip1(n6854), .ip2(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[2]), 
        .s(n6853), .op(n7053) );
  inv_1 U7036 ( .ip(n11251), .op(n11256) );
  mux2_1 U7037 ( .ip1(n6674), .ip2(i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[1]), 
        .s(n6673), .op(n6838) );
  nand2_1 U7038 ( .ip1(n6672), .ip2(n6671), .op(n6673) );
  mux2_1 U7039 ( .ip1(n6862), .ip2(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[1]), 
        .s(n6861), .op(n7055) );
  nor2_1 U7040 ( .ip1(n11253), .ip2(n11252), .op(n11251) );
  nand2_1 U7041 ( .ip1(i_i2c_rx_push_sync), .ip2(n11191), .op(n11197) );
  inv_1 U7042 ( .ip(i_i2c_rx_pop), .op(n11209) );
  mux2_1 U7043 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[0]), .ip2(n6678), 
        .s(n6677), .op(n6988) );
  nor2_1 U7044 ( .ip1(n6676), .ip2(n6675), .op(n6677) );
  inv_1 U7045 ( .ip(n9783), .op(n9766) );
  inv_1 U7046 ( .ip(i_i2c_tx_pop_sync), .op(n11261) );
  or2_1 U7047 ( .ip1(n10011), .ip2(n10010), .op(n10012) );
  nor3_1 U7048 ( .ip1(n9093), .ip2(n9092), .ip3(n9091), .op(n10294) );
  or4_1 U7049 ( .ip1(n6224), .ip2(i_ssi_baudr[14]), .ip3(n11652), .ip4(
        i_ssi_baudr[13]), .op(n9092) );
  nor2_1 U7050 ( .ip1(n10443), .ip2(n10442), .op(n10444) );
  nor2_1 U7051 ( .ip1(n10455), .ip2(n10454), .op(n10456) );
  nor2_1 U7052 ( .ip1(n10449), .ip2(n10448), .op(n10450) );
  nand2_1 U7053 ( .ip1(n5279), .ip2(n5460), .op(n5888) );
  nand2_1 U7054 ( .ip1(n6092), .ip2(n6091), .op(n6093) );
  nor2_1 U7055 ( .ip1(n10461), .ip2(n10460), .op(n10462) );
  nor2_1 U7056 ( .ip1(n10433), .ip2(n10432), .op(n10434) );
  nor2_1 U7057 ( .ip1(n10467), .ip2(n10466), .op(n10468) );
  nand3_1 U7058 ( .ip1(n10024), .ip2(n10108), .ip3(n9374), .op(n6569) );
  inv_1 U7059 ( .ip(n11471), .op(n6570) );
  nor2_1 U7060 ( .ip1(n6564), .ip2(i_apb_U_DW_apb_ahbsif_pipeline_c), .op(
        n6565) );
  or2_1 U7061 ( .ip1(n9927), .ip2(n6961), .op(n9930) );
  nor2_1 U7062 ( .ip1(n11258), .ip2(n6965), .op(n6961) );
  inv_1 U7063 ( .ip(n9627), .op(n8563) );
  nand2_1 U7064 ( .ip1(n7747), .ip2(n8523), .op(n9631) );
  nand2_1 U7065 ( .ip1(n8563), .ip2(n9628), .op(n7747) );
  nand3_1 U7066 ( .ip1(n7746), .ip2(n7754), .ip3(n7745), .op(n9627) );
  nor2_1 U7067 ( .ip1(n7426), .ip2(n7425), .op(n9999) );
  nor2_1 U7068 ( .ip1(n7918), .ip2(n7424), .op(n7425) );
  nand2_1 U7069 ( .ip1(n11772), .ip2(n7421), .op(n8523) );
  nand2_1 U7070 ( .ip1(n7429), .ip2(n7754), .op(n7421) );
  inv_1 U7071 ( .ip(n11772), .op(n11160) );
  nand2_1 U7072 ( .ip1(n6546), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[12]), .op(n10244) );
  inv_1 U7073 ( .ip(n10242), .op(n6546) );
  inv_1 U7074 ( .ip(n10237), .op(n6545) );
  nand2_1 U7075 ( .ip1(n6544), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[10]), .op(n10237) );
  inv_1 U7076 ( .ip(n10228), .op(n6544) );
  inv_1 U7077 ( .ip(n6464), .op(n10275) );
  inv_1 U7078 ( .ip(n10575), .op(n11158) );
  inv_1 U7079 ( .ip(n11717), .op(n11719) );
  nor2_1 U7080 ( .ip1(n11719), .ip2(n11718), .op(n11722) );
  nor2_1 U7081 ( .ip1(n11716), .ip2(n11715), .op(n11717) );
  inv_1 U7082 ( .ip(n11714), .op(n11711) );
  nand2_1 U7083 ( .ip1(n10492), .ip2(n10491), .op(n10493) );
  nor2_1 U7084 ( .ip1(n10488), .ip2(n10487), .op(n10492) );
  nor2_1 U7085 ( .ip1(n10494), .ip2(n10493), .op(n10495) );
  nor2_1 U7086 ( .ip1(n10502), .ip2(n10501), .op(n10516) );
  nand2_1 U7087 ( .ip1(n10500), .ip2(n10499), .op(n10501) );
  nor2_1 U7088 ( .ip1(n10509), .ip2(n10508), .op(n10510) );
  nor2_1 U7089 ( .ip1(n10521), .ip2(n10520), .op(n10522) );
  inv_1 U7090 ( .ip(i_ssi_U_mstfsm_frame_cnt[14]), .op(n6305) );
  inv_1 U7091 ( .ip(i_ssi_U_mstfsm_frame_cnt[15]), .op(n10544) );
  nor2_1 U7092 ( .ip1(n9746), .ip2(n9769), .op(n9745) );
  nor2_1 U7093 ( .ip1(n11194), .ip2(n9746), .op(n9747) );
  inv_1 U7094 ( .ip(n7433), .op(n7434) );
  nand2_1 U7095 ( .ip1(n7435), .ip2(n7436), .op(n8559) );
  or2_1 U7096 ( .ip1(i_i2c_ic_clr_intr_en), .ip2(i_i2c_ic_clr_tx_abrt_en), 
        .op(n7436) );
  nand2_1 U7097 ( .ip1(n7918), .ip2(n7917), .op(n10002) );
  nor2_1 U7098 ( .ip1(n11058), .ip2(n11057), .op(n11059) );
  and4_1 U7099 ( .ip1(n10275), .ip2(n9999), .ip3(n9998), .ip4(n9997), .op(
        n11105) );
  inv_1 U7100 ( .ip(n11099), .op(n10003) );
  inv_1 U7101 ( .ip(n11105), .op(n10004) );
  nor2_1 U7102 ( .ip1(n11043), .ip2(n11042), .op(n11040) );
  nand2_1 U7103 ( .ip1(n11036), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[13]), .op(n11043) );
  nor2_1 U7104 ( .ip1(n7741), .ip2(n7743), .op(n8348) );
  nor2_1 U7105 ( .ip1(n10267), .ip2(n9054), .op(n10268) );
  nor2_1 U7106 ( .ip1(n9053), .ip2(n10984), .op(n10990) );
  nand2_1 U7107 ( .ip1(n10985), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[11]), .op(n9053) );
  nand2_1 U7108 ( .ip1(n10986), .ip2(n10985), .op(n10989) );
  nor2_1 U7109 ( .ip1(n9012), .ip2(n10984), .op(n10983) );
  nor2_1 U7110 ( .ip1(n10980), .ip2(n10979), .op(n10981) );
  nand2_1 U7111 ( .ip1(n10975), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[6]), .op(n10980) );
  nand2_1 U7112 ( .ip1(n10958), .ip2(n5473), .op(n10974) );
  and2_1 U7113 ( .ip1(n10958), .ip2(n5422), .op(n10969) );
  nand2_1 U7114 ( .ip1(n10958), .ip2(n9949), .op(n10965) );
  inv_1 U7115 ( .ip(n11157), .op(n7754) );
  nor2_1 U7116 ( .ip1(n7702), .ip2(n8522), .op(n7753) );
  nor2_1 U7117 ( .ip1(n7751), .ip2(n7750), .op(n7758) );
  nor2_1 U7118 ( .ip1(n10566), .ip2(n9183), .op(n9639) );
  nand2_1 U7119 ( .ip1(n8323), .ip2(n8322), .op(n10565) );
  nor2_1 U7120 ( .ip1(n8357), .ip2(n10575), .op(n10567) );
  nand3_1 U7121 ( .ip1(n8318), .ip2(n9643), .ip3(n9642), .op(n11116) );
  nand2_1 U7122 ( .ip1(n11773), .ip2(n6997), .op(n8359) );
  nor2_1 U7123 ( .ip1(n9643), .ip2(n9632), .op(n11310) );
  nor2_1 U7124 ( .ip1(n9612), .ip2(n8359), .op(n8322) );
  nand3_1 U7125 ( .ip1(n11773), .ip2(n9612), .ip3(n8318), .op(n9645) );
  nor2_1 U7126 ( .ip1(n10571), .ip2(n8321), .op(n8323) );
  inv_1 U7127 ( .ip(n10565), .op(n8357) );
  inv_1 U7128 ( .ip(n9400), .op(n9401) );
  nand2_1 U7129 ( .ip1(n9737), .ip2(n9736), .op(n9738) );
  nand2_1 U7130 ( .ip1(n8554), .ip2(n8259), .op(n11284) );
  inv_1 U7131 ( .ip(n9402), .op(n9403) );
  nor2_1 U7132 ( .ip1(n8336), .ip2(n8335), .op(n9409) );
  nor2_1 U7133 ( .ip1(n10950), .ip2(n7976), .op(n10951) );
  nand2_1 U7134 ( .ip1(n10946), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[11]), .op(n10950) );
  nor2_1 U7135 ( .ip1(n10945), .ip2(n7990), .op(n10946) );
  nand2_1 U7136 ( .ip1(n10941), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[9]), .op(n10945) );
  nor2_1 U7137 ( .ip1(n10940), .ip2(n7981), .op(n10941) );
  nand2_2 U7138 ( .ip1(n10936), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[7]), .op(n10940) );
  inv_1 U7139 ( .ip(n8801), .op(n11170) );
  nor2_1 U7140 ( .ip1(n5245), .ip2(n6483), .op(n11354) );
  nor2_1 U7141 ( .ip1(n8302), .ip2(n9657), .op(n6483) );
  nand2_1 U7142 ( .ip1(n8554), .ip2(n8296), .op(n7924) );
  nand3_1 U7143 ( .ip1(n8554), .ip2(n8219), .ip3(n7922), .op(n8330) );
  nor2_1 U7144 ( .ip1(n11293), .ip2(n8269), .op(n11299) );
  nor2_1 U7145 ( .ip1(n11292), .ip2(n8272), .op(n8444) );
  nand2_1 U7146 ( .ip1(n11769), .ip2(n11115), .op(n11714) );
  nand2_1 U7147 ( .ip1(n8447), .ip2(n9600), .op(n9608) );
  nor2_1 U7148 ( .ip1(n8534), .ip2(n11114), .op(n8417) );
  nor2_1 U7149 ( .ip1(n8525), .ip2(n7922), .op(n11302) );
  nor2_1 U7150 ( .ip1(n7921), .ip2(n9399), .op(n11301) );
  nor4_1 U7151 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[7]), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[6]), .ip3(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[5]), .ip4(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[4]), .op(n8462) );
  inv_1 U7152 ( .ip(n6926), .op(n9723) );
  nand3_1 U7153 ( .ip1(n7422), .ip2(n7922), .ip3(n8527), .op(n9399) );
  or4_1 U7154 ( .ip1(n8302), .ip2(n8344), .ip3(n8301), .ip4(n8300), .op(n8549)
         );
  nor2_1 U7155 ( .ip1(n8299), .ip2(n8534), .op(n8300) );
  inv_1 U7156 ( .ip(n8554), .op(n8534) );
  nor2_1 U7157 ( .ip1(n9625), .ip2(n9633), .op(n9654) );
  nor2_1 U7158 ( .ip1(n11769), .ip2(n9624), .op(n9625) );
  nor2_1 U7159 ( .ip1(n11721), .ip2(n9605), .op(n9636) );
  nor2_1 U7160 ( .ip1(n11769), .ip2(n9570), .op(n9605) );
  inv_1 U7161 ( .ip(n9608), .op(n9638) );
  nand2_1 U7162 ( .ip1(n9566), .ip2(n11328), .op(n9633) );
  inv_1 U7163 ( .ip(n11769), .op(n11113) );
  nor2_1 U7164 ( .ip1(n8447), .ip2(n7677), .op(n11721) );
  nor2_1 U7165 ( .ip1(n11324), .ip2(n11328), .op(n11344) );
  nor2_1 U7166 ( .ip1(n8417), .ip2(n8535), .op(n8447) );
  inv_1 U7167 ( .ip(n11721), .op(n9566) );
  nand3_1 U7168 ( .ip1(n11713), .ip2(n7633), .ip3(n8447), .op(n8278) );
  nand3_1 U7169 ( .ip1(n7921), .ip2(n7922), .ip3(n8527), .op(n8286) );
  nand2_1 U7170 ( .ip1(n6485), .ip2(n6484), .op(n8282) );
  or2_1 U7171 ( .ip1(n6841), .ip2(n11354), .op(n6485) );
  or2_1 U7172 ( .ip1(n9095), .ip2(n11354), .op(n6484) );
  inv_1 U7173 ( .ip(n8259), .op(n11293) );
  nor3_1 U7174 ( .ip1(n11175), .ip2(n6842), .ip3(n7719), .op(n7713) );
  inv_1 U7175 ( .ip(n5109), .op(n11316) );
  inv_1 U7176 ( .ip(n11141), .op(n11147) );
  nor2_1 U7177 ( .ip1(n11142), .ip2(n11143), .op(n11141) );
  nor2_1 U7178 ( .ip1(n11139), .ip2(n11140), .op(n11138) );
  nor2_1 U7179 ( .ip1(n10805), .ip2(n10732), .op(n10804) );
  nor2_1 U7180 ( .ip1(n10809), .ip2(n10906), .op(n10808) );
  nand2_1 U7181 ( .ip1(n10810), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[12]), .op(n10809) );
  nand2_1 U7182 ( .ip1(n10823), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[4]), .op(n10824) );
  nor2_1 U7183 ( .ip1(n10831), .ip2(n10853), .op(n10823) );
  nand2_1 U7184 ( .ip1(n10830), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[2]), .op(n10831) );
  and2_1 U7185 ( .ip1(n10828), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[1]), .op(n10830) );
  and3_1 U7186 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_count_en), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[0]), .ip3(n5450), .op(n10828)
         );
  inv_1 U7187 ( .ip(n10800), .op(n10802) );
  mux2_1 U7188 ( .ip1(n7048), .ip2(n6536), .s(n6535), .op(n10579) );
  nand3_1 U7189 ( .ip1(n7673), .ip2(n9404), .ip3(n9405), .op(n11277) );
  inv_1 U7190 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[3]), .op(
        n10554) );
  nor2_1 U7191 ( .ip1(n10554), .ip2(n10553), .op(n10555) );
  inv_1 U7192 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[2]), .op(
        n10552) );
  nor2_1 U7193 ( .ip1(n10552), .ip2(n10551), .op(n10550) );
  nand2_1 U7194 ( .ip1(n8439), .ip2(n7414), .op(n10561) );
  inv_1 U7195 ( .ip(n11775), .op(n9777) );
  nand2_1 U7196 ( .ip1(n6897), .ip2(n6313), .op(n6618) );
  nor2_1 U7197 ( .ip1(n9724), .ip2(n6900), .op(n10414) );
  nand2_1 U7198 ( .ip1(n6915), .ip2(n7073), .op(n8217) );
  inv_1 U7199 ( .ip(n11048), .op(n8427) );
  nor3_1 U7200 ( .ip1(n6846), .ip2(n6900), .ip3(n6845), .op(n6847) );
  nor2_1 U7201 ( .ip1(n11252), .ip2(n9782), .op(n11255) );
  nor2_1 U7202 ( .ip1(n8332), .ip2(n8421), .op(n8343) );
  nand3_1 U7203 ( .ip1(n6646), .ip2(n6645), .ip3(n6644), .op(n6647) );
  nand4_1 U7204 ( .ip1(n6951), .ip2(n6950), .ip3(n6949), .ip4(n6948), .op(
        n11045) );
  nand4_1 U7205 ( .ip1(n6924), .ip2(n6951), .ip3(n6923), .ip4(n6945), .op(
        n6925) );
  nor2_1 U7206 ( .ip1(n9742), .ip2(n5245), .op(n11051) );
  nor3_1 U7207 ( .ip1(n9096), .ip2(n5245), .ip3(n8329), .op(n11050) );
  nor3_1 U7208 ( .ip1(n11119), .ip2(n6995), .ip3(n10572), .op(n7689) );
  inv_1 U7209 ( .ip(n11773), .op(n10566) );
  nand2_1 U7210 ( .ip1(n6999), .ip2(n9645), .op(n11311) );
  or2_1 U7211 ( .ip1(n7417), .ip2(n8443), .op(n7743) );
  inv_1 U7212 ( .ip(n8418), .op(n7361) );
  nor2_1 U7213 ( .ip1(n7073), .ip2(n9997), .op(n6874) );
  nand2_1 U7214 ( .ip1(n6939), .ip2(n6873), .op(n6883) );
  inv_1 U7215 ( .ip(n8559), .op(n7488) );
  nand2_1 U7216 ( .ip1(n9727), .ip2(n6477), .op(n9414) );
  nand2_1 U7217 ( .ip1(n7494), .ip2(n7493), .op(n9732) );
  inv_1 U7218 ( .ip(n11283), .op(n11110) );
  nand2_1 U7219 ( .ip1(n8427), .ip2(n8425), .op(n8329) );
  nor2_1 U7220 ( .ip1(n9829), .ip2(n7783), .op(n11576) );
  nor2_1 U7221 ( .ip1(n7802), .ip2(n9785), .op(n11691) );
  nor2_1 U7222 ( .ip1(n11615), .ip2(n7783), .op(n11600) );
  nor2_1 U7223 ( .ip1(n11615), .ip2(n9785), .op(n11587) );
  and2_1 U7224 ( .ip1(n5739), .ip2(n10277), .op(n10284) );
  nor2_1 U7225 ( .ip1(n10280), .ip2(n10340), .op(n10282) );
  nand4_1 U7226 ( .ip1(n6013), .ip2(n6012), .ip3(n6011), .ip4(n6010), .op(
        n6014) );
  nor2_1 U7227 ( .ip1(n5929), .ip2(n5928), .op(n10260) );
  nor2_1 U7228 ( .ip1(n5939), .ip2(n5938), .op(n10258) );
  nand4_1 U7229 ( .ip1(n5937), .ip2(n5936), .ip3(n5935), .ip4(n5934), .op(
        n5938) );
  nor2_1 U7230 ( .ip1(n5989), .ip2(n5988), .op(n10246) );
  nand4_1 U7231 ( .ip1(n5987), .ip2(n5986), .ip3(n5985), .ip4(n5984), .op(
        n5988) );
  nand4_1 U7232 ( .ip1(n5824), .ip2(n5823), .ip3(n5822), .ip4(n5821), .op(
        n5825) );
  nor2_1 U7233 ( .ip1(n5592), .ip2(i_ssi_mwcr[0]), .op(n5715) );
  buf_1 U7234 ( .ip(n10170), .op(n10174) );
  buf_1 U7235 ( .ip(n10170), .op(n10175) );
  buf_1 U7236 ( .ip(n10167), .op(n10173) );
  buf_1 U7237 ( .ip(n10167), .op(n10176) );
  buf_1 U7238 ( .ip(n10169), .op(n10172) );
  buf_1 U7239 ( .ip(n10169), .op(n10177) );
  buf_1 U7240 ( .ip(n10168), .op(n10171) );
  buf_1 U7241 ( .ip(n10168), .op(n10178) );
  buf_1 U7242 ( .ip(n10031), .op(n10032) );
  buf_1 U7243 ( .ip(n10031), .op(n10035) );
  buf_1 U7244 ( .ip(n10033), .op(n10037) );
  buf_1 U7245 ( .ip(n10033), .op(n10038) );
  buf_1 U7246 ( .ip(n10034), .op(n10036) );
  buf_1 U7247 ( .ip(n10034), .op(n10039) );
  nand2_1 U7248 ( .ip1(n5552), .ip2(n5551), .op(n5553) );
  nor2_1 U7249 ( .ip1(n7583), .ip2(n9900), .op(n7585) );
  nand2_1 U7250 ( .ip1(n5281), .ip2(n11692), .op(n11654) );
  nand2_1 U7251 ( .ip1(n11652), .ip2(n11691), .op(n11655) );
  nand2_1 U7252 ( .ip1(n7500), .ip2(n11692), .op(n9837) );
  nand2_1 U7253 ( .ip1(n7500), .ip2(n11693), .op(n9896) );
  nor2_1 U7254 ( .ip1(n9900), .ip2(n9899), .op(n9901) );
  nand2_1 U7255 ( .ip1(n7500), .ip2(n11568), .op(n9817) );
  nand2_1 U7256 ( .ip1(n9852), .ip2(n9841), .op(n9843) );
  nand2_1 U7257 ( .ip1(n11573), .ip2(n9841), .op(n9842) );
  and2_1 U7258 ( .ip1(n5868), .ip2(n9335), .op(n9838) );
  nor2_1 U7259 ( .ip1(n9909), .ip2(n11616), .op(n11606) );
  inv_1 U7260 ( .ip(n7612), .op(n7573) );
  or2_1 U7261 ( .ip1(n11476), .ip2(n11475), .op(n11506) );
  nor2_1 U7262 ( .ip1(i_apb_U_DW_apb_ahbsif_use_saved_c), .ip2(n11368), .op(
        n11476) );
  nor3_1 U7263 ( .ip1(n10107), .ip2(n10110), .ip3(n6596), .op(n11466) );
  inv_1 U7264 ( .ip(n9374), .op(n6574) );
  nand2_1 U7265 ( .ip1(n10107), .ip2(n6584), .op(n10011) );
  inv_1 U7266 ( .ip(n10011), .op(n10018) );
  nand2_1 U7267 ( .ip1(n10021), .ip2(n10024), .op(n9897) );
  inv_1 U7268 ( .ip(n11367), .op(n9377) );
  nand2_1 U7269 ( .ip1(n9196), .ip2(n6550), .op(n6555) );
  nand2_1 U7270 ( .ip1(n5648), .ip2(n5647), .op(n7629) );
  nor2_1 U7271 ( .ip1(n7629), .ip2(n7628), .op(n7630) );
  inv_1 U7272 ( .ip(n11607), .op(i_ssi_ssi_rxu_intr_n) );
  inv_1 U7273 ( .ip(n11748), .op(i_ssi_ssi_oe_n) );
  inv_1 U7274 ( .ip(n11724), .op(i_ssi_ss_0_n) );
  nand3_1 U7275 ( .ip1(n9194), .ip2(n9193), .ip3(n9192), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hresp[1]) );
  inv_1 U7276 ( .ip(PRESETn_presetn), .op(n11766) );
  mux2_1 U7277 ( .ip1(i_apb_pwdata_int[0]), .ip2(n5282), .s(n9817), .op(n4637)
         );
  mux2_1 U7278 ( .ip1(i_apb_pwdata_int[10]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[10]), .s(n9896), .op(n4616) );
  mux2_1 U7279 ( .ip1(i_apb_pwdata_int[14]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[14]), .s(n9896), .op(n4612) );
  mux2_1 U7280 ( .ip1(i_apb_pwdata_int[1]), .ip2(n5395), .s(n9896), .op(n4609)
         );
  mux2_1 U7281 ( .ip1(i_apb_pwdata_int[15]), .ip2(n5394), .s(n9896), .op(n4611) );
  mux2_1 U7282 ( .ip1(n5398), .ip2(i_apb_pwdata_int[1]), .s(n9844), .op(n4589)
         );
  mux2_1 U7283 ( .ip1(i_ssi_dfs[0]), .ip2(i_apb_pwdata_int[0]), .s(n9844), 
        .op(n4588) );
  mux2_1 U7284 ( .ip1(i_apb_pwdata_int[11]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[11]), .s(n9896), .op(n4615) );
  mux2_1 U7285 ( .ip1(n10310), .ip2(i_apb_pwdata_int[3]), .s(n9901), .op(n4631) );
  nand2_1 U7286 ( .ip1(n6194), .ip2(n6171), .op(n6198) );
  nor2_1 U7287 ( .ip1(n10542), .ip2(n9087), .op(n4200) );
  nor2_1 U7288 ( .ip1(n10547), .ip2(n10334), .op(n5678) );
  nor2_1 U7289 ( .ip1(n10354), .ip2(n10353), .op(n10359) );
  inv_1 U7290 ( .ip(n10356), .op(n10353) );
  nor2_1 U7291 ( .ip1(n10435), .ip2(n10419), .op(i_ssi_U_sclkgen_N55) );
  mux2_1 U7292 ( .ip1(n9394), .ip2(i_i2c_U_DW_apb_i2c_tx_shift_data_sda_prev_r), .s(n10061), .op(n4941) );
  nand2_1 U7293 ( .ip1(n6169), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[13]), .op(n6173) );
  mux2_1 U7294 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[4]), .ip2(n9719), 
        .s(n6208), .op(n4406) );
  nand2_1 U7295 ( .ip1(n6210), .ip2(n6209), .op(n4407) );
  nand2_1 U7296 ( .ip1(n6207), .ip2(n6206), .op(n6210) );
  mux2_1 U7297 ( .ip1(i_ssi_baudr[4]), .ip2(i_apb_pwdata_int[4]), .s(n9901), 
        .op(n4630) );
  mux2_1 U7298 ( .ip1(i_ssi_baudr[12]), .ip2(i_apb_pwdata_int[12]), .s(n9901), 
        .op(n4622) );
  mux2_1 U7299 ( .ip1(n5257), .ip2(i_apb_pwdata_int[10]), .s(n9901), .op(n4624) );
  nor2_1 U7300 ( .ip1(i_ssi_U_fifo_U_tx_fifo_N37), .ip2(n10194), .op(n10195)
         );
  inv_1 U7301 ( .ip(n11244), .op(n6615) );
  inv_1 U7302 ( .ip(n9953), .op(n9954) );
  and2_1 U7303 ( .ip1(n9079), .ip2(n11166), .op(n9080) );
  nand2_1 U7304 ( .ip1(n11151), .ip2(n9077), .op(n9078) );
  nor3_1 U7305 ( .ip1(n6977), .ip2(n8576), .ip3(n6976), .op(
        i_ssi_U_fifo_U_tx_fifo_N45) );
  nor2_1 U7306 ( .ip1(n6650), .ip2(n6972), .op(i_ssi_U_fifo_U_tx_fifo_N38) );
  and2_1 U7307 ( .ip1(i_i2c_fifo_rst_n), .ip2(n6989), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N49) );
  nor3_1 U7308 ( .ip1(n7059), .ip2(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N37), 
        .ip3(n7058), .op(n7060) );
  nor2_1 U7309 ( .ip1(n11258), .ip2(n7053), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N49) );
  nor2_1 U7310 ( .ip1(n6988), .ip2(n11207), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N47) );
  mux2_1 U7311 ( .ip1(i_apb_pwdata_int[12]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[12]), .s(n9896), .op(n4614) );
  mux2_1 U7312 ( .ip1(n10385), .ip2(i_apb_pwdata_int[1]), .s(n9901), .op(n4633) );
  nand2_1 U7313 ( .ip1(n5233), .ip2(i_ssi_fsm_multi_mst), .op(n5686) );
  nand2_1 U7314 ( .ip1(n5685), .ip2(i_ssi_fsm_multi_mst), .op(n5687) );
  mux2_1 U7315 ( .ip1(n10384), .ip2(i_apb_pwdata_int[2]), .s(n9901), .op(n4632) );
  inv_1 U7316 ( .ip(n10444), .op(n10446) );
  inv_1 U7317 ( .ip(n10434), .op(n10436) );
  inv_1 U7318 ( .ip(n10462), .op(n10464) );
  inv_1 U7319 ( .ip(n10466), .op(n10463) );
  inv_1 U7320 ( .ip(i_ssi_U_sclkgen_ssi_cnt[10]), .op(n10459) );
  inv_1 U7321 ( .ip(n10456), .op(n10458) );
  inv_1 U7322 ( .ip(n10460), .op(n10457) );
  inv_1 U7323 ( .ip(n10450), .op(n10452) );
  mux2_1 U7324 ( .ip1(i_apb_pwdata_int[14]), .ip2(i_ssi_cfs[2]), .s(n9837), 
        .op(n4601) );
  nor2_1 U7325 ( .ip1(n10275), .ip2(n6460), .op(n4159) );
  inv_1 U7326 ( .ip(n6540), .op(i_i2c_U_DW_apb_i2c_toggle_tx_abrt) );
  mux2_1 U7327 ( .ip1(i_ssi_baudr[6]), .ip2(i_apb_pwdata_int[6]), .s(n9901), 
        .op(n4628) );
  mux2_1 U7328 ( .ip1(i_ssi_baudr[5]), .ip2(i_apb_pwdata_int[5]), .s(n9901), 
        .op(n4629) );
  mux2_1 U7329 ( .ip1(i_ssi_baudr[14]), .ip2(i_apb_pwdata_int[14]), .s(n9901), 
        .op(n4620) );
  inv_1 U7330 ( .ip(n10468), .op(n10471) );
  xor2_1 U7331 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[3]), .ip2(n9944), .op(n6458) );
  nor2_1 U7332 ( .ip1(n10275), .ip2(n6654), .op(n4164) );
  nor2_1 U7333 ( .ip1(n10275), .ip2(n6970), .op(n4165) );
  nor3_1 U7334 ( .ip1(n11116), .ip2(n10569), .ip3(n11158), .op(n10573) );
  nor2_1 U7335 ( .ip1(n8573), .ip2(n8572), .op(n4171) );
  and2_1 U7336 ( .ip1(n8571), .ip2(n8570), .op(n8572) );
  nand2_1 U7337 ( .ip1(n5279), .ip2(i_ssi_U_mstfsm_spi0_control), .op(n10241)
         );
  and2_1 U7338 ( .ip1(n10233), .ip2(n6309), .op(n4198) );
  or2_1 U7339 ( .ip1(n9082), .ip2(n6305), .op(n6308) );
  nand2_1 U7340 ( .ip1(n6987), .ip2(n5400), .op(n4201) );
  nor2_1 U7341 ( .ip1(n10480), .ip2(n9367), .op(n4206) );
  inv_1 U7342 ( .ip(n10481), .op(n10477) );
  nor2_1 U7343 ( .ip1(n9191), .ip2(n10480), .op(n4210) );
  mux2_2 U7344 ( .ip1(n6595), .ip2(i_apb_psel_en), .s(n10106), .op(n4212) );
  nor3_1 U7345 ( .ip1(n9643), .ip2(n9642), .ip3(n9645), .op(n9644) );
  mux2_1 U7346 ( .ip1(i_i2c_prdata[30]), .ip2(i_i2c_iprdata[30]), .s(n7435), 
        .op(n4691) );
  mux2_1 U7347 ( .ip1(i_i2c_prdata[28]), .ip2(i_i2c_iprdata[29]), .s(n7435), 
        .op(n4689) );
  mux2_1 U7348 ( .ip1(i_i2c_prdata[26]), .ip2(i_i2c_iprdata[26]), .s(n7435), 
        .op(n4687) );
  mux2_1 U7349 ( .ip1(i_i2c_prdata[25]), .ip2(i_i2c_iprdata[25]), .s(n7435), 
        .op(n4686) );
  mux2_1 U7350 ( .ip1(i_i2c_prdata[12]), .ip2(i_i2c_iprdata[12]), .s(n7435), 
        .op(n4673) );
  mux2_1 U7351 ( .ip1(i_i2c_prdata[11]), .ip2(i_i2c_iprdata[11]), .s(n7435), 
        .op(n4672) );
  mux2_1 U7352 ( .ip1(i_i2c_prdata[10]), .ip2(i_i2c_iprdata[10]), .s(n7435), 
        .op(n4671) );
  mux2_1 U7353 ( .ip1(i_i2c_prdata[8]), .ip2(i_i2c_iprdata[8]), .s(n7435), 
        .op(n4669) );
  mux2_1 U7354 ( .ip1(i_i2c_prdata[7]), .ip2(i_i2c_iprdata[7]), .s(n7435), 
        .op(n4668) );
  mux2_1 U7355 ( .ip1(i_i2c_prdata[6]), .ip2(i_i2c_iprdata[6]), .s(n7435), 
        .op(n4667) );
  mux2_1 U7356 ( .ip1(i_i2c_prdata[5]), .ip2(i_i2c_iprdata[5]), .s(n7435), 
        .op(n4666) );
  mux2_1 U7357 ( .ip1(i_i2c_prdata[4]), .ip2(i_i2c_iprdata[4]), .s(n7435), 
        .op(n4665) );
  mux2_1 U7358 ( .ip1(i_i2c_prdata[3]), .ip2(i_i2c_iprdata[3]), .s(n7435), 
        .op(n4664) );
  mux2_1 U7359 ( .ip1(i_i2c_prdata[2]), .ip2(i_i2c_iprdata[2]), .s(n7435), 
        .op(n4663) );
  mux2_1 U7360 ( .ip1(i_i2c_prdata[1]), .ip2(i_i2c_iprdata[1]), .s(n7435), 
        .op(n4662) );
  mux2_1 U7361 ( .ip1(i_i2c_prdata[0]), .ip2(i_i2c_iprdata[0]), .s(n7435), 
        .op(n4661) );
  or2_1 U7362 ( .ip1(n8500), .ip2(n8499), .op(n8501) );
  or2_1 U7363 ( .ip1(n8506), .ip2(n8505), .op(n8507) );
  or2_1 U7364 ( .ip1(n8518), .ip2(n8517), .op(n8519) );
  or2_1 U7365 ( .ip1(n8512), .ip2(n8511), .op(n8513) );
  nor3_1 U7366 ( .ip1(n11099), .ip2(n7919), .ip3(n10002), .op(
        i_i2c_U_DW_apb_i2c_tx_shift_mst_slv_ack_ext) );
  nor2_1 U7367 ( .ip1(n11041), .ip2(n8879), .op(n5154) );
  xnor2_1 U7368 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[15]), .ip2(
        n11040), .op(n8879) );
  xnor2_1 U7369 ( .ip1(n10631), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[15]), .op(n8388) );
  nor2_1 U7370 ( .ip1(n10994), .ip2(n9055), .op(n5138) );
  xnor2_1 U7371 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[15]), .ip2(
        n10268), .op(n9055) );
  nor2_1 U7372 ( .ip1(n9416), .ip2(n6470), .op(n9421) );
  nor2_1 U7373 ( .ip1(n9428), .ip2(n6470), .op(n9434) );
  nor2_1 U7374 ( .ip1(n9734), .ip2(n6470), .op(n9739) );
  mux2_1 U7375 ( .ip1(n9403), .ip2(n9402), .s(i_i2c_tx_abrt_source[10]), .op(
        n5209) );
  nor2_1 U7376 ( .ip1(n9667), .ip2(n9662), .op(n9663) );
  nor2_1 U7377 ( .ip1(n9699), .ip2(n9737), .op(n9700) );
  xnor2_1 U7378 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[15]), .ip2(
        n10678), .op(n8724) );
  xnor2_1 U7379 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[15]), .ip2(
        n10956), .op(n8210) );
  nand3_1 U7380 ( .ip1(n9636), .ip2(n9653), .ip3(n9609), .op(n9610) );
  nor3_1 U7381 ( .ip1(n9724), .ip2(n9723), .ip3(n9722), .op(n9726) );
  mux2_1 U7382 ( .ip1(i_i2c_slv_debug_cstate[1]), .ip2(i_i2c_slv_rx_2addr), 
        .s(n9399), .op(n5231) );
  nand2_1 U7383 ( .ip1(n9654), .ip2(n9653), .op(n9655) );
  nor2_1 U7384 ( .ip1(n9636), .ip2(n9635), .op(n9637) );
  nor2_1 U7385 ( .ip1(n9634), .ip2(n9633), .op(n9635) );
  nor2_1 U7386 ( .ip1(n9567), .ip2(n9633), .op(n9568) );
  nand3_1 U7387 ( .ip1(n11350), .ip2(n11349), .ip3(n11348), .op(n11353) );
  nand3_1 U7388 ( .ip1(n11344), .ip2(n11349), .ip3(n11348), .op(n11347) );
  nor4_1 U7389 ( .ip1(n8544), .ip2(n8543), .ip3(n8542), .ip4(n8550), .op(n8545) );
  nor2_1 U7390 ( .ip1(n7508), .ip2(n11144), .op(n5096) );
  and2_1 U7391 ( .ip1(n7507), .ip2(n7506), .op(n7508) );
  nor3_1 U7392 ( .ip1(n7050), .ip2(n7505), .ip3(n11144), .op(n5103) );
  nor2_1 U7393 ( .ip1(n6848), .ip2(n7069), .op(n11772) );
  nor2_1 U7394 ( .ip1(n6844), .ip2(n8266), .op(n6848) );
  inv_1 U7395 ( .ip(n6843), .op(n6844) );
  nand3_1 U7396 ( .ip1(n8346), .ip2(n8345), .ip3(n8546), .op(
        i_i2c_U_DW_apb_i2c_tx_shift_N90) );
  and3_1 U7397 ( .ip1(n8343), .ip2(n8342), .ip3(n8341), .op(n8345) );
  nand2_1 U7398 ( .ip1(n6901), .ip2(n6840), .op(n5206) );
  nor2_1 U7399 ( .ip1(n8373), .ip2(n8372), .op(i_i2c_U_DW_apb_i2c_mstfsm_N74)
         );
  inv_1 U7400 ( .ip(n11045), .op(n8373) );
  nor2_1 U7401 ( .ip1(n11044), .ip2(n8372), .op(i_i2c_U_DW_apb_i2c_mstfsm_N73)
         );
  nand2_1 U7402 ( .ip1(n6466), .ip2(n6869), .op(i_i2c_U_DW_apb_i2c_mstfsm_N487) );
  nor2_1 U7403 ( .ip1(n11305), .ip2(n8372), .op(i_i2c_U_DW_apb_i2c_mstfsm_N75)
         );
  nor2_1 U7404 ( .ip1(n11305), .ip2(n11304), .op(n11308) );
  nor2_1 U7405 ( .ip1(n6837), .ip2(n10630), .op(n5200) );
  nor2_1 U7406 ( .ip1(i_i2c_scl_lcnt_cmplt), .ip2(n10589), .op(n6837) );
  nand2_1 U7407 ( .ip1(n6883), .ip2(n6876), .op(n5232) );
  nor2_1 U7408 ( .ip1(n10914), .ip2(n10913), .op(n10916) );
  nor2_1 U7409 ( .ip1(n10912), .ip2(n10911), .op(n10913) );
  nor2_1 U7410 ( .ip1(n7081), .ip2(n7080), .op(n4939) );
  nor2_1 U7411 ( .ip1(n7079), .ip2(n7078), .op(n7081) );
  nand2_1 U7412 ( .ip1(n8377), .ip2(n9920), .op(n4245) );
  nand2_1 U7413 ( .ip1(n9924), .ip2(n9923), .op(n9925) );
  nand2_1 U7414 ( .ip1(n9919), .ip2(n9918), .op(n9924) );
  nand2_1 U7415 ( .ip1(n4645), .ip2(n9922), .op(n9923) );
  nand2_1 U7416 ( .ip1(n11624), .ip2(n11623), .op(n11626) );
  nand2_1 U7417 ( .ip1(n11622), .ip2(n11621), .op(n11623) );
  nand2_1 U7418 ( .ip1(n9920), .ip2(n9913), .op(n9914) );
  nor2_1 U7419 ( .ip1(n5233), .ip2(n5372), .op(n11778) );
  mux2_1 U7420 ( .ip1(i_ssi_U_dff_rx_mem[112]), .ip2(i_ssi_rx_push_data[0]), 
        .s(n9370), .op(n4370) );
  mux2_1 U7421 ( .ip1(i_ssi_rx_push_data[0]), .ip2(i_ssi_U_dff_rx_mem[96]), 
        .s(n10050), .op(n4371) );
  mux2_1 U7422 ( .ip1(i_ssi_U_dff_rx_mem[80]), .ip2(i_ssi_rx_push_data[0]), 
        .s(n9371), .op(n4372) );
  mux2_1 U7423 ( .ip1(i_ssi_U_dff_rx_mem[64]), .ip2(i_ssi_rx_push_data[0]), 
        .s(n5274), .op(n4373) );
  mux2_1 U7424 ( .ip1(i_ssi_U_dff_rx_mem[48]), .ip2(i_ssi_rx_push_data[0]), 
        .s(n9369), .op(n4374) );
  mux2_1 U7425 ( .ip1(i_ssi_rx_push_data[0]), .ip2(i_ssi_U_dff_rx_mem[32]), 
        .s(n10049), .op(n4375) );
  mux2_1 U7426 ( .ip1(i_ssi_rx_push_data[0]), .ip2(i_ssi_U_dff_rx_mem[16]), 
        .s(n9697), .op(n4376) );
  mux2_1 U7427 ( .ip1(i_ssi_U_dff_rx_mem[0]), .ip2(i_ssi_rx_push_data[0]), .s(
        n5275), .op(n4377) );
  mux2_1 U7428 ( .ip1(i_ssi_U_dff_rx_mem[127]), .ip2(i_ssi_rx_push_data[15]), 
        .s(n9370), .op(n4250) );
  mux2_1 U7429 ( .ip1(i_ssi_rx_push_data[15]), .ip2(i_ssi_U_dff_rx_mem[111]), 
        .s(n10050), .op(n4251) );
  mux2_1 U7430 ( .ip1(i_ssi_U_dff_rx_mem[95]), .ip2(i_ssi_rx_push_data[15]), 
        .s(n9371), .op(n4252) );
  mux2_1 U7431 ( .ip1(i_ssi_U_dff_rx_mem[79]), .ip2(i_ssi_rx_push_data[15]), 
        .s(n5274), .op(n4253) );
  mux2_1 U7432 ( .ip1(i_ssi_U_dff_rx_mem[63]), .ip2(i_ssi_rx_push_data[15]), 
        .s(n9369), .op(n4254) );
  mux2_1 U7433 ( .ip1(i_ssi_rx_push_data[15]), .ip2(i_ssi_U_dff_rx_mem[47]), 
        .s(n10049), .op(n4255) );
  mux2_1 U7434 ( .ip1(i_ssi_rx_push_data[15]), .ip2(i_ssi_U_dff_rx_mem[31]), 
        .s(n9697), .op(n4256) );
  mux2_1 U7435 ( .ip1(i_ssi_U_dff_rx_mem[15]), .ip2(i_ssi_rx_push_data[15]), 
        .s(n5275), .op(n4257) );
  mux2_1 U7436 ( .ip1(i_ssi_U_dff_rx_mem[126]), .ip2(i_ssi_rx_push_data[14]), 
        .s(n9370), .op(n4258) );
  mux2_1 U7437 ( .ip1(i_ssi_rx_push_data[14]), .ip2(i_ssi_U_dff_rx_mem[110]), 
        .s(n10050), .op(n4259) );
  mux2_1 U7438 ( .ip1(i_ssi_U_dff_rx_mem[94]), .ip2(i_ssi_rx_push_data[14]), 
        .s(n9371), .op(n4260) );
  mux2_1 U7439 ( .ip1(i_ssi_U_dff_rx_mem[78]), .ip2(i_ssi_rx_push_data[14]), 
        .s(n5274), .op(n4261) );
  mux2_1 U7440 ( .ip1(i_ssi_U_dff_rx_mem[62]), .ip2(i_ssi_rx_push_data[14]), 
        .s(n9369), .op(n4262) );
  mux2_1 U7441 ( .ip1(i_ssi_rx_push_data[14]), .ip2(i_ssi_U_dff_rx_mem[46]), 
        .s(n10049), .op(n4263) );
  mux2_1 U7442 ( .ip1(i_ssi_rx_push_data[14]), .ip2(i_ssi_U_dff_rx_mem[30]), 
        .s(n9697), .op(n4264) );
  mux2_1 U7443 ( .ip1(i_ssi_U_dff_rx_mem[14]), .ip2(i_ssi_rx_push_data[14]), 
        .s(n5275), .op(n4265) );
  mux2_1 U7444 ( .ip1(i_ssi_U_dff_rx_mem[125]), .ip2(i_ssi_rx_push_data[13]), 
        .s(n9370), .op(n4266) );
  mux2_1 U7445 ( .ip1(i_ssi_rx_push_data[13]), .ip2(i_ssi_U_dff_rx_mem[109]), 
        .s(n10050), .op(n4267) );
  mux2_1 U7446 ( .ip1(i_ssi_U_dff_rx_mem[93]), .ip2(i_ssi_rx_push_data[13]), 
        .s(n9371), .op(n4268) );
  mux2_1 U7447 ( .ip1(i_ssi_U_dff_rx_mem[77]), .ip2(i_ssi_rx_push_data[13]), 
        .s(n5274), .op(n4269) );
  mux2_1 U7448 ( .ip1(i_ssi_U_dff_rx_mem[61]), .ip2(i_ssi_rx_push_data[13]), 
        .s(n9369), .op(n4270) );
  mux2_1 U7449 ( .ip1(i_ssi_rx_push_data[13]), .ip2(i_ssi_U_dff_rx_mem[45]), 
        .s(n10049), .op(n4271) );
  mux2_1 U7450 ( .ip1(i_ssi_rx_push_data[13]), .ip2(i_ssi_U_dff_rx_mem[29]), 
        .s(n9697), .op(n4272) );
  mux2_1 U7451 ( .ip1(i_ssi_U_dff_rx_mem[13]), .ip2(i_ssi_rx_push_data[13]), 
        .s(n5275), .op(n4273) );
  mux2_1 U7452 ( .ip1(i_ssi_U_dff_rx_mem[124]), .ip2(i_ssi_rx_push_data[12]), 
        .s(n9370), .op(n4274) );
  mux2_1 U7453 ( .ip1(i_ssi_rx_push_data[12]), .ip2(i_ssi_U_dff_rx_mem[108]), 
        .s(n10050), .op(n4275) );
  mux2_1 U7454 ( .ip1(i_ssi_U_dff_rx_mem[92]), .ip2(i_ssi_rx_push_data[12]), 
        .s(n9371), .op(n4276) );
  mux2_1 U7455 ( .ip1(i_ssi_U_dff_rx_mem[76]), .ip2(i_ssi_rx_push_data[12]), 
        .s(n5274), .op(n4277) );
  mux2_1 U7456 ( .ip1(i_ssi_U_dff_rx_mem[60]), .ip2(i_ssi_rx_push_data[12]), 
        .s(n9369), .op(n4278) );
  mux2_1 U7457 ( .ip1(i_ssi_rx_push_data[12]), .ip2(i_ssi_U_dff_rx_mem[44]), 
        .s(n10049), .op(n4279) );
  mux2_1 U7458 ( .ip1(i_ssi_rx_push_data[12]), .ip2(i_ssi_U_dff_rx_mem[28]), 
        .s(n9697), .op(n4280) );
  mux2_1 U7459 ( .ip1(i_ssi_U_dff_rx_mem[12]), .ip2(i_ssi_rx_push_data[12]), 
        .s(n5275), .op(n4281) );
  mux2_1 U7460 ( .ip1(i_ssi_U_dff_rx_mem[123]), .ip2(i_ssi_rx_push_data[11]), 
        .s(n9370), .op(n4282) );
  mux2_1 U7461 ( .ip1(i_ssi_rx_push_data[11]), .ip2(i_ssi_U_dff_rx_mem[107]), 
        .s(n10050), .op(n4283) );
  mux2_1 U7462 ( .ip1(i_ssi_U_dff_rx_mem[91]), .ip2(i_ssi_rx_push_data[11]), 
        .s(n9371), .op(n4284) );
  mux2_1 U7463 ( .ip1(i_ssi_U_dff_rx_mem[75]), .ip2(i_ssi_rx_push_data[11]), 
        .s(n5274), .op(n4285) );
  mux2_1 U7464 ( .ip1(i_ssi_U_dff_rx_mem[59]), .ip2(i_ssi_rx_push_data[11]), 
        .s(n9369), .op(n4286) );
  mux2_1 U7465 ( .ip1(i_ssi_rx_push_data[11]), .ip2(i_ssi_U_dff_rx_mem[43]), 
        .s(n10049), .op(n4287) );
  mux2_1 U7466 ( .ip1(i_ssi_rx_push_data[11]), .ip2(i_ssi_U_dff_rx_mem[27]), 
        .s(n9697), .op(n4288) );
  mux2_1 U7467 ( .ip1(i_ssi_U_dff_rx_mem[11]), .ip2(i_ssi_rx_push_data[11]), 
        .s(n5275), .op(n4289) );
  mux2_1 U7468 ( .ip1(i_ssi_U_dff_rx_mem[122]), .ip2(i_ssi_rx_push_data[10]), 
        .s(n9370), .op(n4290) );
  mux2_1 U7469 ( .ip1(i_ssi_rx_push_data[10]), .ip2(i_ssi_U_dff_rx_mem[106]), 
        .s(n10050), .op(n4291) );
  mux2_1 U7470 ( .ip1(i_ssi_U_dff_rx_mem[90]), .ip2(i_ssi_rx_push_data[10]), 
        .s(n9371), .op(n4292) );
  mux2_1 U7471 ( .ip1(i_ssi_U_dff_rx_mem[74]), .ip2(i_ssi_rx_push_data[10]), 
        .s(n5274), .op(n4293) );
  mux2_1 U7472 ( .ip1(i_ssi_U_dff_rx_mem[58]), .ip2(i_ssi_rx_push_data[10]), 
        .s(n9369), .op(n4294) );
  mux2_1 U7473 ( .ip1(i_ssi_rx_push_data[10]), .ip2(i_ssi_U_dff_rx_mem[42]), 
        .s(n10049), .op(n4295) );
  mux2_1 U7474 ( .ip1(i_ssi_rx_push_data[10]), .ip2(i_ssi_U_dff_rx_mem[26]), 
        .s(n9697), .op(n4296) );
  mux2_1 U7475 ( .ip1(i_ssi_U_dff_rx_mem[10]), .ip2(i_ssi_rx_push_data[10]), 
        .s(n5275), .op(n4297) );
  mux2_1 U7476 ( .ip1(i_ssi_U_dff_rx_mem[121]), .ip2(i_ssi_rx_push_data[9]), 
        .s(n9370), .op(n4298) );
  mux2_1 U7477 ( .ip1(i_ssi_rx_push_data[9]), .ip2(i_ssi_U_dff_rx_mem[105]), 
        .s(n10050), .op(n4299) );
  mux2_1 U7478 ( .ip1(i_ssi_U_dff_rx_mem[89]), .ip2(i_ssi_rx_push_data[9]), 
        .s(n9371), .op(n4300) );
  mux2_1 U7479 ( .ip1(i_ssi_U_dff_rx_mem[73]), .ip2(i_ssi_rx_push_data[9]), 
        .s(n5274), .op(n4301) );
  mux2_1 U7480 ( .ip1(i_ssi_U_dff_rx_mem[57]), .ip2(i_ssi_rx_push_data[9]), 
        .s(n9369), .op(n4302) );
  mux2_1 U7481 ( .ip1(i_ssi_rx_push_data[9]), .ip2(i_ssi_U_dff_rx_mem[41]), 
        .s(n10049), .op(n4303) );
  mux2_1 U7482 ( .ip1(i_ssi_rx_push_data[9]), .ip2(i_ssi_U_dff_rx_mem[25]), 
        .s(n9697), .op(n4304) );
  mux2_1 U7483 ( .ip1(i_ssi_U_dff_rx_mem[9]), .ip2(i_ssi_rx_push_data[9]), .s(
        n5275), .op(n4305) );
  mux2_1 U7484 ( .ip1(i_ssi_U_dff_rx_mem[120]), .ip2(i_ssi_rx_push_data[8]), 
        .s(n9370), .op(n4306) );
  mux2_1 U7485 ( .ip1(i_ssi_rx_push_data[8]), .ip2(i_ssi_U_dff_rx_mem[104]), 
        .s(n10050), .op(n4307) );
  mux2_1 U7486 ( .ip1(i_ssi_U_dff_rx_mem[88]), .ip2(i_ssi_rx_push_data[8]), 
        .s(n9371), .op(n4308) );
  mux2_1 U7487 ( .ip1(i_ssi_U_dff_rx_mem[72]), .ip2(i_ssi_rx_push_data[8]), 
        .s(n5274), .op(n4309) );
  mux2_1 U7488 ( .ip1(i_ssi_U_dff_rx_mem[56]), .ip2(i_ssi_rx_push_data[8]), 
        .s(n9369), .op(n4310) );
  mux2_1 U7489 ( .ip1(i_ssi_rx_push_data[8]), .ip2(i_ssi_U_dff_rx_mem[40]), 
        .s(n10049), .op(n4311) );
  mux2_1 U7490 ( .ip1(i_ssi_rx_push_data[8]), .ip2(i_ssi_U_dff_rx_mem[24]), 
        .s(n9697), .op(n4312) );
  mux2_1 U7491 ( .ip1(i_ssi_U_dff_rx_mem[8]), .ip2(i_ssi_rx_push_data[8]), .s(
        n5275), .op(n4313) );
  mux2_1 U7492 ( .ip1(i_ssi_U_dff_rx_mem[119]), .ip2(i_ssi_rx_push_data[7]), 
        .s(n9370), .op(n4314) );
  mux2_1 U7493 ( .ip1(i_ssi_rx_push_data[7]), .ip2(i_ssi_U_dff_rx_mem[103]), 
        .s(n10050), .op(n4315) );
  mux2_1 U7494 ( .ip1(i_ssi_U_dff_rx_mem[87]), .ip2(i_ssi_rx_push_data[7]), 
        .s(n9371), .op(n4316) );
  mux2_1 U7495 ( .ip1(i_ssi_U_dff_rx_mem[71]), .ip2(i_ssi_rx_push_data[7]), 
        .s(n5274), .op(n4317) );
  mux2_1 U7496 ( .ip1(i_ssi_U_dff_rx_mem[55]), .ip2(i_ssi_rx_push_data[7]), 
        .s(n9369), .op(n4318) );
  mux2_1 U7497 ( .ip1(i_ssi_rx_push_data[7]), .ip2(i_ssi_U_dff_rx_mem[39]), 
        .s(n10049), .op(n4319) );
  mux2_1 U7498 ( .ip1(i_ssi_rx_push_data[7]), .ip2(i_ssi_U_dff_rx_mem[23]), 
        .s(n9697), .op(n4320) );
  mux2_1 U7499 ( .ip1(i_ssi_U_dff_rx_mem[7]), .ip2(i_ssi_rx_push_data[7]), .s(
        n5275), .op(n4321) );
  mux2_1 U7500 ( .ip1(i_ssi_U_dff_rx_mem[118]), .ip2(i_ssi_rx_push_data[6]), 
        .s(n9370), .op(n4322) );
  mux2_1 U7501 ( .ip1(i_ssi_rx_push_data[6]), .ip2(i_ssi_U_dff_rx_mem[102]), 
        .s(n10050), .op(n4323) );
  mux2_1 U7502 ( .ip1(i_ssi_U_dff_rx_mem[86]), .ip2(i_ssi_rx_push_data[6]), 
        .s(n9371), .op(n4324) );
  mux2_1 U7503 ( .ip1(i_ssi_U_dff_rx_mem[70]), .ip2(i_ssi_rx_push_data[6]), 
        .s(n5274), .op(n4325) );
  mux2_1 U7504 ( .ip1(i_ssi_U_dff_rx_mem[54]), .ip2(i_ssi_rx_push_data[6]), 
        .s(n9369), .op(n4326) );
  mux2_1 U7505 ( .ip1(i_ssi_rx_push_data[6]), .ip2(i_ssi_U_dff_rx_mem[38]), 
        .s(n10049), .op(n4327) );
  mux2_1 U7506 ( .ip1(i_ssi_rx_push_data[6]), .ip2(i_ssi_U_dff_rx_mem[22]), 
        .s(n9697), .op(n4328) );
  mux2_1 U7507 ( .ip1(i_ssi_U_dff_rx_mem[6]), .ip2(i_ssi_rx_push_data[6]), .s(
        n5275), .op(n4329) );
  mux2_1 U7508 ( .ip1(i_ssi_U_dff_rx_mem[117]), .ip2(i_ssi_rx_push_data[5]), 
        .s(n9370), .op(n4330) );
  mux2_1 U7509 ( .ip1(i_ssi_rx_push_data[5]), .ip2(i_ssi_U_dff_rx_mem[101]), 
        .s(n10050), .op(n4331) );
  mux2_1 U7510 ( .ip1(i_ssi_U_dff_rx_mem[85]), .ip2(i_ssi_rx_push_data[5]), 
        .s(n9371), .op(n4332) );
  mux2_1 U7511 ( .ip1(i_ssi_U_dff_rx_mem[69]), .ip2(i_ssi_rx_push_data[5]), 
        .s(n5274), .op(n4333) );
  mux2_1 U7512 ( .ip1(i_ssi_U_dff_rx_mem[53]), .ip2(i_ssi_rx_push_data[5]), 
        .s(n9369), .op(n4334) );
  mux2_1 U7513 ( .ip1(i_ssi_rx_push_data[5]), .ip2(i_ssi_U_dff_rx_mem[37]), 
        .s(n10049), .op(n4335) );
  mux2_1 U7514 ( .ip1(i_ssi_rx_push_data[5]), .ip2(i_ssi_U_dff_rx_mem[21]), 
        .s(n9697), .op(n4336) );
  mux2_1 U7515 ( .ip1(i_ssi_U_dff_rx_mem[5]), .ip2(i_ssi_rx_push_data[5]), .s(
        n5275), .op(n4337) );
  mux2_1 U7516 ( .ip1(i_ssi_U_dff_rx_mem[116]), .ip2(i_ssi_rx_push_data[4]), 
        .s(n9370), .op(n4338) );
  mux2_1 U7517 ( .ip1(i_ssi_rx_push_data[4]), .ip2(i_ssi_U_dff_rx_mem[100]), 
        .s(n10050), .op(n4339) );
  mux2_1 U7518 ( .ip1(i_ssi_U_dff_rx_mem[84]), .ip2(i_ssi_rx_push_data[4]), 
        .s(n9371), .op(n4340) );
  mux2_1 U7519 ( .ip1(i_ssi_U_dff_rx_mem[68]), .ip2(i_ssi_rx_push_data[4]), 
        .s(n5274), .op(n4341) );
  mux2_1 U7520 ( .ip1(i_ssi_U_dff_rx_mem[52]), .ip2(i_ssi_rx_push_data[4]), 
        .s(n9369), .op(n4342) );
  mux2_1 U7521 ( .ip1(i_ssi_rx_push_data[4]), .ip2(i_ssi_U_dff_rx_mem[36]), 
        .s(n10049), .op(n4343) );
  mux2_1 U7522 ( .ip1(i_ssi_rx_push_data[4]), .ip2(i_ssi_U_dff_rx_mem[20]), 
        .s(n9697), .op(n4344) );
  mux2_1 U7523 ( .ip1(i_ssi_U_dff_rx_mem[4]), .ip2(i_ssi_rx_push_data[4]), .s(
        n5275), .op(n4345) );
  mux2_1 U7524 ( .ip1(i_ssi_U_dff_rx_mem[115]), .ip2(i_ssi_rx_push_data[3]), 
        .s(n9370), .op(n4346) );
  mux2_1 U7525 ( .ip1(i_ssi_rx_push_data[3]), .ip2(i_ssi_U_dff_rx_mem[99]), 
        .s(n10050), .op(n4347) );
  mux2_1 U7526 ( .ip1(i_ssi_U_dff_rx_mem[83]), .ip2(i_ssi_rx_push_data[3]), 
        .s(n9371), .op(n4348) );
  mux2_1 U7527 ( .ip1(i_ssi_U_dff_rx_mem[67]), .ip2(i_ssi_rx_push_data[3]), 
        .s(n5274), .op(n4349) );
  mux2_1 U7528 ( .ip1(i_ssi_U_dff_rx_mem[51]), .ip2(i_ssi_rx_push_data[3]), 
        .s(n9369), .op(n4350) );
  mux2_1 U7529 ( .ip1(i_ssi_rx_push_data[3]), .ip2(i_ssi_U_dff_rx_mem[35]), 
        .s(n10049), .op(n4351) );
  mux2_1 U7530 ( .ip1(i_ssi_rx_push_data[3]), .ip2(i_ssi_U_dff_rx_mem[19]), 
        .s(n9697), .op(n4352) );
  mux2_1 U7531 ( .ip1(i_ssi_U_dff_rx_mem[3]), .ip2(i_ssi_rx_push_data[3]), .s(
        n5275), .op(n4353) );
  nor2_1 U7532 ( .ip1(n10068), .ip2(n10067), .op(n10069) );
  nor2_1 U7533 ( .ip1(n11558), .ip2(n10066), .op(n10067) );
  mux2_1 U7534 ( .ip1(i_ssi_U_dff_rx_mem[114]), .ip2(i_ssi_rx_push_data[2]), 
        .s(n9370), .op(n4354) );
  mux2_1 U7535 ( .ip1(i_ssi_rx_push_data[2]), .ip2(i_ssi_U_dff_rx_mem[98]), 
        .s(n10050), .op(n4355) );
  mux2_1 U7536 ( .ip1(i_ssi_U_dff_rx_mem[82]), .ip2(i_ssi_rx_push_data[2]), 
        .s(n9371), .op(n4356) );
  mux2_1 U7537 ( .ip1(i_ssi_U_dff_rx_mem[66]), .ip2(i_ssi_rx_push_data[2]), 
        .s(n5274), .op(n4357) );
  mux2_1 U7538 ( .ip1(i_ssi_U_dff_rx_mem[50]), .ip2(i_ssi_rx_push_data[2]), 
        .s(n9369), .op(n4358) );
  mux2_1 U7539 ( .ip1(i_ssi_rx_push_data[2]), .ip2(i_ssi_U_dff_rx_mem[34]), 
        .s(n10049), .op(n4359) );
  mux2_1 U7540 ( .ip1(i_ssi_rx_push_data[2]), .ip2(i_ssi_U_dff_rx_mem[18]), 
        .s(n9697), .op(n4360) );
  mux2_1 U7541 ( .ip1(i_ssi_U_dff_rx_mem[2]), .ip2(i_ssi_rx_push_data[2]), .s(
        n5275), .op(n4361) );
  mux2_1 U7542 ( .ip1(i_ssi_U_dff_rx_mem[113]), .ip2(i_ssi_rx_push_data[1]), 
        .s(n9370), .op(n4362) );
  mux2_1 U7543 ( .ip1(i_ssi_rx_push_data[1]), .ip2(i_ssi_U_dff_rx_mem[97]), 
        .s(n10050), .op(n4363) );
  mux2_1 U7544 ( .ip1(i_ssi_U_dff_rx_mem[81]), .ip2(i_ssi_rx_push_data[1]), 
        .s(n9371), .op(n4364) );
  mux2_1 U7545 ( .ip1(i_ssi_U_dff_rx_mem[65]), .ip2(i_ssi_rx_push_data[1]), 
        .s(n5274), .op(n4365) );
  mux2_1 U7546 ( .ip1(i_ssi_U_dff_rx_mem[49]), .ip2(i_ssi_rx_push_data[1]), 
        .s(n9369), .op(n4366) );
  mux2_1 U7547 ( .ip1(i_ssi_rx_push_data[1]), .ip2(i_ssi_U_dff_rx_mem[33]), 
        .s(n10049), .op(n4367) );
  mux2_1 U7548 ( .ip1(i_ssi_rx_push_data[1]), .ip2(i_ssi_U_dff_rx_mem[17]), 
        .s(n9697), .op(n4368) );
  mux2_1 U7549 ( .ip1(i_ssi_U_dff_rx_mem[1]), .ip2(i_ssi_rx_push_data[1]), .s(
        n5275), .op(n4369) );
  mux2_1 U7550 ( .ip1(n9682), .ip2(n11526), .s(i_ssi_U_regfile_rxflr[2]), .op(
        n4445) );
  mux2_1 U7551 ( .ip1(n9675), .ip2(n9679), .s(i_ssi_U_regfile_rxflr[0]), .op(
        n4447) );
  nand2_1 U7552 ( .ip1(n9674), .ip2(n9673), .op(n9675) );
  mux2_1 U7553 ( .ip1(i_ssi_txd), .ip2(i_ssi_rxd), .s(n9683), .op(n9691) );
  mux2_1 U7554 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[8]), .ip2(n9713), 
        .s(n9712), .op(n4402) );
  mux2_1 U7555 ( .ip1(n10343), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[15]), 
        .s(n10261), .op(n4412) );
  mux2_1 U7556 ( .ip1(n6189), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[14]), 
        .s(n10261), .op(n4413) );
  mux2_1 U7557 ( .ip1(n6164), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[13]), 
        .s(n10261), .op(n4414) );
  mux2_1 U7558 ( .ip1(n10255), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[12]), 
        .s(n10261), .op(n4415) );
  inv_1 U7559 ( .ip(n10254), .op(n10255) );
  mux2_1 U7560 ( .ip1(n6146), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[11]), 
        .s(n10261), .op(n4416) );
  mux2_1 U7561 ( .ip1(n6156), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[9]), 
        .s(n10261), .op(n4418) );
  inv_1 U7562 ( .ip(n9707), .op(n5791) );
  inv_1 U7563 ( .ip(n6101), .op(n5780) );
  mux2_1 U7564 ( .ip1(n10262), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[6]), 
        .s(n10261), .op(n4421) );
  inv_1 U7565 ( .ip(n10260), .op(n10262) );
  mux2_1 U7566 ( .ip1(n10259), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[5]), 
        .s(n10261), .op(n4422) );
  inv_1 U7567 ( .ip(n10258), .op(n10259) );
  mux2_1 U7568 ( .ip1(n10252), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[4]), 
        .s(n10261), .op(n4423) );
  inv_1 U7569 ( .ip(n10251), .op(n10252) );
  mux2_1 U7570 ( .ip1(n10249), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[3]), 
        .s(n10261), .op(n4424) );
  inv_1 U7571 ( .ip(n10248), .op(n10249) );
  mux2_1 U7572 ( .ip1(n10247), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[2]), 
        .s(n10261), .op(n4425) );
  inv_1 U7573 ( .ip(n10246), .op(n10247) );
  mux2_1 U7574 ( .ip1(n10277), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[1]), 
        .s(n10261), .op(n4426) );
  mux2_1 U7575 ( .ip1(n5458), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[0]), 
        .s(n10261), .op(n4427) );
  nand2_1 U7576 ( .ip1(n11517), .ip2(n11516), .op(n11521) );
  or2_1 U7577 ( .ip1(n11512), .ip2(n11514), .op(n11517) );
  mux2_1 U7578 ( .ip1(n9978), .ip2(n9977), .s(n11514), .op(n4452) );
  nand2_1 U7579 ( .ip1(n11512), .ip2(n9976), .op(n9977) );
  nand3_1 U7580 ( .ip1(n7092), .ip2(n9976), .ip3(n7091), .op(n4453) );
  mux2_1 U7581 ( .ip1(n9948), .ip2(n9947), .s(i_ssi_U_regfile_txflr[0]), .op(
        n4454) );
  mux2_1 U7582 ( .ip1(i_ssi_U_dff_tx_mem[127]), .ip2(i_apb_pwdata_int[15]), 
        .s(n10175), .op(n4456) );
  mux2_1 U7583 ( .ip1(i_ssi_U_dff_tx_mem[126]), .ip2(i_apb_pwdata_int[14]), 
        .s(n10175), .op(n4457) );
  mux2_1 U7584 ( .ip1(i_ssi_U_dff_tx_mem[125]), .ip2(i_apb_pwdata_int[13]), 
        .s(n10175), .op(n4458) );
  mux2_1 U7585 ( .ip1(i_ssi_U_dff_tx_mem[124]), .ip2(i_apb_pwdata_int[12]), 
        .s(n10175), .op(n4459) );
  mux2_1 U7586 ( .ip1(i_ssi_U_dff_tx_mem[123]), .ip2(i_apb_pwdata_int[11]), 
        .s(n10174), .op(n4460) );
  mux2_1 U7587 ( .ip1(i_ssi_U_dff_tx_mem[122]), .ip2(i_apb_pwdata_int[10]), 
        .s(n10174), .op(n4461) );
  mux2_1 U7588 ( .ip1(i_ssi_U_dff_tx_mem[121]), .ip2(i_apb_pwdata_int[9]), .s(
        n10174), .op(n4462) );
  mux2_1 U7589 ( .ip1(i_ssi_U_dff_tx_mem[120]), .ip2(i_apb_pwdata_int[8]), .s(
        n10174), .op(n4463) );
  mux2_1 U7590 ( .ip1(i_ssi_U_dff_tx_mem[119]), .ip2(i_apb_pwdata_int[7]), .s(
        n10174), .op(n4464) );
  mux2_1 U7591 ( .ip1(i_ssi_U_dff_tx_mem[118]), .ip2(i_apb_pwdata_int[6]), .s(
        n10174), .op(n4465) );
  mux2_1 U7592 ( .ip1(i_ssi_U_dff_tx_mem[117]), .ip2(i_apb_pwdata_int[5]), .s(
        n10174), .op(n4466) );
  mux2_1 U7593 ( .ip1(i_ssi_U_dff_tx_mem[116]), .ip2(i_apb_pwdata_int[4]), .s(
        n10174), .op(n4467) );
  mux2_1 U7594 ( .ip1(i_ssi_U_dff_tx_mem[115]), .ip2(i_apb_pwdata_int[3]), .s(
        n10175), .op(n4468) );
  mux2_1 U7595 ( .ip1(i_ssi_U_dff_tx_mem[114]), .ip2(i_apb_pwdata_int[2]), .s(
        n10175), .op(n4469) );
  mux2_1 U7596 ( .ip1(i_ssi_U_dff_tx_mem[113]), .ip2(i_apb_pwdata_int[1]), .s(
        n10175), .op(n4470) );
  mux2_1 U7597 ( .ip1(i_ssi_U_dff_tx_mem[112]), .ip2(i_apb_pwdata_int[0]), .s(
        n10175), .op(n4471) );
  mux2_1 U7598 ( .ip1(i_ssi_U_dff_tx_mem[95]), .ip2(i_apb_pwdata_int[15]), .s(
        n10176), .op(n4488) );
  mux2_1 U7599 ( .ip1(i_ssi_U_dff_tx_mem[94]), .ip2(i_apb_pwdata_int[14]), .s(
        n10176), .op(n4489) );
  mux2_1 U7600 ( .ip1(i_ssi_U_dff_tx_mem[93]), .ip2(i_apb_pwdata_int[13]), .s(
        n10176), .op(n4490) );
  mux2_1 U7601 ( .ip1(i_ssi_U_dff_tx_mem[92]), .ip2(i_apb_pwdata_int[12]), .s(
        n10176), .op(n4491) );
  mux2_1 U7602 ( .ip1(i_ssi_U_dff_tx_mem[91]), .ip2(i_apb_pwdata_int[11]), .s(
        n10173), .op(n4492) );
  mux2_1 U7603 ( .ip1(i_ssi_U_dff_tx_mem[90]), .ip2(i_apb_pwdata_int[10]), .s(
        n10173), .op(n4493) );
  mux2_1 U7604 ( .ip1(i_ssi_U_dff_tx_mem[89]), .ip2(i_apb_pwdata_int[9]), .s(
        n10173), .op(n4494) );
  mux2_1 U7605 ( .ip1(i_ssi_U_dff_tx_mem[88]), .ip2(i_apb_pwdata_int[8]), .s(
        n10173), .op(n4495) );
  mux2_1 U7606 ( .ip1(i_ssi_U_dff_tx_mem[87]), .ip2(i_apb_pwdata_int[7]), .s(
        n10173), .op(n4496) );
  mux2_1 U7607 ( .ip1(i_ssi_U_dff_tx_mem[86]), .ip2(i_apb_pwdata_int[6]), .s(
        n10173), .op(n4497) );
  mux2_1 U7608 ( .ip1(i_ssi_U_dff_tx_mem[85]), .ip2(i_apb_pwdata_int[5]), .s(
        n10173), .op(n4498) );
  mux2_1 U7609 ( .ip1(i_ssi_U_dff_tx_mem[84]), .ip2(i_apb_pwdata_int[4]), .s(
        n10173), .op(n4499) );
  mux2_1 U7610 ( .ip1(i_ssi_U_dff_tx_mem[83]), .ip2(i_apb_pwdata_int[3]), .s(
        n10176), .op(n4500) );
  mux2_1 U7611 ( .ip1(i_ssi_U_dff_tx_mem[82]), .ip2(i_apb_pwdata_int[2]), .s(
        n10176), .op(n4501) );
  mux2_1 U7612 ( .ip1(i_ssi_U_dff_tx_mem[81]), .ip2(i_apb_pwdata_int[1]), .s(
        n10176), .op(n4502) );
  mux2_1 U7613 ( .ip1(i_ssi_U_dff_tx_mem[80]), .ip2(i_apb_pwdata_int[0]), .s(
        n10176), .op(n4503) );
  mux2_1 U7614 ( .ip1(i_ssi_U_dff_tx_mem[63]), .ip2(i_apb_pwdata_int[15]), .s(
        n10177), .op(n4520) );
  mux2_1 U7615 ( .ip1(i_ssi_U_dff_tx_mem[62]), .ip2(i_apb_pwdata_int[14]), .s(
        n10177), .op(n4521) );
  mux2_1 U7616 ( .ip1(i_ssi_U_dff_tx_mem[61]), .ip2(i_apb_pwdata_int[13]), .s(
        n10177), .op(n4522) );
  mux2_1 U7617 ( .ip1(i_ssi_U_dff_tx_mem[60]), .ip2(i_apb_pwdata_int[12]), .s(
        n10177), .op(n4523) );
  mux2_1 U7618 ( .ip1(i_ssi_U_dff_tx_mem[59]), .ip2(i_apb_pwdata_int[11]), .s(
        n10172), .op(n4524) );
  mux2_1 U7619 ( .ip1(i_ssi_U_dff_tx_mem[58]), .ip2(i_apb_pwdata_int[10]), .s(
        n10172), .op(n4525) );
  mux2_1 U7620 ( .ip1(i_ssi_U_dff_tx_mem[57]), .ip2(i_apb_pwdata_int[9]), .s(
        n10172), .op(n4526) );
  mux2_1 U7621 ( .ip1(i_ssi_U_dff_tx_mem[56]), .ip2(i_apb_pwdata_int[8]), .s(
        n10172), .op(n4527) );
  mux2_1 U7622 ( .ip1(i_ssi_U_dff_tx_mem[55]), .ip2(i_apb_pwdata_int[7]), .s(
        n10172), .op(n4528) );
  mux2_1 U7623 ( .ip1(i_ssi_U_dff_tx_mem[54]), .ip2(i_apb_pwdata_int[6]), .s(
        n10172), .op(n4529) );
  mux2_1 U7624 ( .ip1(i_ssi_U_dff_tx_mem[53]), .ip2(i_apb_pwdata_int[5]), .s(
        n10172), .op(n4530) );
  mux2_1 U7625 ( .ip1(i_ssi_U_dff_tx_mem[52]), .ip2(i_apb_pwdata_int[4]), .s(
        n10172), .op(n4531) );
  mux2_1 U7626 ( .ip1(i_ssi_U_dff_tx_mem[51]), .ip2(i_apb_pwdata_int[3]), .s(
        n10177), .op(n4532) );
  mux2_1 U7627 ( .ip1(i_ssi_U_dff_tx_mem[50]), .ip2(i_apb_pwdata_int[2]), .s(
        n10177), .op(n4533) );
  mux2_1 U7628 ( .ip1(i_ssi_U_dff_tx_mem[49]), .ip2(i_apb_pwdata_int[1]), .s(
        n10177), .op(n4534) );
  mux2_1 U7629 ( .ip1(i_ssi_U_dff_tx_mem[48]), .ip2(i_apb_pwdata_int[0]), .s(
        n10177), .op(n4535) );
  mux2_1 U7630 ( .ip1(i_ssi_U_dff_tx_mem[31]), .ip2(i_apb_pwdata_int[15]), .s(
        n10178), .op(n4552) );
  mux2_1 U7631 ( .ip1(i_ssi_U_dff_tx_mem[30]), .ip2(i_apb_pwdata_int[14]), .s(
        n10178), .op(n4553) );
  mux2_1 U7632 ( .ip1(i_ssi_U_dff_tx_mem[29]), .ip2(i_apb_pwdata_int[13]), .s(
        n10178), .op(n4554) );
  mux2_1 U7633 ( .ip1(i_ssi_U_dff_tx_mem[28]), .ip2(i_apb_pwdata_int[12]), .s(
        n10178), .op(n4555) );
  mux2_1 U7634 ( .ip1(i_ssi_U_dff_tx_mem[27]), .ip2(i_apb_pwdata_int[11]), .s(
        n10171), .op(n4556) );
  mux2_1 U7635 ( .ip1(i_ssi_U_dff_tx_mem[26]), .ip2(i_apb_pwdata_int[10]), .s(
        n10171), .op(n4557) );
  mux2_1 U7636 ( .ip1(i_ssi_U_dff_tx_mem[25]), .ip2(i_apb_pwdata_int[9]), .s(
        n10171), .op(n4558) );
  mux2_1 U7637 ( .ip1(i_ssi_U_dff_tx_mem[24]), .ip2(i_apb_pwdata_int[8]), .s(
        n10171), .op(n4559) );
  mux2_1 U7638 ( .ip1(i_ssi_U_dff_tx_mem[23]), .ip2(i_apb_pwdata_int[7]), .s(
        n10171), .op(n4560) );
  mux2_1 U7639 ( .ip1(i_ssi_U_dff_tx_mem[22]), .ip2(i_apb_pwdata_int[6]), .s(
        n10171), .op(n4561) );
  mux2_1 U7640 ( .ip1(i_ssi_U_dff_tx_mem[21]), .ip2(i_apb_pwdata_int[5]), .s(
        n10171), .op(n4562) );
  mux2_1 U7641 ( .ip1(i_ssi_U_dff_tx_mem[20]), .ip2(i_apb_pwdata_int[4]), .s(
        n10171), .op(n4563) );
  mux2_1 U7642 ( .ip1(i_ssi_U_dff_tx_mem[19]), .ip2(i_apb_pwdata_int[3]), .s(
        n10178), .op(n4564) );
  mux2_1 U7643 ( .ip1(i_ssi_U_dff_tx_mem[18]), .ip2(i_apb_pwdata_int[2]), .s(
        n10178), .op(n4565) );
  mux2_1 U7644 ( .ip1(i_ssi_U_dff_tx_mem[17]), .ip2(i_apb_pwdata_int[1]), .s(
        n10178), .op(n4566) );
  mux2_1 U7645 ( .ip1(i_ssi_U_dff_tx_mem[16]), .ip2(i_apb_pwdata_int[0]), .s(
        n10178), .op(n4567) );
  mux2_1 U7646 ( .ip1(i_ssi_U_dff_tx_mem[111]), .ip2(i_apb_pwdata_int[15]), 
        .s(n10035), .op(n4472) );
  mux2_1 U7647 ( .ip1(i_ssi_U_dff_tx_mem[110]), .ip2(i_apb_pwdata_int[14]), 
        .s(n10035), .op(n4473) );
  mux2_1 U7648 ( .ip1(i_ssi_U_dff_tx_mem[109]), .ip2(i_apb_pwdata_int[13]), 
        .s(n10035), .op(n4474) );
  mux2_1 U7649 ( .ip1(i_ssi_U_dff_tx_mem[108]), .ip2(i_apb_pwdata_int[12]), 
        .s(n10035), .op(n4475) );
  mux2_1 U7650 ( .ip1(i_ssi_U_dff_tx_mem[107]), .ip2(i_apb_pwdata_int[11]), 
        .s(n10032), .op(n4476) );
  mux2_1 U7651 ( .ip1(i_ssi_U_dff_tx_mem[106]), .ip2(i_apb_pwdata_int[10]), 
        .s(n10032), .op(n4477) );
  mux2_1 U7652 ( .ip1(i_ssi_U_dff_tx_mem[105]), .ip2(i_apb_pwdata_int[9]), .s(
        n10032), .op(n4478) );
  mux2_1 U7653 ( .ip1(i_ssi_U_dff_tx_mem[104]), .ip2(i_apb_pwdata_int[8]), .s(
        n10032), .op(n4479) );
  mux2_1 U7654 ( .ip1(i_ssi_U_dff_tx_mem[103]), .ip2(i_apb_pwdata_int[7]), .s(
        n10032), .op(n4480) );
  mux2_1 U7655 ( .ip1(i_ssi_U_dff_tx_mem[102]), .ip2(i_apb_pwdata_int[6]), .s(
        n10032), .op(n4481) );
  mux2_1 U7656 ( .ip1(i_ssi_U_dff_tx_mem[101]), .ip2(i_apb_pwdata_int[5]), .s(
        n10032), .op(n4482) );
  mux2_1 U7657 ( .ip1(i_ssi_U_dff_tx_mem[100]), .ip2(i_apb_pwdata_int[4]), .s(
        n10032), .op(n4483) );
  mux2_1 U7658 ( .ip1(i_ssi_U_dff_tx_mem[99]), .ip2(i_apb_pwdata_int[3]), .s(
        n10035), .op(n4484) );
  mux2_1 U7659 ( .ip1(i_ssi_U_dff_tx_mem[98]), .ip2(i_apb_pwdata_int[2]), .s(
        n10035), .op(n4485) );
  mux2_1 U7660 ( .ip1(i_ssi_U_dff_tx_mem[97]), .ip2(i_apb_pwdata_int[1]), .s(
        n10035), .op(n4486) );
  mux2_1 U7661 ( .ip1(i_ssi_U_dff_tx_mem[96]), .ip2(i_apb_pwdata_int[0]), .s(
        n10035), .op(n4487) );
  mux2_1 U7662 ( .ip1(i_ssi_U_dff_tx_mem[79]), .ip2(i_apb_pwdata_int[15]), .s(
        n9696), .op(n4504) );
  mux2_1 U7663 ( .ip1(i_ssi_U_dff_tx_mem[78]), .ip2(i_apb_pwdata_int[14]), .s(
        n9696), .op(n4505) );
  mux2_1 U7664 ( .ip1(i_ssi_U_dff_tx_mem[77]), .ip2(i_apb_pwdata_int[13]), .s(
        n9696), .op(n4506) );
  mux2_1 U7665 ( .ip1(i_ssi_U_dff_tx_mem[76]), .ip2(i_apb_pwdata_int[12]), .s(
        n9696), .op(n4507) );
  mux2_1 U7666 ( .ip1(i_ssi_U_dff_tx_mem[75]), .ip2(i_apb_pwdata_int[11]), .s(
        n9696), .op(n4508) );
  mux2_1 U7667 ( .ip1(i_ssi_U_dff_tx_mem[74]), .ip2(i_apb_pwdata_int[10]), .s(
        n9696), .op(n4509) );
  mux2_1 U7668 ( .ip1(i_ssi_U_dff_tx_mem[73]), .ip2(i_apb_pwdata_int[9]), .s(
        n9696), .op(n4510) );
  mux2_1 U7669 ( .ip1(i_ssi_U_dff_tx_mem[72]), .ip2(i_apb_pwdata_int[8]), .s(
        n9696), .op(n4511) );
  mux2_1 U7670 ( .ip1(i_ssi_U_dff_tx_mem[71]), .ip2(i_apb_pwdata_int[7]), .s(
        n9696), .op(n4512) );
  mux2_1 U7671 ( .ip1(i_ssi_U_dff_tx_mem[70]), .ip2(i_apb_pwdata_int[6]), .s(
        n9696), .op(n4513) );
  mux2_1 U7672 ( .ip1(i_ssi_U_dff_tx_mem[69]), .ip2(i_apb_pwdata_int[5]), .s(
        n9696), .op(n4514) );
  mux2_1 U7673 ( .ip1(i_ssi_U_dff_tx_mem[68]), .ip2(i_apb_pwdata_int[4]), .s(
        n9696), .op(n4515) );
  mux2_1 U7674 ( .ip1(i_ssi_U_dff_tx_mem[67]), .ip2(i_apb_pwdata_int[3]), .s(
        n9696), .op(n4516) );
  mux2_1 U7675 ( .ip1(i_ssi_U_dff_tx_mem[66]), .ip2(i_apb_pwdata_int[2]), .s(
        n9696), .op(n4517) );
  mux2_1 U7676 ( .ip1(i_ssi_U_dff_tx_mem[65]), .ip2(i_apb_pwdata_int[1]), .s(
        n9696), .op(n4518) );
  mux2_1 U7677 ( .ip1(i_ssi_U_dff_tx_mem[64]), .ip2(i_apb_pwdata_int[0]), .s(
        n9696), .op(n4519) );
  mux2_1 U7678 ( .ip1(i_ssi_U_dff_tx_mem[47]), .ip2(i_apb_pwdata_int[15]), .s(
        n10038), .op(n4536) );
  mux2_1 U7679 ( .ip1(i_ssi_U_dff_tx_mem[46]), .ip2(i_apb_pwdata_int[14]), .s(
        n10038), .op(n4537) );
  mux2_1 U7680 ( .ip1(i_ssi_U_dff_tx_mem[45]), .ip2(i_apb_pwdata_int[13]), .s(
        n10038), .op(n4538) );
  mux2_1 U7681 ( .ip1(i_ssi_U_dff_tx_mem[44]), .ip2(i_apb_pwdata_int[12]), .s(
        n10038), .op(n4539) );
  mux2_1 U7682 ( .ip1(i_ssi_U_dff_tx_mem[43]), .ip2(i_apb_pwdata_int[11]), .s(
        n10037), .op(n4540) );
  mux2_1 U7683 ( .ip1(i_ssi_U_dff_tx_mem[42]), .ip2(i_apb_pwdata_int[10]), .s(
        n10037), .op(n4541) );
  mux2_1 U7684 ( .ip1(i_ssi_U_dff_tx_mem[41]), .ip2(i_apb_pwdata_int[9]), .s(
        n10037), .op(n4542) );
  mux2_1 U7685 ( .ip1(i_ssi_U_dff_tx_mem[40]), .ip2(i_apb_pwdata_int[8]), .s(
        n10037), .op(n4543) );
  mux2_1 U7686 ( .ip1(i_ssi_U_dff_tx_mem[39]), .ip2(i_apb_pwdata_int[7]), .s(
        n10037), .op(n4544) );
  mux2_1 U7687 ( .ip1(i_ssi_U_dff_tx_mem[38]), .ip2(i_apb_pwdata_int[6]), .s(
        n10037), .op(n4545) );
  mux2_1 U7688 ( .ip1(i_ssi_U_dff_tx_mem[37]), .ip2(i_apb_pwdata_int[5]), .s(
        n10037), .op(n4546) );
  mux2_1 U7689 ( .ip1(i_ssi_U_dff_tx_mem[36]), .ip2(i_apb_pwdata_int[4]), .s(
        n10037), .op(n4547) );
  mux2_1 U7690 ( .ip1(i_ssi_U_dff_tx_mem[35]), .ip2(i_apb_pwdata_int[3]), .s(
        n10038), .op(n4548) );
  mux2_1 U7691 ( .ip1(i_ssi_U_dff_tx_mem[34]), .ip2(i_apb_pwdata_int[2]), .s(
        n10038), .op(n4549) );
  mux2_1 U7692 ( .ip1(i_ssi_U_dff_tx_mem[33]), .ip2(i_apb_pwdata_int[1]), .s(
        n10038), .op(n4550) );
  mux2_1 U7693 ( .ip1(i_ssi_U_dff_tx_mem[32]), .ip2(i_apb_pwdata_int[0]), .s(
        n10038), .op(n4551) );
  mux2_1 U7694 ( .ip1(i_ssi_U_dff_tx_mem[15]), .ip2(i_apb_pwdata_int[15]), .s(
        n10039), .op(n4568) );
  mux2_1 U7695 ( .ip1(i_ssi_U_dff_tx_mem[14]), .ip2(i_apb_pwdata_int[14]), .s(
        n10039), .op(n4569) );
  mux2_1 U7696 ( .ip1(i_ssi_U_dff_tx_mem[13]), .ip2(i_apb_pwdata_int[13]), .s(
        n10039), .op(n4570) );
  mux2_1 U7697 ( .ip1(i_ssi_U_dff_tx_mem[12]), .ip2(i_apb_pwdata_int[12]), .s(
        n10039), .op(n4571) );
  mux2_1 U7698 ( .ip1(i_ssi_U_dff_tx_mem[11]), .ip2(i_apb_pwdata_int[11]), .s(
        n10036), .op(n4572) );
  mux2_1 U7699 ( .ip1(i_ssi_U_dff_tx_mem[10]), .ip2(i_apb_pwdata_int[10]), .s(
        n10036), .op(n4573) );
  mux2_1 U7700 ( .ip1(i_ssi_U_dff_tx_mem[9]), .ip2(i_apb_pwdata_int[9]), .s(
        n10036), .op(n4574) );
  mux2_1 U7701 ( .ip1(i_ssi_U_dff_tx_mem[8]), .ip2(i_apb_pwdata_int[8]), .s(
        n10036), .op(n4575) );
  mux2_1 U7702 ( .ip1(i_ssi_U_dff_tx_mem[7]), .ip2(i_apb_pwdata_int[7]), .s(
        n10036), .op(n4576) );
  mux2_1 U7703 ( .ip1(i_ssi_U_dff_tx_mem[6]), .ip2(i_apb_pwdata_int[6]), .s(
        n10036), .op(n4577) );
  mux2_1 U7704 ( .ip1(i_ssi_U_dff_tx_mem[5]), .ip2(i_apb_pwdata_int[5]), .s(
        n10036), .op(n4578) );
  mux2_1 U7705 ( .ip1(i_ssi_U_dff_tx_mem[4]), .ip2(i_apb_pwdata_int[4]), .s(
        n10036), .op(n4579) );
  mux2_1 U7706 ( .ip1(i_ssi_U_dff_tx_mem[3]), .ip2(i_apb_pwdata_int[3]), .s(
        n10039), .op(n4580) );
  mux2_1 U7707 ( .ip1(i_ssi_U_dff_tx_mem[2]), .ip2(i_apb_pwdata_int[2]), .s(
        n10039), .op(n4581) );
  mux2_1 U7708 ( .ip1(i_ssi_U_dff_tx_mem[1]), .ip2(i_apb_pwdata_int[1]), .s(
        n10039), .op(n4582) );
  mux2_1 U7709 ( .ip1(i_ssi_U_dff_tx_mem[0]), .ip2(i_apb_pwdata_int[0]), .s(
        n10039), .op(n4583) );
  nor2_1 U7710 ( .ip1(n9966), .ip2(i_ssi_U_mstfsm_c_done_ir), .op(n9968) );
  nor2_1 U7711 ( .ip1(n9965), .ip2(n9964), .op(n9966) );
  nand2_1 U7712 ( .ip1(n9985), .ip2(n9984), .op(n9986) );
  inv_1 U7713 ( .ip(n7087), .op(n11780) );
  mux2_1 U7714 ( .ip1(i_apb_pwdata_int[11]), .ip2(i_ssi_ctrlr0[11]), .s(n9837), 
        .op(n4598) );
  mux2_1 U7715 ( .ip1(i_apb_pwdata_int[9]), .ip2(n5281), .s(n9837), .op(n4596)
         );
  mux2_1 U7716 ( .ip1(i_apb_pwdata_int[8]), .ip2(i_ssi_tmod[0]), .s(n9837), 
        .op(n4595) );
  mux2_1 U7717 ( .ip1(i_apb_pwdata_int[13]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[13]), .s(n9896), .op(n4613) );
  mux2_1 U7718 ( .ip1(i_apb_pwdata_int[9]), .ip2(i_ssi_U_regfile_ctrlr1_int[9]), .s(n9896), .op(n4617) );
  mux2_1 U7719 ( .ip1(i_apb_pwdata_int[8]), .ip2(n5393), .s(n9896), .op(n4618)
         );
  mux2_1 U7720 ( .ip1(i_apb_pwdata_int[6]), .ip2(n5392), .s(n9896), .op(n4604)
         );
  mux2_1 U7721 ( .ip1(i_apb_pwdata_int[5]), .ip2(i_ssi_U_regfile_ctrlr1_int[5]), .s(n9896), .op(n4605) );
  mux2_1 U7722 ( .ip1(i_apb_pwdata_int[4]), .ip2(i_ssi_U_regfile_ctrlr1_int[4]), .s(n9896), .op(n4606) );
  mux2_1 U7723 ( .ip1(i_apb_pwdata_int[3]), .ip2(i_ssi_U_regfile_ctrlr1_int[3]), .s(n9896), .op(n4607) );
  mux2_1 U7724 ( .ip1(i_apb_pwdata_int[2]), .ip2(i_ssi_U_regfile_ctrlr1_int[2]), .s(n9896), .op(n4608) );
  mux2_1 U7725 ( .ip1(i_apb_pwdata_int[0]), .ip2(i_ssi_U_regfile_ctrlr1_int[0]), .s(n9896), .op(n4610) );
  mux2_1 U7726 ( .ip1(i_ssi_baudr[15]), .ip2(i_apb_pwdata_int[15]), .s(n9901), 
        .op(n4619) );
  mux2_1 U7727 ( .ip1(i_ssi_baudr[13]), .ip2(i_apb_pwdata_int[13]), .s(n9901), 
        .op(n4621) );
  mux2_1 U7728 ( .ip1(n6224), .ip2(i_apb_pwdata_int[11]), .s(n9901), .op(n4623) );
  mux2_1 U7729 ( .ip1(n11652), .ip2(i_apb_pwdata_int[9]), .s(n9901), .op(n4625) );
  mux2_1 U7730 ( .ip1(i_ssi_baudr[8]), .ip2(i_apb_pwdata_int[8]), .s(n9901), 
        .op(n4626) );
  mux2_1 U7731 ( .ip1(n5256), .ip2(i_apb_pwdata_int[7]), .s(n9901), .op(n4627)
         );
  mux2_1 U7732 ( .ip1(i_apb_pwdata_int[0]), .ip2(n11569), .s(n9788), .op(n4638) );
  mux2_1 U7733 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[23]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[23]), .s(n9398), .op(n4799) );
  mux2_2 U7734 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[22]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[22]), .s(n9372), .op(n4800) );
  mux2_1 U7735 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[21]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[21]), .s(n9398), .op(n4801) );
  mux2_1 U7736 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[20]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[20]), .s(n9395), .op(n4802) );
  mux2_1 U7737 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[19]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[19]), .s(n9396), .op(n4803) );
  mux2_1 U7738 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[18]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[18]), .s(n9395), .op(n4804) );
  mux2_1 U7739 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[17]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[17]), .s(n9398), .op(n4805) );
  mux2_1 U7740 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[16]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[16]), .s(n9398), .op(n4806) );
  mux2_1 U7741 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[15]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[15]), .s(n9396), .op(n4807) );
  mux2_1 U7742 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[14]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[14]), .s(n9396), .op(n4808) );
  mux2_1 U7743 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[13]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[13]), .s(n9398), .op(n4809) );
  mux2_1 U7744 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[12]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[12]), .s(n9396), .op(n4810) );
  mux2_1 U7745 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[11]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[11]), .s(n9398), .op(n4811) );
  mux2_1 U7746 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[10]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[10]), .s(n9396), .op(n4812) );
  mux2_1 U7747 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[9]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[9]), .s(n9398), .op(n4813) );
  mux2_1 U7748 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[8]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[8]), .s(n9396), .op(n4814) );
  mux2_1 U7749 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[7]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[7]), .s(n9398), .op(n4815) );
  mux2_1 U7750 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[6]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[6]), .s(n9396), .op(n4816) );
  mux2_1 U7751 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[5]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[5]), .s(n9398), .op(n4817) );
  mux2_1 U7752 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[4]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[4]), .s(n9396), .op(n4818) );
  mux2_1 U7753 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[3]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[3]), .s(n9398), .op(n4819) );
  mux2_1 U7754 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[2]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[2]), .s(n9396), .op(n4820) );
  mux2_1 U7755 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[1]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[1]), .s(n9398), .op(n4821) );
  mux2_1 U7756 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[0]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[0]), .s(n9396), .op(n4822) );
  or2_1 U7757 ( .ip1(n11367), .ip2(n11360), .op(n11363) );
  nand2_1 U7758 ( .ip1(n10011), .ip2(n6578), .op(n6575) );
  mux2_1 U7759 ( .ip1(i_apb_U_DW_apb_ahbsif_pipeline_c), .ip2(n9393), .s(n9392), .op(n4854) );
  nor4_1 U7760 ( .ip1(n9391), .ip2(n9390), .ip3(n9389), .ip4(n9388), .op(n9392) );
  mux2_1 U7761 ( .ip1(i_ahb_U_mux_hsel_prev[1]), .ip2(
        ex_i_ahb_AHB_Slave_RAM_hsel), .s(n11355), .op(n4856) );
  mux2_1 U7762 ( .ip1(i_ahb_U_mux_hsel_prev[3]), .ip2(
        ex_i_ahb_AHB_Slave_PWM_hsel), .s(n11355), .op(n4858) );
  mux2_1 U7763 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hsel), .s(n11355), .op(n4859) );
  nand2_1 U7764 ( .ip1(n6549), .ip2(n11182), .op(i_ahb_U_dfltslv_N4) );
  nor2_1 U7765 ( .ip1(n5579), .ip2(n5580), .op(n5588) );
  nand2_1 U7766 ( .ip1(n5588), .ip2(n5587), .op(n5805) );
  mux2_1 U7767 ( .ip1(n9706), .ip2(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[2]), 
        .s(n5330), .op(n4408) );
  or2_1 U7768 ( .ip1(n10355), .ip2(n9705), .op(n5330) );
  nand2_1 U7769 ( .ip1(n5261), .ip2(n6077), .op(n5331) );
  nand2_1 U7770 ( .ip1(n5261), .ip2(n6077), .op(n6060) );
  and2_1 U7771 ( .ip1(n5617), .ip2(n9684), .op(n5408) );
  inv_1 U7772 ( .ip(n10349), .op(n5332) );
  nand2_1 U7773 ( .ip1(n5741), .ip2(n5340), .op(n5333) );
  or2_1 U7774 ( .ip1(n6118), .ip2(n10280), .op(n5869) );
  nand2_1 U7775 ( .ip1(n6208), .ip2(n5426), .op(n6126) );
  nand2_1 U7776 ( .ip1(n5260), .ip2(n5306), .op(n5334) );
  nand2_1 U7777 ( .ip1(n5260), .ip2(n5306), .op(n5335) );
  nand2_1 U7778 ( .ip1(n5377), .ip2(n5306), .op(n6118) );
  or2_1 U7779 ( .ip1(n5454), .ip2(n5761), .op(n6117) );
  nand2_1 U7780 ( .ip1(n5628), .ip2(n5567), .op(n5569) );
  and2_1 U7781 ( .ip1(n5628), .ip2(n6287), .op(n5631) );
  inv_1 U7782 ( .ip(n9704), .op(n5366) );
  nand2_1 U7783 ( .ip1(n5354), .ip2(n5440), .op(n9704) );
  nor3_1 U7784 ( .ip1(n10346), .ip2(i_ssi_load_start_bit), .ip3(n5739), .op(
        n6130) );
  nand2_1 U7785 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[13]), .ip2(
        n5264), .op(n5336) );
  nand2_1 U7786 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[13]), .ip2(
        n5264), .op(n5793) );
  nand2_1 U7787 ( .ip1(n5309), .ip2(n5757), .op(n5758) );
  nand2_1 U7788 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[9]), .ip2(n6131), .op(n5792) );
  nand2_1 U7789 ( .ip1(n5850), .ip2(n5851), .op(n5338) );
  nand2_1 U7790 ( .ip1(n5851), .ip2(n5850), .op(n5809) );
  nand2_1 U7791 ( .ip1(n5740), .ip2(n5356), .op(n5339) );
  nand2_1 U7792 ( .ip1(n5740), .ip2(n5356), .op(n5340) );
  nand2_1 U7793 ( .ip1(n5268), .ip2(n5341), .op(n6175) );
  nand3_2 U7794 ( .ip1(n6144), .ip2(n6132), .ip3(n5373), .op(n5342) );
  nor2_1 U7795 ( .ip1(n5829), .ip2(n5375), .op(n5374) );
  or2_1 U7796 ( .ip1(n10340), .ip2(n6143), .op(n5343) );
  or2_1 U7797 ( .ip1(n5655), .ip2(n5731), .op(n5656) );
  or2_1 U7798 ( .ip1(n5810), .ip2(n5334), .op(n5344) );
  inv_1 U7799 ( .ip(n6107), .op(n5347) );
  nand2_1 U7800 ( .ip1(n6108), .ip2(n5384), .op(n6110) );
  nand2_1 U7801 ( .ip1(n5767), .ip2(n9712), .op(n6155) );
  nor2_1 U7802 ( .ip1(n5347), .ip2(n9712), .op(n5346) );
  inv_1 U7803 ( .ip(n9712), .op(n6106) );
  xnor2_1 U7804 ( .ip1(n5348), .ip2(n5522), .op(n5525) );
  nand2_1 U7805 ( .ip1(n5556), .ip2(n5281), .op(n5507) );
  nand2_1 U7806 ( .ip1(n5742), .ip2(n5350), .op(n5349) );
  nand2_1 U7807 ( .ip1(n5732), .ip2(n5733), .op(n5743) );
  nor2_1 U7808 ( .ip1(n6042), .ip2(n6041), .op(n6043) );
  nor2_1 U7809 ( .ip1(n5967), .ip2(n6168), .op(n5968) );
  nor2_1 U7810 ( .ip1(n10254), .ip2(n6168), .op(n6016) );
  nor2_1 U7811 ( .ip1(n9707), .ip2(n6168), .op(n5902) );
  nor2_1 U7812 ( .ip1(n10251), .ip2(n6168), .op(n5952) );
  nor2_1 U7813 ( .ip1(n5902), .ip2(n5903), .op(n5918) );
  nor2_1 U7814 ( .ip1(n5916), .ip2(n5915), .op(n5917) );
  nor2_1 U7815 ( .ip1(n6017), .ip2(n6016), .op(n6044) );
  nand2_1 U7816 ( .ip1(n5299), .ip2(n9058), .op(n5351) );
  nor2_1 U7817 ( .ip1(n5602), .ip2(n5601), .op(n5352) );
  nor2_1 U7818 ( .ip1(n5602), .ip2(n5601), .op(n5353) );
  inv_1 U7819 ( .ip(n5570), .op(n5573) );
  or2_1 U7820 ( .ip1(n6139), .ip2(n9683), .op(n6141) );
  nor2_1 U7821 ( .ip1(n5598), .ip2(n5690), .op(n7628) );
  inv_1 U7822 ( .ip(n5690), .op(n7626) );
  nor2_1 U7823 ( .ip1(n5969), .ip2(n5968), .op(n5993) );
  nand2_1 U7824 ( .ip1(n5644), .ip2(n5643), .op(n5666) );
  and2_1 U7825 ( .ip1(n5299), .ip2(n9058), .op(n5355) );
  nor2_1 U7826 ( .ip1(n5953), .ip2(n5952), .op(n5954) );
  inv_1 U7827 ( .ip(n11547), .op(n5356) );
  nand2_1 U7828 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[8]), .ip2(n5380), .op(n5357) );
  nand2_1 U7829 ( .ip1(n5380), .ip2(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[8]), .op(n5871) );
  or2_1 U7830 ( .ip1(n5844), .ip2(n5333), .op(n5845) );
  nand2_1 U7831 ( .ip1(n5387), .ip2(n5365), .op(n6207) );
  nand3_1 U7832 ( .ip1(n5365), .ip2(n5387), .ip3(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[3]), .op(n6209) );
  nand2_1 U7833 ( .ip1(n5856), .ip2(n5855), .op(n5857) );
  nand2_1 U7834 ( .ip1(n5366), .ip2(n5367), .op(n5835) );
  inv_1 U7835 ( .ip(n5744), .op(n5358) );
  nand2_1 U7836 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_buffer[6]), .ip2(n6061), 
        .op(n6063) );
  nand2_1 U7837 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_buffer[14]), .ip2(n6061), 
        .op(n6054) );
  nor2_1 U7838 ( .ip1(n5857), .ip2(n5858), .op(n5860) );
  nand3_1 U7839 ( .ip1(n5834), .ip2(n5374), .ip3(n5835), .op(n5858) );
  inv_1 U7840 ( .ip(n5343), .op(n5359) );
  nand2_1 U7841 ( .ip1(n6155), .ip2(n6154), .op(n6161) );
  nand2_1 U7842 ( .ip1(n5345), .ip2(n6153), .op(n6163) );
  nand2_1 U7843 ( .ip1(n5260), .ip2(n5842), .op(n5360) );
  nand2_1 U7844 ( .ip1(n5842), .ip2(n5260), .op(n5839) );
  nand2_1 U7845 ( .ip1(n5792), .ip2(n5336), .op(n5361) );
  nand2_1 U7846 ( .ip1(n5792), .ip2(n5793), .op(n5801) );
  nand2_1 U7847 ( .ip1(n5798), .ip2(n5799), .op(n5800) );
  and2_1 U7848 ( .ip1(n6105), .ip2(n10349), .op(n5364) );
  nand2_1 U7849 ( .ip1(n6144), .ip2(n10349), .op(n5365) );
  nand3_1 U7850 ( .ip1(n5688), .ip2(n5687), .ip3(n5686), .op(n11761) );
  or2_1 U7851 ( .ip1(n5361), .ip2(n5800), .op(n5367) );
  nand2_1 U7852 ( .ip1(n5682), .ip2(n5681), .op(n5688) );
  nor2_1 U7853 ( .ip1(n5680), .ip2(n5372), .op(n5681) );
  or3_1 U7854 ( .ip1(n10355), .ip2(n5332), .ip3(n5377), .op(n6145) );
  nor2_1 U7855 ( .ip1(n5800), .ip2(n5801), .op(n5880) );
  nand2_1 U7856 ( .ip1(n5342), .ip2(n5368), .op(n5424) );
  and2_1 U7857 ( .ip1(n6145), .ip2(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[11]), .op(n5368) );
  nand2_1 U7858 ( .ip1(n6195), .ip2(n6145), .op(n5369) );
  and2_1 U7859 ( .ip1(n5594), .ip2(n5575), .op(n5370) );
  xnor2_1 U7860 ( .ip1(n10381), .ip2(n10380), .op(n5371) );
  or2_1 U7861 ( .ip1(n5766), .ip2(n5765), .op(n5373) );
  and3_1 U7862 ( .ip1(n5638), .ip2(n5637), .ip3(n5636), .op(n5659) );
  inv_1 U7863 ( .ip(n9850), .op(n5376) );
  nand2_1 U7864 ( .ip1(n5355), .ip2(n10231), .op(n5399) );
  nand2_1 U7865 ( .ip1(n9058), .ip2(n5299), .op(n5643) );
  nand2_1 U7866 ( .ip1(n5264), .ip2(n10349), .op(n10352) );
  nand2_1 U7867 ( .ip1(n5264), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[15]), .op(n5832) );
  nand2_1 U7868 ( .ip1(n5264), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[12]), .op(n5870) );
  inv_1 U7869 ( .ip(n5667), .op(n5646) );
  nor2_1 U7870 ( .ip1(n5352), .ip2(n5608), .op(n5378) );
  nand4_1 U7871 ( .ip1(n5872), .ip2(n5871), .ip3(n5849), .ip4(n5870), .op(
        n5854) );
  nand4_1 U7872 ( .ip1(n5357), .ip2(n5869), .ip3(n5870), .ip4(n5872), .op(
        n5873) );
  nand2_1 U7873 ( .ip1(n5378), .ip2(n5673), .op(n5379) );
  nand2_1 U7874 ( .ip1(n10388), .ip2(n5381), .op(n10391) );
  nor2_1 U7875 ( .ip1(n10389), .ip2(n10390), .op(n5381) );
  nand2_1 U7876 ( .ip1(n6111), .ip2(n5836), .op(n5383) );
  nand2_1 U7877 ( .ip1(n6107), .ip2(n6106), .op(n5384) );
  nand2_1 U7878 ( .ip1(n5684), .ip2(n10240), .op(n5685) );
  and2_1 U7879 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[1]), .ip2(n5385), .op(n5386) );
  inv_1 U7880 ( .ip(i_ssi_U_sclkgen_ssi_cnt[0]), .op(n5385) );
  and2_1 U7881 ( .ip1(n5307), .ip2(n5385), .op(n11781) );
  nand2_1 U7882 ( .ip1(n5504), .ip2(n5503), .op(n5505) );
  or2_1 U7883 ( .ip1(n10355), .ip2(n6182), .op(n5387) );
  xor2_1 U7884 ( .ip1(i_ssi_U_mstfsm_frame_cnt[10]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[10]), .op(n5526) );
  inv_1 U7885 ( .ip(n5590), .op(n5388) );
  or2_1 U7886 ( .ip1(n5847), .ip2(n5846), .op(n5389) );
  xnor2_1 U7887 ( .ip1(n5390), .ip2(n5483), .op(n5487) );
  and2_1 U7888 ( .ip1(i_ssi_U_regfile_ctrlr1_int[1]), .ip2(n10498), .op(n5390)
         );
  nand2_1 U7889 ( .ip1(n10409), .ip2(n11569), .op(n5391) );
  nand2_1 U7890 ( .ip1(n10409), .ip2(n11569), .op(n10435) );
  xnor2_1 U7891 ( .ip1(n5502), .ip2(n5501), .op(n5503) );
  nand2_1 U7892 ( .ip1(n5690), .ip2(n5581), .op(n5586) );
  nand2_1 U7893 ( .ip1(n5351), .ip2(n5582), .op(n5585) );
  xnor2_1 U7894 ( .ip1(n5527), .ip2(n5526), .op(n5531) );
  xnor2_1 U7895 ( .ip1(n5396), .ip2(n5509), .op(n5513) );
  xnor2_1 U7896 ( .ip1(n5500), .ip2(n5499), .op(n5504) );
  or2_1 U7897 ( .ip1(n5360), .ip2(n5397), .op(n5798) );
  xor2_1 U7898 ( .ip1(i_ssi_U_mstfsm_frame_cnt[15]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[15]), .op(n5488) );
  nand2_1 U7899 ( .ip1(n10544), .ip2(i_ssi_U_regfile_ctrlr1_int[15]), .op(
        n5495) );
  inv_1 U7900 ( .ip(n11543), .op(n5398) );
  inv_1 U7901 ( .ip(n5683), .op(n5684) );
  nand3_1 U7902 ( .ip1(n10288), .ip2(n5650), .ip3(n5649), .op(n5651) );
  nor2_1 U7903 ( .ip1(n7629), .ip2(n5651), .op(n5652) );
  nor2_1 U7904 ( .ip1(n5400), .ip2(n8382), .op(n8383) );
  inv_1 U7905 ( .ip(n5599), .op(n5542) );
  inv_2 U7906 ( .ip(i_ssi_dfs[0]), .op(n10198) );
  inv_1 U7907 ( .ip(n6297), .op(n10483) );
  xor2_2 U7908 ( .ip1(i_ssi_U_mstfsm_bit_cnt[0]), .ip2(n10198), .op(n6297) );
  nand4_1 U7909 ( .ip1(i_ssi_U_mstfsm_frame_cnt[16]), .ip2(n10541), .ip3(n9082), .ip4(n10536), .op(n9086) );
  nand3_1 U7910 ( .ip1(n9082), .ip2(n6305), .ip3(n10536), .op(n6306) );
  or2_1 U7911 ( .ip1(n10536), .ip2(i_ssi_U_mstfsm_frame_cnt[16]), .op(n9085)
         );
  nand2_1 U7912 ( .ip1(i_ssi_U_mstfsm_frame_cnt[12]), .ip2(n10536), .op(n10538) );
  nand2_1 U7913 ( .ip1(n6162), .ip2(n6163), .op(n4401) );
  nand2_1 U7914 ( .ip1(n6160), .ip2(n6161), .op(n6162) );
  nand2_1 U7915 ( .ip1(n6110), .ip2(n6109), .op(n4403) );
  nand2_1 U7916 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[7]), .ip2(n5346), .op(n6109) );
  or2_1 U7917 ( .ip1(n5260), .ip2(n5843), .op(n5844) );
  nor2_1 U7918 ( .ip1(n5533), .ip2(n5532), .op(n5558) );
  nand3_1 U7919 ( .ip1(n6077), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[9]), 
        .ip3(n5261), .op(n6084) );
  inv_1 U7920 ( .ip(n5666), .op(n5645) );
  inv_1 U7921 ( .ip(n5252), .op(n9985) );
  nor2_1 U7922 ( .ip1(n10258), .ip2(n5331), .op(n5940) );
  nor2_1 U7923 ( .ip1(n10256), .ip2(n5331), .op(n6042) );
  nor2_1 U7924 ( .ip1(n10276), .ip2(n6060), .op(n5969) );
  nor2_1 U7925 ( .ip1(n10257), .ip2(n6060), .op(n5915) );
  inv_1 U7926 ( .ip(n6078), .op(n6079) );
  nand2_1 U7927 ( .ip1(i_ssi_mwcr[1]), .ip2(n5477), .op(n5615) );
  inv_1 U7928 ( .ip(i_ssi_mwcr[0]), .op(n6978) );
  inv_1 U7929 ( .ip(n6076), .op(n5403) );
  and2_1 U7930 ( .ip1(n10533), .ip2(i_ssi_U_regfile_ctrlr1_int[11]), .op(n5405) );
  xor2_1 U7931 ( .ip1(i_ssi_rx_push), .ip2(n5266), .op(n4451) );
  nand2_1 U7932 ( .ip1(n6177), .ip2(n6176), .op(n6184) );
  nor2_4 U7933 ( .ip1(n6230), .ip2(n5414), .op(n6236) );
  inv_2 U7934 ( .ip(n10104), .op(n11369) );
  and2_1 U7935 ( .ip1(i_i2c_fifo_rst_n), .ip2(n6693), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N36) );
  and3_1 U7936 ( .ip1(n6618), .ip2(n6461), .ip3(n6462), .op(n5412) );
  xor2_1 U7937 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[10]), .ip2(n6235), .op(n5414) );
  and2_1 U7938 ( .ip1(n6222), .ip2(n6236), .op(n5415) );
  inv_2 U7939 ( .ip(n5442), .op(n11497) );
  or3_1 U7940 ( .ip1(n6442), .ip2(n6441), .ip3(n6440), .op(n5416) );
  or3_1 U7941 ( .ip1(n6385), .ip2(n6384), .ip3(n6383), .op(n5417) );
  ab_or_c_or_d U7942 ( .ip1(n6410), .ip2(n6409), .ip3(n6408), .ip4(n6407), 
        .op(n5418) );
  and2_1 U7943 ( .ip1(n10719), .ip2(n7716), .op(n5419) );
  xor2_1 U7944 ( .ip1(n8181), .ip2(n8005), .op(n5420) );
  inv_1 U7945 ( .ip(n6470), .op(n9449) );
  or2_1 U7946 ( .ip1(n10108), .ip2(n9381), .op(n5421) );
  and2_1 U7947 ( .ip1(n9949), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[3]), .op(n5422) );
  and2_1 U7948 ( .ip1(i_ssi_rxd), .ip2(n5593), .op(n5423) );
  and2_1 U7949 ( .ip1(n10541), .ip2(n10540), .op(n5425) );
  and2_1 U7950 ( .ip1(n6123), .ip2(n6122), .op(n5426) );
  or2_1 U7951 ( .ip1(n10350), .ip2(n6188), .op(n5427) );
  and2_1 U7952 ( .ip1(n6184), .ip2(n6181), .op(n5428) );
  inv_1 U7953 ( .ip(n6169), .op(n6172) );
  and2_1 U7954 ( .ip1(n6341), .ip2(n6465), .op(n5431) );
  or2_1 U7955 ( .ip1(n5803), .ip2(n5379), .op(n5432) );
  or2_1 U7956 ( .ip1(n5803), .ip2(n5379), .op(n5435) );
  nand2_1 U7957 ( .ip1(n5263), .ip2(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[3]), .op(n5436) );
  inv_1 U7958 ( .ip(n5281), .op(n5482) );
  or2_1 U7959 ( .ip1(n6315), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_hcnt_cmplt_int), .op(n5437) );
  inv_1 U7960 ( .ip(n6060), .op(n6051) );
  and2_1 U7961 ( .ip1(n5261), .ip2(n9714), .op(n5440) );
  inv_1 U7962 ( .ip(n5566), .op(n6287) );
  or2_1 U7963 ( .ip1(n11369), .ip2(n10109), .op(n5442) );
  and2_1 U7964 ( .ip1(n6289), .ip2(n10490), .op(n5443) );
  and2_1 U7965 ( .ip1(n5377), .ip2(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[15]), .op(n5444) );
  and2_1 U7966 ( .ip1(n8108), .ip2(n8107), .op(n5445) );
  nor2_1 U7967 ( .ip1(n10430), .ip2(n11093), .op(n5446) );
  and2_1 U7968 ( .ip1(n8163), .ip2(n8013), .op(n5447) );
  and2_1 U7969 ( .ip1(n6136), .ip2(n11569), .op(n5448) );
  nand3_1 U7970 ( .ip1(n6221), .ip2(n6220), .ip3(n6219), .op(n6222) );
  and2_1 U7971 ( .ip1(n6217), .ip2(n6218), .op(n5451) );
  or2_1 U7972 ( .ip1(n8151), .ip2(n8027), .op(n5452) );
  and2_1 U7973 ( .ip1(n11760), .ip2(n9672), .op(n5453) );
  or3_1 U7974 ( .ip1(i_ssi_cfs[2]), .ip2(i_ssi_cfs[3]), .ip3(n5760), .op(n5454) );
  and2_1 U7975 ( .ip1(n5593), .ip2(n5627), .op(n5455) );
  and2_1 U7976 ( .ip1(n8905), .ip2(n8904), .op(n5456) );
  nor2_1 U7977 ( .ip1(n5966), .ip2(n5965), .op(n10276) );
  inv_1 U7978 ( .ip(n10276), .op(n10277) );
  nor2_1 U7979 ( .ip1(n6039), .ip2(n6038), .op(n10250) );
  inv_1 U7980 ( .ip(n10250), .op(n6189) );
  nor2_1 U7981 ( .ip1(n6027), .ip2(n6026), .op(n10256) );
  inv_1 U7982 ( .ip(n10256), .op(n6164) );
  nor2_1 U7983 ( .ip1(n5914), .ip2(n5913), .op(n10257) );
  inv_1 U7984 ( .ip(n10257), .op(n6156) );
  nor2_1 U7985 ( .ip1(n5713), .ip2(n5712), .op(n5904) );
  inv_1 U7986 ( .ip(n5904), .op(n5714) );
  or2_1 U7987 ( .ip1(n5826), .ip2(n5825), .op(n5458) );
  nor2_1 U7988 ( .ip1(n6005), .ip2(n6004), .op(n10342) );
  inv_1 U7989 ( .ip(n10342), .op(n10343) );
  nor2_1 U7990 ( .ip1(n5901), .ip2(n5900), .op(n10253) );
  inv_1 U7991 ( .ip(n10253), .op(n6146) );
  and2_1 U7992 ( .ip1(n9017), .ip2(n9016), .op(n5459) );
  inv_2 U7993 ( .ip(n9714), .op(n10340) );
  and2_1 U7994 ( .ip1(n6072), .ip2(n10278), .op(n5460) );
  xor2_1 U7995 ( .ip1(n8083), .ip2(n8097), .op(n5461) );
  or2_1 U7996 ( .ip1(n6443), .ip2(n6361), .op(n5463) );
  and2_1 U7997 ( .ip1(n8977), .ip2(n10977), .op(n5464) );
  inv_1 U7998 ( .ip(n8966), .op(n6727) );
  xor2_1 U7999 ( .ip1(n8132), .ip2(n8131), .op(n8921) );
  xor2_1 U8000 ( .ip1(n8168), .ip2(n8167), .op(n5465) );
  inv_1 U8001 ( .ip(n8967), .op(n6734) );
  and2_1 U8002 ( .ip1(n6394), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[5]), .op(n5466) );
  nand2_1 U8003 ( .ip1(n8039), .ip2(n8038), .op(n8093) );
  xor2_1 U8004 ( .ip1(n7979), .ip2(n6764), .op(n9022) );
  xor2_1 U8005 ( .ip1(n8155), .ip2(n8154), .op(n5467) );
  and2_1 U8006 ( .ip1(n6422), .ip2(n6423), .op(n5468) );
  and2_1 U8007 ( .ip1(n6424), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[7]), .op(n5469) );
  inv_1 U8008 ( .ip(n8079), .op(n8094) );
  nand2_1 U8009 ( .ip1(n10981), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[8]), .op(n10984) );
  inv_1 U8010 ( .ip(n10984), .op(n10986) );
  inv_1 U8011 ( .ip(n8988), .op(n6802) );
  nor2_1 U8012 ( .ip1(n8940), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[0]), .op(n5470) );
  and2_1 U8013 ( .ip1(n7114), .ip2(n7252), .op(n5471) );
  inv_1 U8014 ( .ip(n10843), .op(n10749) );
  and2_1 U8015 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[2]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[1]), .op(n5472) );
  and2_1 U8016 ( .ip1(n5422), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[4]), .op(n5473) );
  or2_1 U8017 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_hwrite_c), .ip2(n9381), .op(
        n5474) );
  inv_1 U8018 ( .ip(i_ahb_U_dfltslv_current_state), .op(n6549) );
  nor2_1 U8019 ( .ip1(n5538), .ip2(n9059), .op(n9684) );
  inv_1 U8020 ( .ip(n5641), .op(n5642) );
  inv_1 U8021 ( .ip(n5575), .op(n6137) );
  nor2_1 U8022 ( .ip1(n5536), .ip2(n9056), .op(n5575) );
  nand2_1 U8023 ( .ip1(n10473), .ip2(n6281), .op(n6298) );
  inv_1 U8024 ( .ip(n6298), .op(n10486) );
  nand2_1 U8025 ( .ip1(n6138), .ip2(i_ssi_sclk_re), .op(n5475) );
  nand2_1 U8026 ( .ip1(i_ssi_U_mstfsm_c_done_ir), .ip2(i_ssi_sclk_re), .op(
        n5476) );
  nand2_1 U8027 ( .ip1(i_ssi_U_mstfsm_c_done_ir), .ip2(i_ssi_sclk_fe), .op(
        n5477) );
  and2_1 U8028 ( .ip1(n6980), .ip2(n5749), .op(n5478) );
  inv_1 U8029 ( .ip(i_ssi_U_mstfsm_last_frame), .op(n5574) );
  nand2_1 U8030 ( .ip1(n5547), .ip2(n5546), .op(n10287) );
  nand2_1 U8031 ( .ip1(n6286), .ip2(n6285), .op(n10542) );
  or2_1 U8032 ( .ip1(n10541), .ip2(i_ssi_U_mstfsm_frame_cnt[16]), .op(n5479)
         );
  and2_1 U8033 ( .ip1(n5479), .ip2(n9083), .op(n5480) );
  nor2_1 U8034 ( .ip1(n10539), .ip2(n10535), .op(n9082) );
  inv_1 U8035 ( .ip(n9082), .op(n10537) );
  inv_1 U8036 ( .ip(i_ssi_U_mstfsm_frame_cnt[16]), .op(n9084) );
  inv_1 U8037 ( .ip(i_ssi_U_mstfsm_bit_cnt[2]), .op(n5565) );
  inv_1 U8038 ( .ip(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[11]), .op(n5874)
         );
  inv_1 U8039 ( .ip(i_i2c_ic_rst_n), .op(n11747) );
  inv_1 U8040 ( .ip(i_i2c_ic_rst_n), .op(n11726) );
  inv_1 U8041 ( .ip(i_ssi_ser_0_), .op(n10547) );
  inv_1 U8042 ( .ip(i_ssi_U_mstfsm_frame_cnt[1]), .op(n10498) );
  xor2_1 U8043 ( .ip1(i_ssi_U_mstfsm_frame_cnt[2]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[2]), .op(n5483) );
  inv_1 U8044 ( .ip(i_ssi_U_mstfsm_frame_cnt[5]), .op(n10513) );
  nand2_1 U8045 ( .ip1(n10513), .ip2(i_ssi_U_regfile_ctrlr1_int[5]), .op(n5485) );
  xor2_1 U8046 ( .ip1(i_ssi_U_mstfsm_frame_cnt[6]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[6]), .op(n5484) );
  nand2_1 U8047 ( .ip1(n6305), .ip2(i_ssi_U_regfile_ctrlr1_int[14]), .op(n5489) );
  inv_1 U8048 ( .ip(i_ssi_U_mstfsm_frame_cnt[11]), .op(n10533) );
  fulladder U8049 ( .a(n10498), .b(i_ssi_U_regfile_ctrlr1_int[1]), .ci(
        i_ssi_U_regfile_ctrlr1_int[0]), .s(n5498) );
  xnor2_1 U8050 ( .ip1(i_ssi_U_mstfsm_frame_cnt[16]), .ip2(n5495), .op(n5496)
         );
  nand2_1 U8051 ( .ip1(n5497), .ip2(n5498), .op(n5506) );
  inv_1 U8052 ( .ip(i_ssi_U_mstfsm_frame_cnt[6]), .op(n10519) );
  inv_1 U8053 ( .ip(i_ssi_U_mstfsm_frame_cnt[3]), .op(n10507) );
  xor2_1 U8054 ( .ip1(i_ssi_U_mstfsm_frame_cnt[4]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[4]), .op(n5501) );
  inv_1 U8055 ( .ip(i_ssi_U_mstfsm_frame_cnt[10]), .op(n10531) );
  inv_1 U8056 ( .ip(i_ssi_U_mstfsm_frame_cnt[12]), .op(n10535) );
  inv_1 U8057 ( .ip(i_ssi_U_mstfsm_frame_cnt[2]), .op(n10504) );
  nand2_1 U8058 ( .ip1(n10504), .ip2(i_ssi_U_regfile_ctrlr1_int[2]), .op(n5515) );
  xor2_1 U8059 ( .ip1(i_ssi_U_mstfsm_frame_cnt[3]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[3]), .op(n5514) );
  inv_1 U8060 ( .ip(i_ssi_U_mstfsm_frame_cnt[4]), .op(n10509) );
  nand2_1 U8061 ( .ip1(n10509), .ip2(i_ssi_U_regfile_ctrlr1_int[4]), .op(n5517) );
  xor2_1 U8062 ( .ip1(i_ssi_U_mstfsm_frame_cnt[5]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[5]), .op(n5516) );
  inv_1 U8063 ( .ip(i_ssi_U_mstfsm_frame_cnt[7]), .op(n10521) );
  xor2_1 U8064 ( .ip1(i_ssi_U_mstfsm_frame_cnt[8]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[8]), .op(n5522) );
  inv_1 U8065 ( .ip(i_ssi_U_mstfsm_frame_cnt[13]), .op(n10539) );
  inv_1 U8066 ( .ip(i_ssi_U_mstfsm_frame_cnt[9]), .op(n10527) );
  inv_1 U8067 ( .ip(i_ssi_U_mstfsm_frame_cnt[8]), .op(n10525) );
  nand2_1 U8068 ( .ip1(n10525), .ip2(i_ssi_U_regfile_ctrlr1_int[8]), .op(n5529) );
  xor2_1 U8069 ( .ip1(i_ssi_U_mstfsm_frame_cnt[9]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[9]), .op(n5528) );
  xor2_2 U8070 ( .ip1(n5529), .ip2(n5528), .op(n5530) );
  inv_1 U8071 ( .ip(i_ssi_U_mstfsm_c_state[1]), .op(n5543) );
  nand2_1 U8072 ( .ip1(n5543), .ip2(i_ssi_U_mstfsm_c_state[0]), .op(n5536) );
  nand2_1 U8073 ( .ip1(n6281), .ip2(i_ssi_U_mstfsm_c_state[2]), .op(n9056) );
  nor2_1 U8074 ( .ip1(i_ssi_U_mstfsm_c_state[2]), .ip2(n6281), .op(n6284) );
  inv_1 U8075 ( .ip(i_ssi_U_mstfsm_c_state[0]), .op(n5647) );
  nand2_1 U8076 ( .ip1(n5537), .ip2(i_ssi_U_mstfsm_c_state[1]), .op(n5541) );
  nand2_1 U8077 ( .ip1(i_ssi_U_mstfsm_c_state[0]), .ip2(
        i_ssi_U_mstfsm_c_state[1]), .op(n9686) );
  nor2_1 U8078 ( .ip1(n6281), .ip2(n9686), .op(n5611) );
  inv_2 U8079 ( .ip(i_ssi_ssi_en_int), .op(n11148) );
  and2_1 U8080 ( .ip1(n5611), .ip2(n11148), .op(n5635) );
  nand2_1 U8081 ( .ip1(n6281), .ip2(i_ssi_U_mstfsm_c_state[1]), .op(n5538) );
  inv_1 U8082 ( .ip(i_ssi_U_mstfsm_c_state[2]), .op(n6283) );
  nand2_1 U8083 ( .ip1(n6283), .ip2(i_ssi_U_mstfsm_c_state[0]), .op(n9059) );
  and2_1 U8084 ( .ip1(n9684), .ip2(i_ssi_U_mstfsm_c_done_ir), .op(n5610) );
  nor2_1 U8085 ( .ip1(n5578), .ip2(n5400), .op(n5540) );
  not_ab_or_c_or_d U8086 ( .ip1(n6284), .ip2(n5541), .ip3(n5635), .ip4(n5540), 
        .op(n5552) );
  nor2_1 U8087 ( .ip1(i_ssi_U_mstfsm_c_state[0]), .ip2(n5543), .op(n9057) );
  and2_1 U8088 ( .ip1(i_ssi_U_mstfsm_c_state[2]), .ip2(
        i_ssi_U_mstfsm_c_state[3]), .op(n5568) );
  nand2_1 U8089 ( .ip1(n9057), .ip2(n5568), .op(n5601) );
  nand2_1 U8090 ( .ip1(n5299), .ip2(n5545), .op(n5548) );
  nor2_1 U8091 ( .ip1(i_ssi_U_mstfsm_c_state[1]), .ip2(n6281), .op(n5547) );
  and2_1 U8092 ( .ip1(i_ssi_U_mstfsm_c_state[0]), .ip2(
        i_ssi_U_mstfsm_c_state[2]), .op(n5546) );
  nor2_1 U8093 ( .ip1(n9686), .ip2(n9056), .op(n10231) );
  nor3_1 U8094 ( .ip1(n5550), .ip2(n5570), .ip3(n5549), .op(n5551) );
  nand2_1 U8095 ( .ip1(n5556), .ip2(n5555), .op(n5560) );
  inv_1 U8096 ( .ip(n5755), .op(n5561) );
  inv_1 U8097 ( .ip(n5665), .op(n5562) );
  or2_1 U8098 ( .ip1(i_ssi_U_mstfsm_bit_cnt[4]), .ip2(n5663), .op(n5563) );
  nor2_1 U8099 ( .ip1(i_ssi_U_mstfsm_c_state[1]), .ip2(
        i_ssi_U_mstfsm_c_state[0]), .op(n6282) );
  nand2_1 U8100 ( .ip1(n5568), .ip2(n6282), .op(n5641) );
  nor2_1 U8101 ( .ip1(i_ssi_U_mstfsm_c_state[0]), .ip2(n9056), .op(n5576) );
  nand2_1 U8102 ( .ip1(n5599), .ip2(n5583), .op(n5584) );
  inv_1 U8103 ( .ip(n5715), .op(n5595) );
  inv_1 U8104 ( .ip(n10287), .op(n5593) );
  inv_1 U8105 ( .ip(n9057), .op(n5598) );
  buf_1 U8106 ( .ip(i_ssi_baud2), .op(n5624) );
  nand2_1 U8107 ( .ip1(n10288), .ip2(i_ssi_sclk_fe), .op(n5600) );
  nor2_1 U8108 ( .ip1(n7628), .ip2(n5353), .op(n5603) );
  nand2_1 U8109 ( .ip1(n5438), .ip2(n5603), .op(n10303) );
  inv_1 U8110 ( .ip(n10303), .op(n5604) );
  or2_1 U8111 ( .ip1(n10306), .ip2(n5604), .op(n5605) );
  nand2_1 U8112 ( .ip1(n5611), .ip2(n11148), .op(n5612) );
  inv_1 U8113 ( .ip(i_ssi_mwcr[1]), .op(n5614) );
  nand2_1 U8114 ( .ip1(n5476), .ip2(n5614), .op(n5616) );
  inv_1 U8115 ( .ip(n9684), .op(n9967) );
  nand2_1 U8116 ( .ip1(i_ssi_baud2), .ip2(i_ssi_U_mstfsm_c_done_ir), .op(n5617) );
  nor3_1 U8117 ( .ip1(n5608), .ip2(n7628), .ip3(n5803), .op(n5620) );
  nor2_1 U8118 ( .ip1(n7626), .ip2(n10232), .op(n5623) );
  nand2_1 U8119 ( .ip1(n5624), .ip2(n5595), .op(n5625) );
  nand2_1 U8120 ( .ip1(i_ssi_rxd), .ip2(n5626), .op(n5627) );
  inv_1 U8121 ( .ip(n6282), .op(n5629) );
  nor2_1 U8122 ( .ip1(n9056), .ip2(n5629), .op(n5630) );
  nand2_1 U8123 ( .ip1(n5631), .ip2(n5630), .op(n5638) );
  nand2_1 U8124 ( .ip1(n6284), .ip2(n6282), .op(n8378) );
  nor2_1 U8125 ( .ip1(n7626), .ip2(n8378), .op(n5634) );
  inv_1 U8126 ( .ip(n5632), .op(n5633) );
  xor2_2 U8127 ( .ip1(i_ssi_U_mstfsm_bit_cnt[0]), .ip2(i_ssi_dfs[0]), .op(
        n5664) );
  nor2_1 U8128 ( .ip1(n5734), .ip2(n5732), .op(n5657) );
  nor2_1 U8129 ( .ip1(i_ssi_U_mstfsm_c_state[3]), .ip2(
        i_ssi_U_mstfsm_c_state[2]), .op(n5648) );
  inv_1 U8130 ( .ip(i_ssi_mst_contention), .op(n5650) );
  nor2_1 U8131 ( .ip1(i_ssi_U_mstfsm_c_state[1]), .ip2(n5654), .op(n5655) );
  or2_1 U8132 ( .ip1(n5455), .ip2(n5660), .op(n5661) );
  inv_1 U8164 ( .ip(HRESETn_hresetn), .op(n11759) );
  inv_1 U8165 ( .ip(i_ssi_U_mstfsm_ss_in_n_sync), .op(n10240) );
  nand2_1 U8166 ( .ip1(n5642), .ip2(n5351), .op(n6139) );
  nand2_1 U8167 ( .ip1(i_ssi_U_mstfsm_c_state[1]), .ip2(i_ssi_sclk_re), .op(
        n5691) );
  nand2_1 U8168 ( .ip1(n5755), .ip2(n5692), .op(n5698) );
  inv_1 U8169 ( .ip(i_ssi_U_mstfsm_tx_load_en_int), .op(n5749) );
  nand2_1 U8170 ( .ip1(i_ssi_U_mstfsm_c_state[0]), .ip2(i_ssi_sclk_re), .op(
        n5693) );
  nor2_1 U8171 ( .ip1(n5693), .ip2(n9056), .op(n6980) );
  nand2_1 U8172 ( .ip1(i_ssi_U_mstfsm_c_state[1]), .ip2(
        i_ssi_U_mstfsm_abort_ir), .op(n5694) );
  inv_1 U8173 ( .ip(i_ssi_tx_rd_addr[1]), .op(n5699) );
  nand2_1 U8174 ( .ip1(n5699), .ip2(i_ssi_tx_rd_addr[2]), .op(n5705) );
  nand2_1 U8175 ( .ip1(n5812), .ip2(i_ssi_U_dff_tx_mem[42]), .op(n5704) );
  nor2_1 U8176 ( .ip1(i_ssi_tx_rd_addr[2]), .ip2(i_ssi_tx_rd_addr[1]), .op(
        n5700) );
  and2_1 U8177 ( .ip1(n5700), .ip2(i_ssi_tx_rd_addr[0]), .op(n6028) );
  nand2_1 U8178 ( .ip1(n6028), .ip2(i_ssi_U_dff_tx_mem[106]), .op(n5703) );
  nand2_1 U8179 ( .ip1(n5769), .ip2(i_ssi_U_dff_tx_mem[90]), .op(n5702) );
  nand2_1 U8180 ( .ip1(n6029), .ip2(i_ssi_U_dff_tx_mem[122]), .op(n5701) );
  nand4_1 U8181 ( .ip1(n5704), .ip2(n5703), .ip3(n5702), .ip4(n5701), .op(
        n5713) );
  nand2_1 U8182 ( .ip1(n5817), .ip2(i_ssi_U_dff_tx_mem[58]), .op(n5711) );
  nand2_1 U8183 ( .ip1(i_ssi_tx_rd_addr[0]), .ip2(i_ssi_tx_rd_addr[1]), .op(
        n5706) );
  nand2_1 U8184 ( .ip1(n5818), .ip2(i_ssi_U_dff_tx_mem[74]), .op(n5710) );
  nand2_1 U8185 ( .ip1(i_ssi_tx_rd_addr[1]), .ip2(i_ssi_tx_rd_addr[2]), .op(
        n9953) );
  nand2_1 U8186 ( .ip1(n5819), .ip2(i_ssi_U_dff_tx_mem[26]), .op(n5709) );
  inv_1 U8187 ( .ip(i_ssi_tx_rd_addr[2]), .op(n5707) );
  nor2_2 U8188 ( .ip1(n5707), .ip2(n5706), .op(n5820) );
  nand2_1 U8189 ( .ip1(n5820), .ip2(i_ssi_U_dff_tx_mem[10]), .op(n5708) );
  nand4_1 U8190 ( .ip1(n5711), .ip2(n5710), .ip3(n5709), .ip4(n5708), .op(
        n5712) );
  nor3_2 U8191 ( .ip1(n5715), .ip2(n5481), .ip3(n10287), .op(
        i_ssi_load_start_bit) );
  inv_2 U8192 ( .ip(i_ssi_load_start_bit), .op(n9717) );
  nand2_1 U8193 ( .ip1(n10346), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[10]), 
        .op(n5729) );
  inv_1 U8194 ( .ip(i_ssi_tmod[0]), .op(n5722) );
  nor2_1 U8195 ( .ip1(i_ssi_U_mstfsm_spi1_control), .ip2(
        i_ssi_U_mstfsm_spi0_control), .op(n5721) );
  and2_1 U8196 ( .ip1(i_ssi_U_mstfsm_c_state[2]), .ip2(i_ssi_sclk_re), .op(
        n5724) );
  and2_1 U8197 ( .ip1(n6282), .ip2(n5724), .op(n10473) );
  and2_1 U8198 ( .ip1(n9684), .ip2(i_ssi_sclk_re), .op(n11702) );
  nand2_2 U8199 ( .ip1(n5727), .ip2(n5726), .op(n9714) );
  nand2_1 U8200 ( .ip1(n9714), .ip2(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[9]), .op(n5728) );
  nand4_1 U8201 ( .ip1(n5730), .ip2(n9717), .ip3(n5729), .ip4(n5728), .op(
        n5768) );
  inv_1 U8202 ( .ip(n5736), .op(n5735) );
  nand2_1 U8203 ( .ip1(n5736), .ip2(n5398), .op(n5737) );
  nand2_2 U8204 ( .ip1(n5737), .ip2(n5738), .op(n6188) );
  nor4_1 U8205 ( .ip1(n10346), .ip2(i_ssi_load_start_bit), .ip3(n6188), .ip4(
        n5739), .op(n5748) );
  inv_1 U8206 ( .ip(i_ssi_dfs[3]), .op(n5744) );
  nand2_1 U8207 ( .ip1(n5744), .ip2(n5349), .op(n5747) );
  inv_1 U8208 ( .ip(i_ssi_cfs[3]), .op(n5745) );
  nand2_1 U8209 ( .ip1(n5748), .ip2(n5403), .op(n5767) );
  nor2_2 U8210 ( .ip1(n6111), .ip2(n10232), .op(n5887) );
  nand2_1 U8211 ( .ip1(n5751), .ip2(i_ssi_U_mstfsm_tx_load_en_int), .op(n5811)
         );
  inv_1 U8212 ( .ip(i_ssi_cfs[1]), .op(n5759) );
  inv_1 U8213 ( .ip(i_ssi_cfs[0]), .op(n5806) );
  nand2_1 U8214 ( .ip1(n5759), .ip2(n5806), .op(n5760) );
  nor2_1 U8215 ( .ip1(n5398), .ip2(i_ssi_dfs[0]), .op(n5762) );
  nor2_1 U8216 ( .ip1(i_ssi_dfs[3]), .ip2(i_ssi_dfs[2]), .op(n10205) );
  nand2_1 U8217 ( .ip1(n5762), .ip2(n10205), .op(n6659) );
  mux2_1 U8218 ( .ip1(n5768), .ip2(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[10]), .s(n5345), .op(n4400) );
  nand2_1 U8219 ( .ip1(n5812), .ip2(i_ssi_U_dff_tx_mem[39]), .op(n5773) );
  nand2_1 U8220 ( .ip1(n6028), .ip2(i_ssi_U_dff_tx_mem[103]), .op(n5772) );
  nand2_1 U8221 ( .ip1(n5769), .ip2(i_ssi_U_dff_tx_mem[87]), .op(n5771) );
  nand2_1 U8222 ( .ip1(n6029), .ip2(i_ssi_U_dff_tx_mem[119]), .op(n5770) );
  nand4_1 U8223 ( .ip1(n5773), .ip2(n5772), .ip3(n5771), .ip4(n5770), .op(
        n5779) );
  nand2_1 U8224 ( .ip1(n5817), .ip2(i_ssi_U_dff_tx_mem[55]), .op(n5777) );
  nand2_1 U8225 ( .ip1(n5818), .ip2(i_ssi_U_dff_tx_mem[71]), .op(n5776) );
  nand2_1 U8226 ( .ip1(n5819), .ip2(i_ssi_U_dff_tx_mem[23]), .op(n5775) );
  nand2_1 U8227 ( .ip1(n5820), .ip2(i_ssi_U_dff_tx_mem[7]), .op(n5774) );
  nand4_1 U8228 ( .ip1(n5777), .ip2(n5776), .ip3(n5775), .ip4(n5774), .op(
        n5778) );
  mux2_1 U8229 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_buffer[7]), .ip2(n5780), 
        .s(n5739), .op(n4420) );
  nand2_1 U8230 ( .ip1(n5812), .ip2(i_ssi_U_dff_tx_mem[40]), .op(n5784) );
  nand2_1 U8231 ( .ip1(n6028), .ip2(i_ssi_U_dff_tx_mem[104]), .op(n5783) );
  nand2_1 U8232 ( .ip1(n5769), .ip2(i_ssi_U_dff_tx_mem[88]), .op(n5782) );
  nand2_1 U8233 ( .ip1(n6029), .ip2(i_ssi_U_dff_tx_mem[120]), .op(n5781) );
  nand4_1 U8234 ( .ip1(n5784), .ip2(n5783), .ip3(n5782), .ip4(n5781), .op(
        n5790) );
  nand2_1 U8235 ( .ip1(n5817), .ip2(i_ssi_U_dff_tx_mem[56]), .op(n5788) );
  nand2_1 U8236 ( .ip1(n5818), .ip2(i_ssi_U_dff_tx_mem[72]), .op(n5787) );
  nand2_1 U8237 ( .ip1(n5819), .ip2(i_ssi_U_dff_tx_mem[24]), .op(n5786) );
  nand2_1 U8238 ( .ip1(n5820), .ip2(i_ssi_U_dff_tx_mem[8]), .op(n5785) );
  nand4_1 U8239 ( .ip1(n5788), .ip2(n5787), .ip3(n5786), .ip4(n5785), .op(
        n5789) );
  mux2_1 U8240 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_buffer[8]), .ip2(n5791), 
        .s(n5739), .op(n4419) );
  mux2_1 U8241 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_buffer[10]), .ip2(n5714), 
        .s(n5739), .op(n4417) );
  nand2_1 U8242 ( .ip1(n5328), .ip2(n5794), .op(n5795) );
  or2_1 U8243 ( .ip1(n5887), .ip2(n5886), .op(n10348) );
  nand2_1 U8244 ( .ip1(n5812), .ip2(i_ssi_U_dff_tx_mem[32]), .op(n5816) );
  nand2_1 U8245 ( .ip1(n6028), .ip2(i_ssi_U_dff_tx_mem[96]), .op(n5815) );
  nand2_1 U8246 ( .ip1(n5769), .ip2(i_ssi_U_dff_tx_mem[80]), .op(n5814) );
  nand2_1 U8247 ( .ip1(n6029), .ip2(i_ssi_U_dff_tx_mem[112]), .op(n5813) );
  nand4_1 U8248 ( .ip1(n5816), .ip2(n5815), .ip3(n5814), .ip4(n5813), .op(
        n5826) );
  nand2_1 U8249 ( .ip1(n5817), .ip2(i_ssi_U_dff_tx_mem[48]), .op(n5824) );
  nand2_1 U8250 ( .ip1(n5818), .ip2(i_ssi_U_dff_tx_mem[64]), .op(n5823) );
  nand2_1 U8251 ( .ip1(n5819), .ip2(i_ssi_U_dff_tx_mem[16]), .op(n5822) );
  nand2_1 U8252 ( .ip1(n5820), .ip2(i_ssi_U_dff_tx_mem[0]), .op(n5821) );
  nand2_1 U8253 ( .ip1(n10346), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[0]), 
        .op(n5827) );
  nand2_1 U8254 ( .ip1(n5380), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[11]), .op(n5831) );
  nand2_1 U8255 ( .ip1(n5263), .ip2(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[7]), .op(n5830) );
  nand3_1 U8256 ( .ip1(n5832), .ip2(n5831), .ip3(n5830), .op(n5833) );
  or2_1 U8257 ( .ip1(n5360), .ip2(n5838), .op(n5840) );
  nand2_1 U8258 ( .ip1(n5850), .ip2(n5851), .op(n6078) );
  nand2_1 U8259 ( .ip1(n5852), .ip2(n6078), .op(n6085) );
  nor2_1 U8260 ( .ip1(n6168), .ip2(n10340), .op(n5853) );
  inv_1 U8261 ( .ip(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[0]), .op(n10280)
         );
  nor2_1 U8262 ( .ip1(n5859), .ip2(n5860), .op(n4410) );
  and3_1 U8263 ( .ip1(i_apb_penable), .ip2(i_apb_pwrite), .ip3(i_apb_psel_en), 
        .op(n5868) );
  inv_1 U8264 ( .ip(i_apb_paddr[17]), .op(n5862) );
  inv_1 U8265 ( .ip(i_apb_paddr[12]), .op(n5867) );
  nand2_1 U8266 ( .ip1(n9838), .ip2(n11148), .op(n9899) );
  inv_1 U8267 ( .ip(i_ssi_reg_addr[1]), .op(n9820) );
  inv_1 U8268 ( .ip(i_ssi_reg_addr[2]), .op(n6199) );
  nor2_1 U8269 ( .ip1(i_ssi_reg_addr[5]), .ip2(i_ssi_reg_addr[4]), .op(n7778)
         );
  inv_1 U8270 ( .ip(i_ssi_reg_addr[3]), .op(n7607) );
  nand3_1 U8271 ( .ip1(i_ssi_reg_addr[0]), .ip2(n7778), .ip3(n7607), .op(n7802) );
  nand2_1 U8272 ( .ip1(n6051), .ip2(n5873), .op(n5885) );
  inv_1 U8273 ( .ip(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[14]), .op(n10341)
         );
  not_ab_or_c_or_d U8274 ( .ip1(n6131), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[7]), .ip3(n5877), .ip4(n5876), 
        .op(n5878) );
  nand2_1 U8275 ( .ip1(n5878), .ip2(n5436), .op(n5879) );
  nand2_1 U8276 ( .ip1(n6177), .ip2(n5879), .op(n5884) );
  or2_1 U8277 ( .ip1(n5880), .ip2(n6040), .op(n5883) );
  or2_1 U8278 ( .ip1(n5881), .ip2(n5332), .op(n5882) );
  nand4_1 U8279 ( .ip1(n5885), .ip2(n5884), .ip3(n5883), .ip4(n5882), .op(
        n5890) );
  inv_1 U8280 ( .ip(i_ssi_U_shift_U_tx_shifter_load_start_bit_ir), .op(n6072)
         );
  nor2_1 U8281 ( .ip1(n5888), .ip2(n10281), .op(n5889) );
  nand2_1 U8282 ( .ip1(n5889), .ip2(n5890), .op(n6100) );
  nand2_1 U8283 ( .ip1(n5812), .ip2(i_ssi_U_dff_tx_mem[43]), .op(n5895) );
  nand2_1 U8284 ( .ip1(n6028), .ip2(i_ssi_U_dff_tx_mem[107]), .op(n5894) );
  nand2_1 U8285 ( .ip1(n5769), .ip2(i_ssi_U_dff_tx_mem[91]), .op(n5893) );
  nand2_1 U8286 ( .ip1(n6029), .ip2(i_ssi_U_dff_tx_mem[123]), .op(n5892) );
  nand4_1 U8287 ( .ip1(n5895), .ip2(n5894), .ip3(n5893), .ip4(n5892), .op(
        n5901) );
  nand2_1 U8288 ( .ip1(n5817), .ip2(i_ssi_U_dff_tx_mem[59]), .op(n5899) );
  nand2_1 U8289 ( .ip1(n5818), .ip2(i_ssi_U_dff_tx_mem[75]), .op(n5898) );
  nand2_1 U8290 ( .ip1(n5819), .ip2(i_ssi_U_dff_tx_mem[27]), .op(n5897) );
  nand2_1 U8291 ( .ip1(n5820), .ip2(i_ssi_U_dff_tx_mem[11]), .op(n5896) );
  nand4_1 U8292 ( .ip1(n5899), .ip2(n5898), .ip3(n5897), .ip4(n5896), .op(
        n5900) );
  nor2_1 U8293 ( .ip1(n10253), .ip2(n6143), .op(n5903) );
  nand2_1 U8294 ( .ip1(n5812), .ip2(i_ssi_U_dff_tx_mem[41]), .op(n5908) );
  nand2_1 U8295 ( .ip1(n6028), .ip2(i_ssi_U_dff_tx_mem[105]), .op(n5907) );
  nand2_1 U8296 ( .ip1(n5769), .ip2(i_ssi_U_dff_tx_mem[89]), .op(n5906) );
  nand2_1 U8297 ( .ip1(n6029), .ip2(i_ssi_U_dff_tx_mem[121]), .op(n5905) );
  nand4_1 U8298 ( .ip1(n5908), .ip2(n5907), .ip3(n5906), .ip4(n5905), .op(
        n5914) );
  nand2_1 U8299 ( .ip1(n5817), .ip2(i_ssi_U_dff_tx_mem[57]), .op(n5912) );
  nand2_1 U8300 ( .ip1(n5818), .ip2(i_ssi_U_dff_tx_mem[73]), .op(n5911) );
  nand2_1 U8301 ( .ip1(n5819), .ip2(i_ssi_U_dff_tx_mem[25]), .op(n5910) );
  nand2_1 U8302 ( .ip1(n5820), .ip2(i_ssi_U_dff_tx_mem[9]), .op(n5909) );
  nand2_1 U8303 ( .ip1(n5918), .ip2(n5917), .op(n5919) );
  nand2_1 U8304 ( .ip1(n5403), .ip2(n5919), .op(n6049) );
  nand2_1 U8305 ( .ip1(n5812), .ip2(i_ssi_U_dff_tx_mem[38]), .op(n5923) );
  nand2_1 U8306 ( .ip1(n6028), .ip2(i_ssi_U_dff_tx_mem[102]), .op(n5922) );
  nand2_1 U8307 ( .ip1(n5769), .ip2(i_ssi_U_dff_tx_mem[86]), .op(n5921) );
  nand2_1 U8308 ( .ip1(n6029), .ip2(i_ssi_U_dff_tx_mem[118]), .op(n5920) );
  nand4_1 U8309 ( .ip1(n5923), .ip2(n5922), .ip3(n5921), .ip4(n5920), .op(
        n5929) );
  nand2_1 U8310 ( .ip1(n5817), .ip2(i_ssi_U_dff_tx_mem[54]), .op(n5927) );
  nand2_1 U8311 ( .ip1(n5818), .ip2(i_ssi_U_dff_tx_mem[70]), .op(n5926) );
  nand2_1 U8312 ( .ip1(n5819), .ip2(i_ssi_U_dff_tx_mem[22]), .op(n5925) );
  nand2_1 U8313 ( .ip1(n5820), .ip2(i_ssi_U_dff_tx_mem[6]), .op(n5924) );
  nand4_1 U8314 ( .ip1(n5927), .ip2(n5926), .ip3(n5925), .ip4(n5924), .op(
        n5928) );
  nor2_1 U8315 ( .ip1(n10260), .ip2(n6040), .op(n5941) );
  nand2_1 U8316 ( .ip1(n5812), .ip2(i_ssi_U_dff_tx_mem[37]), .op(n5933) );
  nand2_1 U8317 ( .ip1(n6028), .ip2(i_ssi_U_dff_tx_mem[101]), .op(n5932) );
  nand2_1 U8318 ( .ip1(n5769), .ip2(i_ssi_U_dff_tx_mem[85]), .op(n5931) );
  nand2_1 U8319 ( .ip1(n6029), .ip2(i_ssi_U_dff_tx_mem[117]), .op(n5930) );
  nand4_1 U8320 ( .ip1(n5933), .ip2(n5932), .ip3(n5931), .ip4(n5930), .op(
        n5939) );
  nand2_1 U8321 ( .ip1(n5817), .ip2(i_ssi_U_dff_tx_mem[53]), .op(n5937) );
  nand2_1 U8322 ( .ip1(n5818), .ip2(i_ssi_U_dff_tx_mem[69]), .op(n5936) );
  nand2_1 U8323 ( .ip1(n5819), .ip2(i_ssi_U_dff_tx_mem[21]), .op(n5935) );
  nand2_1 U8324 ( .ip1(n5820), .ip2(i_ssi_U_dff_tx_mem[5]), .op(n5934) );
  nor2_1 U8325 ( .ip1(n5940), .ip2(n5941), .op(n5955) );
  nor2_1 U8326 ( .ip1(n6101), .ip2(n6143), .op(n5953) );
  nand2_1 U8327 ( .ip1(n5812), .ip2(i_ssi_U_dff_tx_mem[36]), .op(n5945) );
  nand2_1 U8328 ( .ip1(n6028), .ip2(i_ssi_U_dff_tx_mem[100]), .op(n5944) );
  nand2_1 U8329 ( .ip1(n5769), .ip2(i_ssi_U_dff_tx_mem[84]), .op(n5943) );
  nand2_1 U8330 ( .ip1(n6029), .ip2(i_ssi_U_dff_tx_mem[116]), .op(n5942) );
  nand4_1 U8331 ( .ip1(n5945), .ip2(n5944), .ip3(n5943), .ip4(n5942), .op(
        n5951) );
  nand2_1 U8332 ( .ip1(n5817), .ip2(i_ssi_U_dff_tx_mem[52]), .op(n5949) );
  nand2_1 U8333 ( .ip1(n5818), .ip2(i_ssi_U_dff_tx_mem[68]), .op(n5948) );
  nand2_1 U8334 ( .ip1(n5819), .ip2(i_ssi_U_dff_tx_mem[20]), .op(n5947) );
  nand2_1 U8335 ( .ip1(n5820), .ip2(i_ssi_U_dff_tx_mem[4]), .op(n5946) );
  nand2_1 U8336 ( .ip1(n5954), .ip2(n5955), .op(n5956) );
  nand2_1 U8337 ( .ip1(n5263), .ip2(n5956), .op(n6048) );
  nand2_1 U8338 ( .ip1(n5812), .ip2(i_ssi_U_dff_tx_mem[33]), .op(n5960) );
  nand2_1 U8339 ( .ip1(n6028), .ip2(i_ssi_U_dff_tx_mem[97]), .op(n5959) );
  nand2_1 U8340 ( .ip1(n5769), .ip2(i_ssi_U_dff_tx_mem[81]), .op(n5958) );
  nand2_1 U8341 ( .ip1(n6029), .ip2(i_ssi_U_dff_tx_mem[113]), .op(n5957) );
  nand4_1 U8342 ( .ip1(n5960), .ip2(n5959), .ip3(n5958), .ip4(n5957), .op(
        n5966) );
  nand2_1 U8343 ( .ip1(n5817), .ip2(i_ssi_U_dff_tx_mem[49]), .op(n5964) );
  nand2_1 U8344 ( .ip1(n5818), .ip2(i_ssi_U_dff_tx_mem[65]), .op(n5963) );
  nand2_1 U8345 ( .ip1(n5819), .ip2(i_ssi_U_dff_tx_mem[17]), .op(n5962) );
  nand2_1 U8346 ( .ip1(n5820), .ip2(i_ssi_U_dff_tx_mem[1]), .op(n5961) );
  inv_1 U8347 ( .ip(n5458), .op(n5967) );
  nand2_1 U8348 ( .ip1(n5812), .ip2(i_ssi_U_dff_tx_mem[35]), .op(n5973) );
  nand2_1 U8349 ( .ip1(n6028), .ip2(i_ssi_U_dff_tx_mem[99]), .op(n5972) );
  nand2_1 U8350 ( .ip1(n5769), .ip2(i_ssi_U_dff_tx_mem[83]), .op(n5971) );
  nand2_1 U8351 ( .ip1(n6029), .ip2(i_ssi_U_dff_tx_mem[115]), .op(n5970) );
  nand4_1 U8352 ( .ip1(n5973), .ip2(n5972), .ip3(n5971), .ip4(n5970), .op(
        n5979) );
  nand2_1 U8353 ( .ip1(n5817), .ip2(i_ssi_U_dff_tx_mem[51]), .op(n5977) );
  nand2_1 U8354 ( .ip1(n5818), .ip2(i_ssi_U_dff_tx_mem[67]), .op(n5976) );
  nand2_1 U8355 ( .ip1(n5819), .ip2(i_ssi_U_dff_tx_mem[19]), .op(n5975) );
  nand2_1 U8356 ( .ip1(n5820), .ip2(i_ssi_U_dff_tx_mem[3]), .op(n5974) );
  nand4_1 U8357 ( .ip1(n5977), .ip2(n5976), .ip3(n5975), .ip4(n5974), .op(
        n5978) );
  nand2_1 U8358 ( .ip1(n5812), .ip2(i_ssi_U_dff_tx_mem[34]), .op(n5983) );
  nand2_1 U8359 ( .ip1(n6028), .ip2(i_ssi_U_dff_tx_mem[98]), .op(n5982) );
  nand2_1 U8360 ( .ip1(n5769), .ip2(i_ssi_U_dff_tx_mem[82]), .op(n5981) );
  nand2_1 U8361 ( .ip1(n6029), .ip2(i_ssi_U_dff_tx_mem[114]), .op(n5980) );
  nand4_1 U8362 ( .ip1(n5983), .ip2(n5982), .ip3(n5981), .ip4(n5980), .op(
        n5989) );
  nand2_1 U8363 ( .ip1(n5817), .ip2(i_ssi_U_dff_tx_mem[50]), .op(n5987) );
  nand2_1 U8364 ( .ip1(n5818), .ip2(i_ssi_U_dff_tx_mem[66]), .op(n5986) );
  nand2_1 U8365 ( .ip1(n5819), .ip2(i_ssi_U_dff_tx_mem[18]), .op(n5985) );
  nand2_1 U8366 ( .ip1(n5820), .ip2(i_ssi_U_dff_tx_mem[2]), .op(n5984) );
  nand2_1 U8367 ( .ip1(n5992), .ip2(n5993), .op(n5995) );
  inv_1 U8368 ( .ip(n5334), .op(n5994) );
  nand2_1 U8369 ( .ip1(n5995), .ip2(n5994), .op(n6047) );
  nand2_1 U8370 ( .ip1(n5812), .ip2(i_ssi_U_dff_tx_mem[47]), .op(n5999) );
  nand2_1 U8371 ( .ip1(n6028), .ip2(i_ssi_U_dff_tx_mem[111]), .op(n5998) );
  nand2_1 U8372 ( .ip1(n5769), .ip2(i_ssi_U_dff_tx_mem[95]), .op(n5997) );
  nand2_1 U8373 ( .ip1(n6029), .ip2(i_ssi_U_dff_tx_mem[127]), .op(n5996) );
  nand4_1 U8374 ( .ip1(n5999), .ip2(n5998), .ip3(n5997), .ip4(n5996), .op(
        n6005) );
  nand2_1 U8375 ( .ip1(n5817), .ip2(i_ssi_U_dff_tx_mem[63]), .op(n6003) );
  nand2_1 U8376 ( .ip1(n5818), .ip2(i_ssi_U_dff_tx_mem[79]), .op(n6002) );
  nand2_1 U8377 ( .ip1(n5819), .ip2(i_ssi_U_dff_tx_mem[31]), .op(n6001) );
  nand2_1 U8378 ( .ip1(n5820), .ip2(i_ssi_U_dff_tx_mem[15]), .op(n6000) );
  nand4_1 U8379 ( .ip1(n6003), .ip2(n6002), .ip3(n6001), .ip4(n6000), .op(
        n6004) );
  nor2_1 U8380 ( .ip1(n10342), .ip2(n6143), .op(n6017) );
  nand2_1 U8381 ( .ip1(n5812), .ip2(i_ssi_U_dff_tx_mem[44]), .op(n6009) );
  nand2_1 U8382 ( .ip1(n6028), .ip2(i_ssi_U_dff_tx_mem[108]), .op(n6008) );
  nand2_1 U8383 ( .ip1(n5769), .ip2(i_ssi_U_dff_tx_mem[92]), .op(n6007) );
  nand2_1 U8384 ( .ip1(n6029), .ip2(i_ssi_U_dff_tx_mem[124]), .op(n6006) );
  nand4_1 U8385 ( .ip1(n6009), .ip2(n6008), .ip3(n6007), .ip4(n6006), .op(
        n6015) );
  nand2_1 U8386 ( .ip1(n5817), .ip2(i_ssi_U_dff_tx_mem[60]), .op(n6013) );
  nand2_1 U8387 ( .ip1(n5818), .ip2(i_ssi_U_dff_tx_mem[76]), .op(n6012) );
  nand2_1 U8388 ( .ip1(n5819), .ip2(i_ssi_U_dff_tx_mem[28]), .op(n6011) );
  nand2_1 U8389 ( .ip1(n5820), .ip2(i_ssi_U_dff_tx_mem[12]), .op(n6010) );
  nand2_1 U8390 ( .ip1(n5812), .ip2(i_ssi_U_dff_tx_mem[45]), .op(n6021) );
  nand2_1 U8391 ( .ip1(n6028), .ip2(i_ssi_U_dff_tx_mem[109]), .op(n6020) );
  nand2_1 U8392 ( .ip1(n5769), .ip2(i_ssi_U_dff_tx_mem[93]), .op(n6019) );
  nand2_1 U8393 ( .ip1(n6029), .ip2(i_ssi_U_dff_tx_mem[125]), .op(n6018) );
  nand4_1 U8394 ( .ip1(n6021), .ip2(n6020), .ip3(n6019), .ip4(n6018), .op(
        n6027) );
  nand2_1 U8395 ( .ip1(n5817), .ip2(i_ssi_U_dff_tx_mem[61]), .op(n6025) );
  nand2_1 U8396 ( .ip1(n5818), .ip2(i_ssi_U_dff_tx_mem[77]), .op(n6024) );
  nand2_1 U8397 ( .ip1(n5819), .ip2(i_ssi_U_dff_tx_mem[29]), .op(n6023) );
  nand2_1 U8398 ( .ip1(n5820), .ip2(i_ssi_U_dff_tx_mem[13]), .op(n6022) );
  nand2_1 U8399 ( .ip1(n5812), .ip2(i_ssi_U_dff_tx_mem[46]), .op(n6033) );
  nand2_1 U8400 ( .ip1(n6028), .ip2(i_ssi_U_dff_tx_mem[110]), .op(n6032) );
  nand2_1 U8401 ( .ip1(n5769), .ip2(i_ssi_U_dff_tx_mem[94]), .op(n6031) );
  nand2_1 U8402 ( .ip1(n6029), .ip2(i_ssi_U_dff_tx_mem[126]), .op(n6030) );
  nand4_1 U8403 ( .ip1(n6033), .ip2(n6032), .ip3(n6031), .ip4(n6030), .op(
        n6039) );
  nand2_1 U8404 ( .ip1(n5817), .ip2(i_ssi_U_dff_tx_mem[62]), .op(n6037) );
  nand2_1 U8405 ( .ip1(n5818), .ip2(i_ssi_U_dff_tx_mem[78]), .op(n6036) );
  nand2_1 U8406 ( .ip1(n5819), .ip2(i_ssi_U_dff_tx_mem[30]), .op(n6035) );
  nand2_1 U8407 ( .ip1(n5820), .ip2(i_ssi_U_dff_tx_mem[14]), .op(n6034) );
  nand2_1 U8408 ( .ip1(n6044), .ip2(n6043), .op(n6045) );
  nand2_1 U8409 ( .ip1(n5264), .ip2(n6045), .op(n6046) );
  nand4_1 U8410 ( .ip1(n6048), .ip2(n6046), .ip3(n6049), .ip4(n6047), .op(
        n6050) );
  nand2_1 U8411 ( .ip1(n5891), .ip2(n6050), .op(n6099) );
  nand2_1 U8412 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_buffer[15]), .ip2(n10349), 
        .op(n6055) );
  nand2_1 U8413 ( .ip1(n6051), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[13]), 
        .op(n6053) );
  nand4_1 U8414 ( .ip1(n6055), .ip2(n6054), .ip3(n6053), .ip4(n6052), .op(
        n6058) );
  or2_1 U8415 ( .ip1(i_ssi_U_shift_U_tx_shifter_load_start_bit_ir), .ip2(n6056), .op(n6075) );
  nor2_1 U8416 ( .ip1(n6075), .ip2(n5300), .op(n6057) );
  nand2_1 U8417 ( .ip1(n6057), .ip2(n6058), .op(n6069) );
  or2_1 U8418 ( .ip1(n6059), .ip2(n5331), .op(n6065) );
  nor2_1 U8419 ( .ip1(n6075), .ip2(n5839), .op(n6066) );
  nand2_1 U8420 ( .ip1(n6066), .ip2(n6067), .op(n6068) );
  nand2_1 U8421 ( .ip1(n6069), .ip2(n6068), .op(n6097) );
  nor2_1 U8422 ( .ip1(n5334), .ip2(n6075), .op(n6071) );
  nand3_1 U8423 ( .ip1(n10281), .ip2(i_ssi_txd), .ip3(n6072), .op(n6074) );
  nand2_1 U8424 ( .ip1(i_ssi_U_shift_U_tx_shifter_load_start_bit_ir), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[15]), .op(n6073) );
  and2_1 U8425 ( .ip1(n6074), .ip2(n6073), .op(n6094) );
  inv_1 U8426 ( .ip(n5380), .op(n6076) );
  nor2_1 U8427 ( .ip1(n6076), .ip2(n6075), .op(n6092) );
  inv_1 U8428 ( .ip(i_ssi_U_shift_U_tx_shifter_tx_buffer[10]), .op(n6080) );
  nand2_1 U8429 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_buffer[8]), .ip2(n5261), 
        .op(n6086) );
  nand2_1 U8430 ( .ip1(n10349), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[11]), 
        .op(n6089) );
  nand3_1 U8431 ( .ip1(n6100), .ip2(n6098), .ip3(n6099), .op(n4395) );
  or2_1 U8432 ( .ip1(n6101), .ip2(n5279), .op(n6104) );
  nand2_1 U8433 ( .ip1(n9708), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[7]), 
        .op(n6103) );
  nand2_1 U8434 ( .ip1(n9714), .ip2(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[6]), .op(n6102) );
  nand4_1 U8435 ( .ip1(n6104), .ip2(n9717), .ip3(n6103), .ip4(n6102), .op(
        n6108) );
  inv_1 U8436 ( .ip(n5363), .op(n6105) );
  inv_1 U8437 ( .ip(n6111), .op(n6112) );
  nor2_1 U8438 ( .ip1(n6112), .ip2(n9708), .op(n6113) );
  nand2_1 U8439 ( .ip1(n6176), .ip2(n5261), .op(n6123) );
  or2_1 U8440 ( .ip1(n10260), .ip2(n5279), .op(n6121) );
  nand2_1 U8441 ( .ip1(n10346), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[6]), 
        .op(n6120) );
  nand2_1 U8442 ( .ip1(n9714), .ip2(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[5]), .op(n6119) );
  nand4_1 U8443 ( .ip1(n6121), .ip2(n9717), .ip3(n6120), .ip4(n6119), .op(
        n6122) );
  nand2_1 U8444 ( .ip1(n6123), .ip2(n6208), .op(n6124) );
  nand2_1 U8445 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[6]), .ip2(n6124), .op(n6125) );
  nand2_1 U8446 ( .ip1(n6126), .ip2(n6125), .op(n4404) );
  or2_1 U8447 ( .ip1(n10254), .ip2(n5279), .op(n6129) );
  nand2_1 U8448 ( .ip1(n10346), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[12]), 
        .op(n6128) );
  nand2_1 U8449 ( .ip1(n9714), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[11]), .op(n6127) );
  nand4_1 U8450 ( .ip1(n6129), .ip2(n9717), .ip3(n6128), .ip4(n6127), .op(
        n6133) );
  nand2_1 U8451 ( .ip1(n5380), .ip2(n6130), .op(n6132) );
  mux2_1 U8452 ( .ip1(n6133), .ip2(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[12]), .s(n5342), .op(n4398) );
  inv_1 U8453 ( .ip(i_ssi_U_mstfsm_spi1_control), .op(n6134) );
  nand2_1 U8454 ( .ip1(n6135), .ip2(i_ssi_tmod[0]), .op(n6136) );
  nand2_1 U8455 ( .ip1(n6137), .ip2(n8378), .op(n6138) );
  inv_1 U8456 ( .ip(i_ssi_ctrlr0[11]), .op(n9683) );
  nand2_1 U8457 ( .ip1(n10346), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[11]), 
        .op(n6148) );
  nand2_1 U8458 ( .ip1(n9714), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[10]), .op(n6147) );
  nand4_1 U8459 ( .ip1(n6149), .ip2(n9717), .ip3(n6148), .ip4(n6147), .op(
        n6150) );
  nand2_1 U8460 ( .ip1(n5369), .ip2(n6150), .op(n6151) );
  nand2_1 U8461 ( .ip1(n5424), .ip2(n6151), .op(n4399) );
  nand2_1 U8462 ( .ip1(n10346), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[9]), 
        .op(n6158) );
  nand2_1 U8463 ( .ip1(n9714), .ip2(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[8]), .op(n6157) );
  nand4_1 U8464 ( .ip1(n6159), .ip2(n9717), .ip3(n6158), .ip4(n6157), .op(
        n6160) );
  inv_1 U8465 ( .ip(n5342), .op(n6171) );
  nand2_1 U8466 ( .ip1(n10346), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[13]), 
        .op(n6166) );
  nand2_1 U8467 ( .ip1(n9714), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[12]), .op(n6165) );
  nand4_1 U8468 ( .ip1(n6167), .ip2(n9717), .ip3(n6166), .ip4(n6165), .op(
        n6170) );
  nor2_1 U8469 ( .ip1(n6168), .ip2(n10350), .op(n6169) );
  nand2_1 U8470 ( .ip1(n5342), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[13]), .op(n6174) );
  nand3_1 U8471 ( .ip1(n6173), .ip2(n6175), .ip3(n6174), .op(n4397) );
  or2_1 U8472 ( .ip1(n10258), .ip2(n5279), .op(n6180) );
  nand2_1 U8473 ( .ip1(n10346), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[5]), 
        .op(n6179) );
  nand2_1 U8474 ( .ip1(n9714), .ip2(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[4]), .op(n6178) );
  nand4_1 U8475 ( .ip1(n6180), .ip2(n9717), .ip3(n6179), .ip4(n6178), .op(
        n6181) );
  nand2_1 U8476 ( .ip1(n5428), .ip2(n6208), .op(n6187) );
  inv_1 U8477 ( .ip(n6182), .op(n6183) );
  nand3_1 U8478 ( .ip1(n6144), .ip2(n6184), .ip3(n6183), .op(n6185) );
  nand2_1 U8479 ( .ip1(n6185), .ip2(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[5]), .op(n6186) );
  nand2_1 U8480 ( .ip1(n6187), .ip2(n6186), .op(n4405) );
  nand2_1 U8481 ( .ip1(n10346), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[14]), 
        .op(n6191) );
  nand2_1 U8482 ( .ip1(n9714), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[13]), .op(n6190) );
  nand4_1 U8483 ( .ip1(n6192), .ip2(n9717), .ip3(n6191), .ip4(n6190), .op(
        n6193) );
  nand2_1 U8484 ( .ip1(n5268), .ip2(n5427), .op(n6196) );
  nand2_1 U8485 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[14]), .ip2(
        n6196), .op(n6197) );
  nand2_1 U8486 ( .ip1(n6197), .ip2(n6198), .op(n4411) );
  nand2_1 U8487 ( .ip1(n6199), .ip2(i_ssi_reg_addr[1]), .op(n7783) );
  inv_1 U8488 ( .ip(n9817), .op(n6200) );
  nand2_1 U8489 ( .ip1(n6200), .ip2(i_apb_pwdata_int[1]), .op(n6202) );
  nand2_1 U8490 ( .ip1(n9817), .ip2(n5376), .op(n6201) );
  nand2_1 U8491 ( .ip1(n6202), .ip2(n6201), .op(n4636) );
  or2_1 U8492 ( .ip1(n10248), .ip2(n5279), .op(n6205) );
  nand2_1 U8493 ( .ip1(n10346), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[3]), 
        .op(n6204) );
  nand2_1 U8494 ( .ip1(n9714), .ip2(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[2]), .op(n6203) );
  nand4_1 U8495 ( .ip1(n6205), .ip2(n9717), .ip3(n6204), .ip4(n6203), .op(
        n6206) );
  inv_1 U8496 ( .ip(i_ssi_U_sclkgen_ssi_cnt[11]), .op(n10461) );
  inv_1 U8497 ( .ip(n6238), .op(n11652) );
  nor2_1 U8498 ( .ip1(n5257), .ip2(n11652), .op(n6267) );
  nand2_1 U8499 ( .ip1(n6231), .ip2(n6216), .op(n6220) );
  inv_1 U8500 ( .ip(i_ssi_U_sclkgen_ssi_cnt[12]), .op(n10465) );
  inv_1 U8501 ( .ip(i_ssi_baudr[13]), .op(n6223) );
  inv_1 U8502 ( .ip(n6232), .op(n6233) );
  nand2_1 U8503 ( .ip1(n10395), .ip2(n6238), .op(n10378) );
  xor2_1 U8504 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[3]), .ip2(i_ssi_baudr[4]), .op(
        n10321) );
  inv_1 U8505 ( .ip(i_ssi_U_sclkgen_ssi_cnt[2]), .op(n10433) );
  buf_1 U8506 ( .ip(i_ssi_baudr[1]), .op(n10385) );
  xor2_1 U8507 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[0]), .ip2(n10385), .op(n10323)
         );
  nor2_1 U8508 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[15]), .ip2(n11148), .op(n6245)
         );
  inv_1 U8509 ( .ip(i_ssi_U_sclkgen_ssi_cnt[1]), .op(n10416) );
  buf_1 U8510 ( .ip(i_ssi_baudr[2]), .op(n10384) );
  fulladder U8511 ( .a(i_ssi_U_sclkgen_ssi_cnt[1]), .b(n10385), .ci(n10384), 
        .s(n6244) );
  inv_1 U8512 ( .ip(n6248), .op(n6263) );
  xor2_1 U8513 ( .ip1(n6263), .ip2(i_ssi_baudr[5]), .op(n6249) );
  xor2_2 U8514 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[4]), .ip2(n6249), .op(n6250) );
  nand2_1 U8515 ( .ip1(n6252), .ip2(n6251), .op(n6256) );
  nand2_1 U8516 ( .ip1(n5267), .ip2(n6240), .op(n10382) );
  nor2_1 U8517 ( .ip1(i_ssi_baudr[5]), .ip2(i_ssi_baudr[6]), .op(n9088) );
  xnor2_1 U8518 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[6]), .ip2(n6254), .op(n6255) );
  nor2_1 U8519 ( .ip1(n6256), .ip2(n6255), .op(n6257) );
  nand3_1 U8520 ( .ip1(n5415), .ip2(n6239), .ip3(n6257), .op(n6280) );
  inv_1 U8521 ( .ip(i_ssi_baudr[5]), .op(n6259) );
  xor2_1 U8522 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[5]), .ip2(i_ssi_baudr[6]), .op(
        n10322) );
  inv_1 U8523 ( .ip(i_ssi_U_sclkgen_ssi_cnt[8]), .op(n10453) );
  xor2_2 U8524 ( .ip1(n10453), .ip2(n6260), .op(n6276) );
  inv_1 U8525 ( .ip(i_ssi_U_sclkgen_ssi_cnt[7]), .op(n10449) );
  xor2_1 U8526 ( .ip1(n10449), .ip2(n6265), .op(n6266) );
  xor2_1 U8527 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[14]), .ip2(i_ssi_baudr[15]), 
        .op(n10320) );
  xor2_1 U8528 ( .ip1(n10320), .ip2(n6272), .op(n6273) );
  nand2_4 U8529 ( .ip1(n6266), .ip2(n6273), .op(n6274) );
  inv_1 U8530 ( .ip(n6274), .op(n6275) );
  nand2_1 U8531 ( .ip1(n6258), .ip2(n6278), .op(n6279) );
  nor2_1 U8532 ( .ip1(n6280), .ip2(n6279), .op(i_ssi_U_sclkgen_N74) );
  and2_1 U8533 ( .ip1(n6282), .ip2(n6281), .op(n8381) );
  nand2_1 U8534 ( .ip1(n8381), .ip2(n6283), .op(n6286) );
  nand2_1 U8535 ( .ip1(n6284), .ip2(n9057), .op(n6285) );
  nand3_1 U8536 ( .ip1(i_ssi_U_mstfsm_frame_cnt[9]), .ip2(
        i_ssi_U_mstfsm_frame_cnt[8]), .ip3(i_ssi_U_mstfsm_frame_cnt[7]), .op(
        n6288) );
  nand4_1 U8537 ( .ip1(i_ssi_U_mstfsm_frame_cnt[6]), .ip2(
        i_ssi_U_mstfsm_frame_cnt[5]), .ip3(i_ssi_U_mstfsm_frame_cnt[3]), .ip4(
        i_ssi_U_mstfsm_frame_cnt[4]), .op(n10514) );
  inv_2 U8538 ( .ip(i_ssi_dfs[2]), .op(n11547) );
  inv_1 U8539 ( .ip(i_ssi_U_mstfsm_bit_cnt[4]), .op(n9366) );
  nand2_1 U8540 ( .ip1(i_ssi_U_mstfsm_bit_cnt[1]), .ip2(
        i_ssi_U_mstfsm_bit_cnt[2]), .op(n6290) );
  nand2_1 U8541 ( .ip1(n6290), .ip2(n5358), .op(n6291) );
  inv_1 U8542 ( .ip(i_ssi_U_mstfsm_bit_cnt[3]), .op(n10482) );
  nand2_1 U8543 ( .ip1(n6292), .ip2(n10482), .op(n6296) );
  inv_1 U8544 ( .ip(i_ssi_U_mstfsm_bit_cnt[1]), .op(n10475) );
  nor2_1 U8545 ( .ip1(i_ssi_dfs[2]), .ip2(n10475), .op(n6293) );
  nand2_1 U8546 ( .ip1(n6294), .ip2(i_ssi_U_mstfsm_bit_cnt[3]), .op(n6295) );
  and3_1 U8547 ( .ip1(i_ssi_U_mstfsm_spi1_control), .ip2(i_ssi_tmod[0]), .ip3(
        n5281), .op(n10484) );
  nand3_1 U8548 ( .ip1(i_ssi_U_mstfsm_frame_cnt[2]), .ip2(
        i_ssi_U_mstfsm_frame_cnt[1]), .ip3(i_ssi_U_mstfsm_frame_cnt[0]), .op(
        n6299) );
  or2_1 U8549 ( .ip1(n10536), .ip2(n6305), .op(n6307) );
  nand3_1 U8550 ( .ip1(n6308), .ip2(n6307), .ip3(n6306), .op(n6309) );
  nor2_1 U8551 ( .ip1(i_i2c_scl_hcnt_en), .ip2(i_i2c_rx_scl_hcnt_en), .op(
        n6341) );
  inv_1 U8552 ( .ip(i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv), .op(n6897) );
  inv_1 U8553 ( .ip(i_i2c_U_DW_apb_i2c_mstfsm_N252), .op(n6937) );
  nor2_1 U8554 ( .ip1(i_i2c_ic_tar[10]), .ip2(n6937), .op(n6619) );
  inv_1 U8555 ( .ip(i_i2c_mst_debug_cstate[1]), .op(n6867) );
  inv_1 U8556 ( .ip(n6310), .op(n6311) );
  nand2_1 U8557 ( .ip1(i_i2c_mst_debug_cstate[0]), .ip2(n6905), .op(n6913) );
  inv_1 U8558 ( .ip(i_i2c_mst_debug_cstate[2]), .op(n6702) );
  nor2_1 U8559 ( .ip1(i_i2c_mst_debug_cstate[4]), .ip2(n6702), .op(n6468) );
  nand2_1 U8560 ( .ip1(i_i2c_mst_debug_cstate[1]), .ip2(n6468), .op(n6695) );
  nor2_1 U8561 ( .ip1(i_i2c_mst_debug_cstate[0]), .ip2(n6695), .op(n6312) );
  ab_or_c_or_d U8562 ( .ip1(n6619), .ip2(n6469), .ip3(n6880), .ip4(n6312), 
        .op(n6313) );
  nor2_1 U8563 ( .ip1(i_i2c_mst_debug_cstate[3]), .ip2(n10413), .op(n9740) );
  nand2_1 U8564 ( .ip1(n6618), .ip2(n9725), .op(n6314) );
  inv_1 U8565 ( .ip(i_i2c_ic_fs_sync), .op(n7716) );
  inv_1 U8566 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_scl_clk_int), .op(n6315) );
  nor3_4 U8567 ( .ip1(i_i2c_ic_fs_sync), .ip2(
        i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv), .ip3(n7384), .op(n7410) );
  inv_1 U8568 ( .ip(i_i2c_ic_fs_spklen[4]), .op(n6487) );
  inv_1 U8569 ( .ip(i_i2c_ic_fs_spklen[3]), .op(n6321) );
  inv_1 U8570 ( .ip(i_i2c_ic_fs_spklen[1]), .op(n8004) );
  inv_1 U8571 ( .ip(i_i2c_ic_fs_spklen[6]), .op(n7100) );
  nand2_1 U8572 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[6]), 
        .ip2(n7100), .op(n7393) );
  nor4_2 U8573 ( .ip1(n7410), .ip2(n7400), .ip3(n7396), .ip4(n6320), .op(n6328) );
  nor2_1 U8574 ( .ip1(n7394), .ip2(n7389), .op(n6327) );
  inv_1 U8575 ( .ip(i_i2c_ic_fs_spklen[2]), .op(n7118) );
  nor2_1 U8576 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[2]), 
        .ip2(n7118), .op(n6323) );
  nor2_2 U8577 ( .ip1(n5314), .ip2(n8004), .op(n7387) );
  nor4_2 U8578 ( .ip1(n7387), .ip2(n7404), .ip3(n6325), .ip4(n6324), .op(n6326) );
  nand4_1 U8579 ( .ip1(n6328), .ip2(n6327), .ip3(n7398), .ip4(n6326), .op(
        n6339) );
  inv_1 U8580 ( .ip(i_i2c_ic_hs_spklen[2]), .op(n7117) );
  not_ab_or_c_or_d U8581 ( .ip1(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[2]), .ip2(n7117), .ip3(
        n6329), .ip4(n7370), .op(n7375) );
  inv_1 U8582 ( .ip(i_i2c_ic_hs_spklen[7]), .op(n6507) );
  inv_1 U8583 ( .ip(i_i2c_ic_hs_spklen[6]), .op(n7099) );
  nor2_1 U8584 ( .ip1(n5316), .ip2(n7099), .op(n6330) );
  or2_1 U8585 ( .ip1(n6331), .ip2(n6330), .op(n7381) );
  nand2_1 U8586 ( .ip1(i_i2c_ic_hs_spklen[3]), .ip2(n10554), .op(n6333) );
  nand2_1 U8587 ( .ip1(i_i2c_ic_hs_spklen[2]), .ip2(n10552), .op(n6332) );
  nand2_1 U8588 ( .ip1(n6333), .ip2(n6332), .op(n7368) );
  nor2_1 U8589 ( .ip1(n7381), .ip2(n7368), .op(n6337) );
  nand2_1 U8590 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[6]), 
        .ip2(n7099), .op(n6334) );
  inv_1 U8591 ( .ip(i_i2c_ic_hs_spklen[5]), .op(n6515) );
  nand3_1 U8592 ( .ip1(n7375), .ip2(n6337), .ip3(n6336), .op(n6338) );
  nor2_2 U8593 ( .ip1(n5437), .ip2(n6463), .op(n6344) );
  or2_1 U8594 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_hcnt_cmplt_int), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_int_d), .op(n6340) );
  nand3_1 U8595 ( .ip1(i_i2c_mst_tx_ack_vld), .ip2(i_i2c_scl_lcnt_cmplt), 
        .ip3(n6340), .op(n6342) );
  inv_1 U8596 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_hcnt_cmplt_int), .op(n6465)
         );
  nor2_2 U8597 ( .ip1(n6344), .ip2(n6343), .op(n6462) );
  inv_1 U8598 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_data_d_int_0_), 
        .op(n8437) );
  or2_4 U8599 ( .ip1(n6345), .ip2(n5412), .op(n6717) );
  mux2_2 U8600 ( .ip1(i_i2c_ic_fs_hcnt[6]), .ip2(i_i2c_ic_hcnt[6]), .s(n6346), 
        .op(n8023) );
  mux2_2 U8601 ( .ip1(i_i2c_ic_fs_hcnt[5]), .ip2(i_i2c_ic_hcnt[5]), .s(n6717), 
        .op(n8031) );
  mux2_2 U8602 ( .ip1(i_i2c_ic_fs_hcnt[4]), .ip2(i_i2c_ic_hcnt[4]), .s(n6717), 
        .op(n8029) );
  nor2_1 U8603 ( .ip1(n8031), .ip2(n8029), .op(n6416) );
  mux2_2 U8604 ( .ip1(i_i2c_ic_fs_hcnt[1]), .ip2(i_i2c_ic_hcnt[1]), .s(n6717), 
        .op(n8005) );
  mux2_2 U8605 ( .ip1(i_i2c_ic_fs_hcnt[0]), .ip2(i_i2c_ic_hcnt[0]), .s(n6717), 
        .op(n8181) );
  mux2_2 U8606 ( .ip1(i_i2c_ic_fs_hcnt[3]), .ip2(i_i2c_ic_hcnt[3]), .s(n6717), 
        .op(n8010) );
  mux2_2 U8607 ( .ip1(i_i2c_ic_fs_hcnt[2]), .ip2(i_i2c_ic_hcnt[2]), .s(n6717), 
        .op(n8012) );
  nor2_1 U8608 ( .ip1(n8010), .ip2(n8012), .op(n6348) );
  nand2_1 U8609 ( .ip1(n6396), .ip2(n6348), .op(n6390) );
  nor2_1 U8610 ( .ip1(n8065), .ip2(n8100), .op(n6350) );
  inv_1 U8611 ( .ip(n6363), .op(n6351) );
  nand2_1 U8612 ( .ip1(n6376), .ip2(n6351), .op(n6352) );
  inv_1 U8613 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[12]), .op(n6446)
         );
  nor2_1 U8614 ( .ip1(n8003), .ip2(n8070), .op(n6357) );
  inv_1 U8615 ( .ip(n6357), .op(n6353) );
  nor2_1 U8616 ( .ip1(n6363), .ip2(n6353), .op(n6354) );
  nand2_1 U8617 ( .ip1(n6376), .ip2(n6354), .op(n6355) );
  inv_1 U8618 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[14]), .op(n6442)
         );
  nand2_1 U8619 ( .ip1(n6357), .ip2(n8051), .op(n6358) );
  nor2_1 U8620 ( .ip1(n6363), .ip2(n6358), .op(n6359) );
  nand2_1 U8621 ( .ip1(n6376), .ip2(n6359), .op(n6360) );
  inv_1 U8622 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[15]), .op(n6361)
         );
  ab_or_c_or_d U8623 ( .ip1(n6444), .ip2(n6446), .ip3(n6450), .ip4(n6445), 
        .op(n6435) );
  inv_1 U8624 ( .ip(n8039), .op(n6367) );
  nand2_1 U8625 ( .ip1(n6376), .ip2(n6367), .op(n6368) );
  inv_1 U8626 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[8]), .op(n6429)
         );
  xor2_1 U8627 ( .ip1(n6376), .ip2(n8039), .op(n6430) );
  nor2_1 U8628 ( .ip1(n6369), .ip2(n5313), .op(n6371) );
  nor2_1 U8629 ( .ip1(n6369), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[9]), .op(n6370) );
  or2_1 U8630 ( .ip1(n6371), .ip2(n6370), .op(n6381) );
  nand2_1 U8631 ( .ip1(n6376), .ip2(n6373), .op(n6372) );
  inv_1 U8632 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[10]), .op(n6385)
         );
  inv_1 U8633 ( .ip(n6373), .op(n6374) );
  nor2_1 U8634 ( .ip1(n6374), .ip2(n8100), .op(n6375) );
  nand2_1 U8635 ( .ip1(n6376), .ip2(n6375), .op(n6377) );
  inv_1 U8636 ( .ip(n6383), .op(n6379) );
  nor2_1 U8637 ( .ip1(n6381), .ip2(n6428), .op(n6388) );
  inv_1 U8638 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[4]), .op(n6409)
         );
  inv_1 U8639 ( .ip(n6390), .op(n6417) );
  inv_1 U8640 ( .ip(n8029), .op(n6391) );
  nand2_1 U8641 ( .ip1(n6417), .ip2(n6391), .op(n6392) );
  nor2_1 U8642 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[5]), .ip2(n6394), .op(n6408) );
  xor2_1 U8643 ( .ip1(n6417), .ip2(n8029), .op(n6410) );
  inv_1 U8644 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[2]), .op(n6404)
         );
  not_ab_or_c_or_d U8645 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[1]), 
        .ip2(n5420), .ip3(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[0]), .ip4(
        n8181), .op(n6400) );
  nor2_1 U8646 ( .ip1(n5420), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[1]), .op(n6399) );
  nor3_1 U8647 ( .ip1(n6404), .ip2(n6403), .ip3(n6402), .op(n6405) );
  not_ab_or_c_or_d U8648 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[3]), 
        .ip2(n5430), .ip3(n6406), .ip4(n6405), .op(n6407) );
  inv_1 U8649 ( .ip(n6416), .op(n6412) );
  nor2_1 U8650 ( .ip1(n6412), .ip2(n8023), .op(n6413) );
  nand2_1 U8651 ( .ip1(n6413), .ip2(n6417), .op(n6414) );
  nand2_1 U8652 ( .ip1(n6417), .ip2(n6416), .op(n6418) );
  inv_1 U8653 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[6]), .op(n6423)
         );
  nor3_1 U8654 ( .ip1(n6423), .ip2(n6422), .ip3(n6421), .op(n6425) );
  and2_1 U8655 ( .ip1(n6430), .ip2(n6429), .op(n6432) );
  inv_1 U8656 ( .ip(n6439), .op(n6440) );
  nor2_1 U8657 ( .ip1(n6366), .ip2(n6447), .op(n6449) );
  or2_1 U8658 ( .ip1(n6448), .ip2(n6449), .op(n6451) );
  xor2_1 U8659 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[6]), .ip2(n9982), .op(n6460) );
  inv_1 U8660 ( .ip(n6619), .op(n8336) );
  and2_1 U8661 ( .ip1(n6462), .ip2(n6461), .op(n6616) );
  inv_1 U8662 ( .ip(i_i2c_scl_lcnt_cmplt), .op(n11119) );
  nor2_1 U8663 ( .ip1(i_i2c_mst_debug_cstate[3]), .ip2(
        i_i2c_mst_debug_cstate[0]), .op(n6869) );
  nand2_1 U8664 ( .ip1(n6632), .ip2(n6869), .op(n6928) );
  nor2_1 U8665 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_mst_arb_lost), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_slv_arb_lost), .op(n11283) );
  inv_1 U8666 ( .ip(i_i2c_tx_fifo_data_buf[8]), .op(n9096) );
  inv_1 U8667 ( .ip(i_i2c_ack_det), .op(n10582) );
  inv_1 U8668 ( .ip(n6881), .op(n6466) );
  inv_1 U8669 ( .ip(i_i2c_mst_activity), .op(n7080) );
  nand2_1 U8670 ( .ip1(n7080), .ip2(i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_sync_d), 
        .op(n6467) );
  nand3_1 U8671 ( .ip1(n11053), .ip2(i_i2c_ic_abort_sync), .ip3(n6467), .op(
        n9400) );
  nand2_1 U8672 ( .ip1(n6468), .ip2(n6867), .op(n7072) );
  nor2_1 U8673 ( .ip1(n6905), .ip2(n7072), .op(n9724) );
  nand2_1 U8674 ( .ip1(i_i2c_mst_debug_cstate[0]), .ip2(n9724), .op(n6901) );
  nand3_1 U8675 ( .ip1(n9735), .ip2(i_i2c_tx_fifo_data_buf[8]), .ip3(
        i_i2c_U_DW_apb_i2c_sync_ic_rstrt_en_sync_inv), .op(n9402) );
  not_ab_or_c_or_d U8676 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_N487), .ip2(n11110), 
        .ip3(n9401), .ip4(n9403), .op(n6480) );
  nand2_1 U8677 ( .ip1(n6468), .ip2(n6869), .op(n6926) );
  nor2_1 U8678 ( .ip1(n6867), .ip2(n6926), .op(n6694) );
  xor2_1 U8679 ( .ip1(i_i2c_ack_det), .ip2(n8336), .op(n6631) );
  nor2_1 U8680 ( .ip1(n8266), .ip2(n6843), .op(n6899) );
  nor2_1 U8681 ( .ip1(i_i2c_ack_det), .ip2(n8266), .op(n9410) );
  inv_1 U8682 ( .ip(i_i2c_mst_debug_cstate[0]), .op(n7073) );
  inv_1 U8683 ( .ip(n6469), .op(n6470) );
  nand2_1 U8684 ( .ip1(n9410), .ip2(n6471), .op(n6478) );
  mux2_1 U8685 ( .ip1(i_i2c_U_DW_apb_i2c_sync_tx_empty_int_inv), .ip2(
        i_i2c_U_DW_apb_i2c_mstfsm_tx_empty_hld), .s(
        i_i2c_U_DW_apb_i2c_mstfsm_mst_tx_flush), .op(n6473) );
  inv_1 U8686 ( .ip(i_i2c_ic_abort_sync), .op(n6472) );
  nand3_1 U8687 ( .ip1(n6473), .ip2(i_i2c_ic_bus_idle), .ip3(n6472), .op(n6474) );
  nand2_1 U8688 ( .ip1(i_i2c_ic_tar[10]), .ip2(i_i2c_U_DW_apb_i2c_mstfsm_N252), 
        .op(n9188) );
  nand2_1 U8689 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv), .ip2(n9188), 
        .op(n6475) );
  and2_1 U8690 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_rstrt_en_sync_inv), .ip2(
        n6475), .op(n6476) );
  nor2_1 U8691 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv), .ip2(n6476), 
        .op(n6887) );
  inv_1 U8692 ( .ip(n6887), .op(n6477) );
  inv_1 U8693 ( .ip(i_i2c_U_DW_apb_i2c_sync_tx_empty_int_inv), .op(n5245) );
  nor2_1 U8694 ( .ip1(i_i2c_p_det), .ip2(i_i2c_s_det), .op(n8554) );
  inv_1 U8695 ( .ip(i_i2c_slv_debug_cstate[2]), .op(n8527) );
  inv_1 U8696 ( .ip(i_i2c_slv_debug_cstate[3]), .op(n7422) );
  inv_1 U8697 ( .ip(i_i2c_slv_debug_cstate[1]), .op(n7921) );
  inv_1 U8698 ( .ip(i_i2c_slv_debug_cstate[0]), .op(n7922) );
  nor2_1 U8699 ( .ip1(i_i2c_rx_gen_call), .ip2(n8536), .op(n8539) );
  and3_1 U8700 ( .ip1(n8539), .ip2(i_i2c_rx_addr_match), .ip3(
        i_i2c_rx_slv_read), .op(n8302) );
  nand3_1 U8701 ( .ip1(n7422), .ip2(i_i2c_slv_debug_cstate[0]), .ip3(
        i_i2c_slv_debug_cstate[2]), .op(n7634) );
  nand3_1 U8702 ( .ip1(n8294), .ip2(i_i2c_slv_tx_cmplt), .ip3(n6482), .op(
        n9658) );
  nor2_1 U8703 ( .ip1(i_i2c_slv_ack_det), .ip2(n9658), .op(n9657) );
  inv_1 U8704 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_sda_data_int), .op(n6534) );
  inv_1 U8705 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[5]), .op(
        n11276) );
  nor2_1 U8706 ( .ip1(i_i2c_ic_fs_spklen[5]), .ip2(n11276), .op(n6486) );
  or2_1 U8707 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[4]), .ip2(
        n6486), .op(n6489) );
  or2_1 U8708 ( .ip1(n6487), .ip2(n6486), .op(n6488) );
  inv_1 U8709 ( .ip(i_i2c_ic_fs_spklen[0]), .op(n6504) );
  inv_1 U8710 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[3]), .op(
        n11269) );
  nand2_1 U8711 ( .ip1(i_i2c_ic_fs_spklen[3]), .ip2(n11269), .op(n6491) );
  inv_1 U8712 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[2]), .op(
        n11266) );
  nand2_1 U8713 ( .ip1(i_i2c_ic_fs_spklen[2]), .ip2(n11266), .op(n6490) );
  nand2_1 U8714 ( .ip1(n6491), .ip2(n6490), .op(n7640) );
  inv_1 U8715 ( .ip(n7410), .op(n6493) );
  inv_1 U8716 ( .ip(i_i2c_ic_fs_spklen[7]), .op(n7411) );
  nand2_1 U8717 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[7]), 
        .ip2(n7411), .op(n6492) );
  nand2_1 U8718 ( .ip1(n6493), .ip2(n6492), .op(n7650) );
  inv_1 U8719 ( .ip(n7650), .op(n6502) );
  inv_1 U8720 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[4]), .op(
        n11272) );
  and2_1 U8721 ( .ip1(n11276), .ip2(i_i2c_ic_fs_spklen[5]), .op(n7645) );
  nor2_1 U8722 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[6]), 
        .ip2(n7100), .op(n6495) );
  nor2_1 U8723 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[7]), 
        .ip2(n7411), .op(n6494) );
  or2_1 U8724 ( .ip1(n6495), .ip2(n6494), .op(n7646) );
  not_ab_or_c_or_d U8725 ( .ip1(i_i2c_ic_fs_spklen[4]), .ip2(n11272), .ip3(
        n7645), .ip4(n7646), .op(n7653) );
  nor2_1 U8726 ( .ip1(i_i2c_ic_fs_spklen[2]), .ip2(n11266), .op(n6496) );
  or2_1 U8727 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[1]), .ip2(
        n6496), .op(n6498) );
  or2_1 U8728 ( .ip1(n8004), .ip2(n6496), .op(n6497) );
  nand2_1 U8729 ( .ip1(n6498), .ip2(n6497), .op(n7636) );
  nor2_1 U8730 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[1]), 
        .ip2(n8004), .op(n6499) );
  or2_1 U8731 ( .ip1(i_i2c_ic_fs_spklen[0]), .ip2(n6499), .op(n6501) );
  inv_1 U8732 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[0]), .op(
        n11263) );
  or2_1 U8733 ( .ip1(n11263), .ip2(n6499), .op(n6500) );
  nand2_1 U8734 ( .ip1(n6501), .ip2(n6500), .op(n7638) );
  not_ab_or_c_or_d U8735 ( .ip1(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[0]), .ip2(n6504), .ip3(
        n7640), .ip4(n6503), .op(n6505) );
  nand2_1 U8736 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[6]), 
        .ip2(n7100), .op(n7643) );
  or2_1 U8737 ( .ip1(n11269), .ip2(i_i2c_ic_fs_spklen[3]), .op(n7642) );
  inv_1 U8738 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[1]), .op(
        n11262) );
  nor2_1 U8739 ( .ip1(i_i2c_ic_hs_spklen[1]), .ip2(n11262), .op(n6506) );
  nor2_1 U8740 ( .ip1(i_i2c_ic_hs_spklen[3]), .ip2(n11269), .op(n7657) );
  not_ab_or_c_or_d U8741 ( .ip1(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[2]), .ip2(n7117), .ip3(
        n6506), .ip4(n7657), .op(n7655) );
  nor2_1 U8742 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[7]), 
        .ip2(n6507), .op(n7671) );
  and2_1 U8743 ( .ip1(n6507), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[7]), .op(n7666) );
  nand2_1 U8744 ( .ip1(i_i2c_ic_hs_spklen[3]), .ip2(n11269), .op(n6509) );
  nand2_1 U8745 ( .ip1(i_i2c_ic_hs_spklen[2]), .ip2(n11266), .op(n6508) );
  nand2_1 U8746 ( .ip1(n6509), .ip2(n6508), .op(n7659) );
  nand2_1 U8747 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[6]), 
        .ip2(n7099), .op(n6510) );
  nand2_1 U8748 ( .ip1(n7672), .ip2(n6510), .op(n7665) );
  inv_1 U8749 ( .ip(n7665), .op(n6522) );
  nor2_1 U8750 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[5]), 
        .ip2(n6515), .op(n6511) );
  or2_1 U8751 ( .ip1(i_i2c_ic_hs_spklen[6]), .ip2(n6511), .op(n6513) );
  inv_1 U8752 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[6]), .op(
        n11280) );
  or2_1 U8753 ( .ip1(n11280), .ip2(n6511), .op(n6512) );
  nand2_1 U8754 ( .ip1(n6513), .ip2(n6512), .op(n7668) );
  nor2_1 U8755 ( .ip1(i_i2c_ic_hs_spklen[4]), .ip2(n11272), .op(n6514) );
  or2_1 U8756 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[5]), .ip2(
        n6514), .op(n6517) );
  or2_1 U8757 ( .ip1(n6515), .ip2(n6514), .op(n6516) );
  nand2_1 U8758 ( .ip1(n6517), .ip2(n6516), .op(n7664) );
  inv_1 U8759 ( .ip(i_i2c_ic_hs_spklen[1]), .op(n6518) );
  nor2_1 U8760 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[1]), 
        .ip2(n6518), .op(n6519) );
  or2_1 U8761 ( .ip1(i_i2c_ic_hs_spklen[0]), .ip2(n6519), .op(n6521) );
  or2_1 U8762 ( .ip1(n11263), .ip2(n6519), .op(n6520) );
  nand2_1 U8763 ( .ip1(n6521), .ip2(n6520), .op(n7654) );
  inv_1 U8764 ( .ip(i_i2c_ic_hs_spklen[0]), .op(n6524) );
  nand2_1 U8765 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[0]), 
        .ip2(n6524), .op(n6525) );
  nand2_1 U8766 ( .ip1(i_i2c_ic_hs_spklen[4]), .ip2(n11272), .op(n7661) );
  nor4_1 U8767 ( .ip1(n5320), .ip2(n5317), .ip3(n5316), .ip4(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[2]), .op(n6530) );
  nor2_1 U8768 ( .ip1(n5314), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[0]), .op(n7415) );
  inv_1 U8769 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[7]), .op(
        n6529) );
  nand4_1 U8770 ( .ip1(n6530), .ip2(n7415), .ip3(n10554), .ip4(n6529), .op(
        n6531) );
  nand3_1 U8771 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_scl_clk_int), .ip2(n8437), 
        .ip3(n6531), .op(n9404) );
  inv_1 U8772 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_sda_post_hold_done), .op(
        n6536) );
  nor2_1 U8773 ( .ip1(i_i2c_ic_sda_rx_hold_sync[4]), .ip2(n7002), .op(n7001)
         );
  or2_1 U8774 ( .ip1(i_i2c_ic_sda_rx_hold_sync[5]), .ip2(n7005), .op(n7032) );
  nor2_1 U8775 ( .ip1(i_i2c_ic_sda_rx_hold_sync[6]), .ip2(n7032), .op(n7031)
         );
  nor2_1 U8776 ( .ip1(i_i2c_ic_sda_rx_hold_sync[7]), .ip2(n7044), .op(n7046)
         );
  nor2_1 U8777 ( .ip1(n7046), .ip2(n10584), .op(n6535) );
  nand2_1 U8778 ( .ip1(n11776), .ip2(i_i2c_sda_int), .op(n10800) );
  nor2_1 U8779 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_sda_int_q), .ip2(n10800), 
        .op(n11775) );
  or2_1 U8780 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_scl_int_q), .ip2(n10584), 
        .op(n11167) );
  inv_1 U8781 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_hs_mcode_fed_dtctd_r), .op(
        n6537) );
  nor3_1 U8782 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv), .ip2(n11167), 
        .ip3(n6537), .op(n6538) );
  nor2_1 U8783 ( .ip1(n7672), .ip2(n6538), .op(n6539) );
  nor2_1 U8784 ( .ip1(n11775), .ip2(n6539), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_hs) );
  inv_1 U8785 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_scl_int_q), .op(n6541) );
  nor2_1 U8786 ( .ip1(n11776), .ip2(n6541), .op(n11769) );
  inv_1 U8787 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[13]), .op(n6547)
         );
  inv_1 U8788 ( .ip(i_apb_U_DW_apb_ahbsif_state[2]), .op(n10024) );
  nor3_1 U8789 ( .ip1(i_ahb_U_mux_hsel_prev[2]), .ip2(i_ahb_U_mux_hsel_prev[3]), .ip3(i_ahb_U_mux_hsel_prev[4]), .op(n9196) );
  inv_1 U8790 ( .ip(i_ahb_U_mux_hsel_prev[1]), .op(n9195) );
  inv_1 U8791 ( .ip(i_ahb_U_mux_hsel_prev[2]), .op(n11356) );
  inv_1 U8792 ( .ip(i_ahb_U_mux_hsel_prev[3]), .op(n6551) );
  nand2_1 U8793 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hready_resp), .op(
        n6553) );
  nand2_1 U8794 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hready_resp), .op(n6552) );
  inv_1 U8795 ( .ip(n6569), .op(n6568) );
  inv_1 U8796 ( .ip(i_apb_U_DW_apb_ahbsif_state[1]), .op(n9378) );
  inv_1 U8797 ( .ip(i_apb_U_DW_apb_ahbsif_state[0]), .op(n9381) );
  nor3_1 U8798 ( .ip1(n9378), .ip2(n9381), .ip3(i_apb_U_DW_apb_ahbsif_state[2]), .op(n6586) );
  nor2_1 U8799 ( .ip1(i_apb_U_DW_apb_ahbsif_state[0]), .ip2(n9378), .op(n10021) );
  nand2_1 U8800 ( .ip1(i_apb_U_DW_apb_ahbsif_state[2]), .ip2(n10021), .op(
        n6584) );
  or2_1 U8801 ( .ip1(n10106), .ip2(n9379), .op(n6563) );
  inv_1 U8802 ( .ip(ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite), .op(n6561) );
  or2_1 U8803 ( .ip1(n6561), .ip2(n9379), .op(n6562) );
  nand2_1 U8804 ( .ip1(n6563), .ip2(n6562), .op(n6564) );
  not_ab_or_c_or_d U8805 ( .ip1(i_apb_U_DW_apb_ahbsif_pipeline_c), .ip2(n6566), 
        .ip3(n10018), .ip4(n6565), .op(n6567) );
  nor2_1 U8806 ( .ip1(n9381), .ip2(i_apb_U_DW_apb_ahbsif_state[1]), .op(n11367) );
  nor2_1 U8807 ( .ip1(i_apb_pclk_en), .ip2(n9377), .op(n10020) );
  not_ab_or_c_or_d U8808 ( .ip1(n6568), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite), .ip3(n6567), .ip4(n10020), .op(
        n6573) );
  nand3_1 U8809 ( .ip1(n9897), .ip2(n6570), .ip3(n6569), .op(n6571) );
  nand2_1 U8810 ( .ip1(i_apb_pclk_en), .ip2(n6571), .op(n6572) );
  nand2_1 U8811 ( .ip1(i_apb_U_DW_apb_ahbsif_pipeline_c), .ip2(
        i_apb_U_DW_apb_ahbsif_piped_hwrite_c), .op(n6578) );
  not_ab_or_c_or_d U8812 ( .ip1(n6575), .ip2(n6574), .ip3(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite), .ip4(n9379), .op(n6577) );
  inv_1 U8813 ( .ip(i_apb_U_DW_apb_ahbsif_pipeline_c), .op(n10110) );
  nor3_1 U8814 ( .ip1(n10018), .ip2(i_apb_U_DW_apb_ahbsif_piped_hwrite_c), 
        .ip3(n10110), .op(n6576) );
  ab_or_c_or_d U8815 ( .ip1(i_apb_U_DW_apb_ahbsif_state[2]), .ip2(n9378), 
        .ip3(n6577), .ip4(n6576), .op(i_apb_U_DW_apb_ahbsif_nextstate[2]) );
  nand3_1 U8816 ( .ip1(n6580), .ip2(n6579), .ip3(i_apb_pclk_en), .op(n6581) );
  or2_1 U8817 ( .ip1(i_apb_U_DW_apb_ahbsif_nextstate[0]), .ip2(n10105), .op(
        n9384) );
  inv_1 U8818 ( .ip(n6589), .op(n6583) );
  or2_1 U8819 ( .ip1(n9384), .ip2(n6583), .op(n10041) );
  nor2_4 U8820 ( .ip1(n10009), .ip2(i_apb_U_DW_apb_ahbsif_nextstate[2]), .op(
        n10026) );
  nor2_1 U8821 ( .ip1(n6585), .ip2(n6596), .op(n11365) );
  nand2_1 U8822 ( .ip1(n6586), .ip2(i_apb_U_DW_apb_ahbsif_pipeline_c), .op(
        n6587) );
  nand2_1 U8823 ( .ip1(n11365), .ip2(n6587), .op(n10040) );
  nand2_2 U8824 ( .ip1(n10041), .ip2(n10040), .op(n11465) );
  nand2_1 U8825 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[3]), .ip2(n11465), 
        .op(n6594) );
  nand2_1 U8826 ( .ip1(n9384), .ip2(n6596), .op(n6588) );
  nand2_1 U8827 ( .ip1(n6589), .ip2(n6588), .op(n10042) );
  nand2_1 U8828 ( .ip1(n5270), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[3]), 
        .op(n6591) );
  nand2_1 U8829 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[3]), .ip2(n11466), 
        .op(n6590) );
  nand2_1 U8830 ( .ip1(n6591), .ip2(n6590), .op(n6592) );
  inv_1 U8831 ( .ip(n6592), .op(n6593) );
  nand2_1 U8832 ( .ip1(n6594), .ip2(n6593), .op(n4758) );
  nand2_1 U8833 ( .ip1(n10105), .ip2(n10017), .op(n6595) );
  nor2_1 U8834 ( .ip1(i_apb_U_DW_apb_ahbsif_state[2]), .ip2(n9374), .op(n10019) );
  nand2_1 U8835 ( .ip1(i_apb_U_DW_apb_ahbsif_pipeline_c), .ip2(n10019), .op(
        n6597) );
  not_ab_or_c_or_d U8836 ( .ip1(n9377), .ip2(n6597), .ip3(
        i_apb_U_DW_apb_ahbsif_use_saved_data), .ip4(n6596), .op(n9372) );
  xor2_2 U8837 ( .ip1(i_ssi_U_fifo_tx_pop_edge), .ip2(i_ssi_tx_pop), .op(
        i_ssi_tx_pop_sync) );
  and4_1 U8838 ( .ip1(i_ssi_reg_addr[5]), .ip2(i_ssi_reg_addr[3]), .ip3(
        i_ssi_reg_addr[4]), .ip4(i_ssi_reg_addr[2]), .op(n6599) );
  nor2_1 U8839 ( .ip1(i_ssi_reg_addr[5]), .ip2(i_ssi_reg_addr[3]), .op(n6598)
         );
  nor3_1 U8840 ( .ip1(i_ssi_reg_addr[0]), .ip2(i_ssi_reg_addr[5]), .ip3(
        i_ssi_reg_addr[4]), .op(n6600) );
  nand2_1 U8841 ( .ip1(n9838), .ip2(n11567), .op(n9788) );
  inv_1 U8842 ( .ip(n9788), .op(n6602) );
  inv_1 U8843 ( .ip(i_apb_pwdata_int[0]), .op(n6601) );
  nand2_2 U8844 ( .ip1(i_ssi_U_fifo_U_tx_fifo_empty_n), .ip2(i_ssi_tx_pop_sync), .op(n9692) );
  nand2_1 U8845 ( .ip1(i_ssi_tx_full), .ip2(i_ssi_U_fifo_U_tx_fifo_empty_n), 
        .op(n6604) );
  nand2_2 U8846 ( .ip1(n6972), .ip2(n7087), .op(n9071) );
  inv_1 U8847 ( .ip(i_ssi_U_fifo_unconnected_tx_wrd_count[0]), .op(n6606) );
  nand2_2 U8848 ( .ip1(n10052), .ip2(n6606), .op(n10055) );
  nand2_2 U8849 ( .ip1(n10055), .ip2(n6605), .op(n9074) );
  nand2_1 U8850 ( .ip1(n9071), .ip2(n6606), .op(n6607) );
  xor2_2 U8851 ( .ip1(i_ssi_U_fifo_unconnected_tx_wrd_count[1]), .ip2(n6608), 
        .op(n10184) );
  nor2_2 U8852 ( .ip1(n11227), .ip2(n10184), .op(i_ssi_U_fifo_U_tx_fifo_N48)
         );
  inv_1 U8853 ( .ip(i_ssi_U_fifo_unconnected_rx_wrd_count[2]), .op(n6614) );
  inv_1 U8854 ( .ip(i_ssi_U_fifo_unconnected_rx_wrd_count[0]), .op(n6612) );
  inv_1 U8855 ( .ip(i_apb_psel_en), .op(n6609) );
  nor3_1 U8856 ( .ip1(i_apb_penable), .ip2(i_apb_pwrite), .ip3(n6609), .op(
        n7433) );
  inv_1 U8857 ( .ip(n11165), .op(n11782) );
  not_ab_or_c_or_d U8858 ( .ip1(i_ssi_U_fifo_U_rx_fifo_empty_n), .ip2(
        i_ssi_rx_full), .ip3(n11164), .ip4(n5413), .op(n6610) );
  nor2_1 U8859 ( .ip1(n6610), .ip2(n10220), .op(n10225) );
  nor2_1 U8860 ( .ip1(n10223), .ip2(i_ssi_U_fifo_unconnected_rx_wrd_count[1]), 
        .op(n6611) );
  not_ab_or_c_or_d U8861 ( .ip1(i_ssi_U_fifo_unconnected_rx_wrd_count[1]), 
        .ip2(n6612), .ip3(n10225), .ip4(n6611), .op(n6613) );
  nor2_2 U8862 ( .ip1(n11227), .ip2(n6615), .op(i_ssi_U_fifo_U_rx_fifo_N49) );
  xor2_1 U8863 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_rx_push_flg_sync), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_rx_push_flg_sync_q), .op(i_i2c_rx_push_sync)
         );
  nand2_1 U8864 ( .ip1(n9740), .ip2(n8266), .op(n6617) );
  nand2_1 U8865 ( .ip1(n6618), .ip2(n6617), .op(i_i2c_hs_mcode_en) );
  nor2_1 U8866 ( .ip1(n6619), .ip2(n6648), .op(n6626) );
  inv_1 U8867 ( .ip(i_i2c_U_DW_apb_i2c_sync_ic_10bit_mst_sync_inv), .op(n6703)
         );
  nand2_1 U8868 ( .ip1(n6927), .ip2(i_i2c_U_DW_apb_i2c_mstfsm_addr_2byte_sent), 
        .op(n6910) );
  inv_1 U8869 ( .ip(i_i2c_U_DW_apb_i2c_mstfsm_addr_1byte_sent), .op(n6625) );
  nand2_1 U8870 ( .ip1(n6910), .ip2(n6625), .op(n6620) );
  nand2_1 U8871 ( .ip1(n9096), .ip2(n6946), .op(n6621) );
  nor3_1 U8872 ( .ip1(i_i2c_ic_abort_sync), .ip2(n5245), .ip3(n6470), .op(
        n8337) );
  nor2_1 U8873 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_rstrt_en_sync_inv), .ip2(
        n6703), .op(n6623) );
  and2_1 U8874 ( .ip1(n9096), .ip2(n6623), .op(n6624) );
  nor2_1 U8875 ( .ip1(n6913), .ip2(n6695), .op(n8418) );
  nand2_1 U8876 ( .ip1(n8418), .ip2(i_i2c_U_DW_apb_i2c_mstfsm_byte_waiting_q), 
        .op(n11048) );
  nand2_1 U8877 ( .ip1(i_i2c_ic_abort_sync), .ip2(
        i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_chk_win), .op(n8425) );
  nor2_1 U8878 ( .ip1(n6624), .ip2(n8329), .op(n6641) );
  nand2_1 U8879 ( .ip1(i_i2c_scl_lcnt_cmplt), .ip2(i_i2c_scl_p_setup_cmplt), 
        .op(n9997) );
  inv_1 U8880 ( .ip(n6695), .op(n6870) );
  nand2_1 U8881 ( .ip1(i_i2c_mst_debug_cstate[3]), .ip2(n6870), .op(n7075) );
  nor2_1 U8882 ( .ip1(n6874), .ip2(n7075), .op(n6639) );
  nand2_1 U8883 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_10bit_mst_sync_inv), .ip2(
        n6626), .op(n6929) );
  or2_1 U8884 ( .ip1(n6927), .ip2(n6894), .op(n6629) );
  inv_1 U8885 ( .ip(i_i2c_U_DW_apb_i2c_sync_ic_rstrt_en_sync_inv), .op(n6903)
         );
  or2_1 U8886 ( .ip1(n6903), .ip2(n6894), .op(n6628) );
  and2_1 U8887 ( .ip1(i_i2c_scl_s_hld_cmplt), .ip2(i_i2c_scl_s_setup_cmplt), 
        .op(n6941) );
  inv_1 U8888 ( .ip(i_i2c_mst_rxbyte_rdy), .op(n6630) );
  nand2_1 U8889 ( .ip1(n8418), .ip2(n6630), .op(n6636) );
  nand2_1 U8890 ( .ip1(n6880), .ip2(i_i2c_scl_s_hld_cmplt), .op(n6634) );
  nand3_1 U8891 ( .ip1(i_i2c_mst_debug_cstate[3]), .ip2(n6632), .ip3(n7073), 
        .op(n6936) );
  or2_1 U8892 ( .ip1(n6941), .ip2(n6936), .op(n6633) );
  not_ab_or_c_or_d U8893 ( .ip1(i_i2c_ack_det), .ip2(n8337), .ip3(n6641), 
        .ip4(n6640), .op(n6646) );
  nor2_1 U8894 ( .ip1(n6903), .ip2(n9096), .op(n6642) );
  nor2_1 U8895 ( .ip1(n6642), .ip2(n6901), .op(n6846) );
  inv_1 U8896 ( .ip(n6846), .op(n9662) );
  inv_1 U8897 ( .ip(n9448), .op(n9664) );
  nand2_1 U8898 ( .ip1(n9724), .ip2(n7073), .op(n9666) );
  nand2_1 U8899 ( .ip1(n8339), .ip2(n6643), .op(n6645) );
  nand2_1 U8900 ( .ip1(n8266), .ip2(n6845), .op(n6644) );
  not_ab_or_c_or_d U8901 ( .ip1(n6912), .ip2(n6648), .ip3(n6715), .ip4(n6647), 
        .op(n11044) );
  inv_1 U8902 ( .ip(i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv), .op(n9773) );
  or2_1 U8903 ( .ip1(i_i2c_ic_enable_sync), .ip2(i_i2c_mst_activity), .op(
        n6649) );
  nand3_1 U8904 ( .ip1(n11283), .ip2(n9773), .ip3(n6649), .op(n8372) );
  inv_1 U8905 ( .ip(n11227), .op(n11219) );
  nand3_1 U8906 ( .ip1(n11219), .ip2(i_ssi_tx_full), .ip3(n11780), .op(n6650)
         );
  inv_1 U8907 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[1]), .op(n6652)
         );
  nand2_1 U8908 ( .ip1(n6969), .ip2(n6652), .op(n6653) );
  nand2_1 U8909 ( .ip1(n9942), .ip2(n6653), .op(n6654) );
  inv_1 U8910 ( .ip(i_ssi_dfs[1]), .op(n11543) );
  nand2_1 U8911 ( .ip1(n10205), .ip2(n11543), .op(n6656) );
  nand3_1 U8912 ( .ip1(n5266), .ip2(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[2]), .ip3(n6656), .op(n6658) );
  nand2_1 U8913 ( .ip1(n6655), .ip2(i_ssi_rx_push_data[2]), .op(n6657) );
  nand2_1 U8914 ( .ip1(n6658), .ip2(n6657), .op(n4443) );
  nand2_1 U8915 ( .ip1(n6655), .ip2(i_ssi_rx_push_data[1]), .op(n6661) );
  nand3_1 U8916 ( .ip1(n5266), .ip2(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[1]), .ip3(n6659), .op(n6660) );
  nand2_1 U8917 ( .ip1(n6661), .ip2(n6660), .op(n4444) );
  inv_1 U8918 ( .ip(i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[0]), .op(n6678) );
  inv_1 U8919 ( .ip(i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[1]), .op(n6674) );
  inv_1 U8920 ( .ip(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_empty_n), .op(n5247) );
  or2_1 U8921 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[1]), .ip2(n6664), 
        .op(n6666) );
  inv_1 U8922 ( .ip(i_i2c_rx_full), .op(n11180) );
  nand2_1 U8923 ( .ip1(n11209), .ip2(n11180), .op(n11204) );
  nand2_1 U8924 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_empty_n), .ip2(n11204), .op(n6663) );
  nand2_1 U8925 ( .ip1(i_i2c_rx_push_sync), .ip2(n6663), .op(n6669) );
  nand2_1 U8926 ( .ip1(i_i2c_ic_rx_tl[0]), .ip2(i_i2c_ic_rx_tl[1]), .op(n6680)
         );
  inv_1 U8927 ( .ip(i_i2c_ic_rx_tl[2]), .op(n6668) );
  nand2_1 U8928 ( .ip1(n6680), .ip2(n6668), .op(n6690) );
  or2_1 U8929 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[0]), .ip2(n6670), 
        .op(n6672) );
  inv_1 U8930 ( .ip(n6669), .op(n6675) );
  or2_1 U8931 ( .ip1(n6675), .ip2(n6670), .op(n6671) );
  nor2_1 U8932 ( .ip1(i_i2c_rx_push_sync), .ip2(n11205), .op(n6676) );
  nand3_1 U8933 ( .ip1(i_i2c_ic_rx_tl[0]), .ip2(i_i2c_ic_rx_tl[1]), .ip3(
        i_i2c_ic_rx_tl[2]), .op(n11177) );
  nand2_1 U8934 ( .ip1(i_i2c_ic_rx_tl[0]), .ip2(n11177), .op(n6679) );
  nand2_1 U8935 ( .ip1(n6988), .ip2(n6679), .op(n6683) );
  nor2_1 U8936 ( .ip1(n6838), .ip2(n6683), .op(n6685) );
  nor2_1 U8937 ( .ip1(i_i2c_ic_rx_tl[0]), .ip2(i_i2c_ic_rx_tl[1]), .op(n6682)
         );
  nor2_1 U8938 ( .ip1(i_i2c_ic_rx_tl[2]), .ip2(n6680), .op(n6681) );
  not_ab_or_c_or_d U8939 ( .ip1(n6683), .ip2(n6838), .ip3(n6682), .ip4(n6681), 
        .op(n6684) );
  or2_1 U8940 ( .ip1(n6685), .ip2(n6684), .op(n6689) );
  nand2_1 U8941 ( .ip1(n6690), .ip2(n6689), .op(n6692) );
  nand4_1 U8942 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[0]), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[1]), .ip3(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[2]), .ip4(n11209), .op(n6686)
         );
  nand2_1 U8943 ( .ip1(n6686), .ip2(n11180), .op(n6687) );
  nand2_1 U8944 ( .ip1(n6687), .ip2(i_i2c_rx_push_sync), .op(n6688) );
  nand2_1 U8945 ( .ip1(i_i2c_rx_full), .ip2(n11209), .op(n11191) );
  nand2_1 U8946 ( .ip1(n6688), .ip2(n11191), .op(n6839) );
  nor2_1 U8947 ( .ip1(n6690), .ip2(n6689), .op(n6691) );
  ab_or_c_or_d U8948 ( .ip1(n6989), .ip2(n6692), .ip3(n6839), .ip4(n6691), 
        .op(n6693) );
  nand2_1 U8949 ( .ip1(n9725), .ip2(n9737), .op(n6711) );
  nor2_1 U8950 ( .ip1(n7073), .ip2(n6695), .op(n6907) );
  nor2_1 U8951 ( .ip1(n6616), .ip2(n8217), .op(n6697) );
  nor2_1 U8952 ( .ip1(n6941), .ip2(n6881), .op(n6696) );
  not_ab_or_c_or_d U8953 ( .ip1(n6907), .ip2(n9997), .ip3(n6697), .ip4(n6696), 
        .op(n6698) );
  nor2_1 U8954 ( .ip1(n6698), .ip2(n6905), .op(n6710) );
  nand3_1 U8955 ( .ip1(n9096), .ip2(n8425), .ip3(i_i2c_mst_rxbyte_rdy), .op(
        n6902) );
  nor2_1 U8956 ( .ip1(n6902), .ip2(n11048), .op(n6707) );
  nor3_1 U8957 ( .ip1(i_i2c_mst_debug_cstate[0]), .ip2(n6941), .ip3(n7075), 
        .op(n6701) );
  nor3_1 U8958 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_addr_1byte_sent), .ip2(n6888), 
        .ip3(n6928), .op(n6700) );
  inv_1 U8959 ( .ip(i_i2c_mst_debug_cstate[4]), .op(n6868) );
  nor4_1 U8960 ( .ip1(i_i2c_mst_debug_cstate[1]), .ip2(n6868), .ip3(n6913), 
        .ip4(n6702), .op(n6939) );
  inv_1 U8961 ( .ip(i_i2c_U_DW_apb_i2c_mstfsm_N382), .op(n6954) );
  nand4_1 U8962 ( .ip1(n6939), .ip2(i_i2c_scl_s_hld_cmplt), .ip3(n6954), .ip4(
        n6703), .op(n6704) );
  not_ab_or_c_or_d U8963 ( .ip1(n9410), .ip2(n6711), .ip3(n6710), .ip4(n6709), 
        .op(n6714) );
  nand2_1 U8964 ( .ip1(n6846), .ip2(n9667), .op(n6713) );
  nand3_1 U8965 ( .ip1(n9448), .ip2(n8339), .ip3(n9096), .op(n6712) );
  mux2_2 U8966 ( .ip1(i_i2c_ic_fs_lcnt[6]), .ip2(i_i2c_ic_lcnt[6]), .s(n6717), 
        .op(n7965) );
  nand2_1 U8967 ( .ip1(n6716), .ip2(n6782), .op(n6719) );
  mux2_2 U8968 ( .ip1(i_i2c_ic_fs_lcnt[1]), .ip2(i_i2c_ic_lcnt[1]), .s(n6717), 
        .op(n7942) );
  nor2_2 U8969 ( .ip1(n6719), .ip2(n6766), .op(n6764) );
  nor2_2 U8970 ( .ip1(n7979), .ip2(n7938), .op(n6756) );
  inv_1 U8971 ( .ip(n7934), .op(n6723) );
  nand2_1 U8972 ( .ip1(n6728), .ip2(n6723), .op(n6724) );
  nor2_1 U8973 ( .ip1(n6738), .ip2(n6724), .op(n6725) );
  nand2_1 U8974 ( .ip1(n6727), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[15]), .op(n6755) );
  inv_1 U8975 ( .ip(n6728), .op(n6729) );
  nor2_1 U8976 ( .ip1(n6738), .ip2(n6729), .op(n6730) );
  nand2_1 U8977 ( .ip1(n6734), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[14]), .op(n6737) );
  nor2_1 U8978 ( .ip1(n6738), .ip2(n7977), .op(n6732) );
  nand2_1 U8979 ( .ip1(n8730), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[13]), .op(n6735) );
  nor2_2 U8980 ( .ip1(n6734), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[14]), .op(n6748) );
  or2_1 U8981 ( .ip1(n6735), .ip2(n6748), .op(n6736) );
  nand2_1 U8982 ( .ip1(n6737), .ip2(n6736), .op(n6752) );
  inv_1 U8983 ( .ip(n6738), .op(n6739) );
  nand2_1 U8984 ( .ip1(n6744), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[12]), .op(n6747) );
  inv_1 U8985 ( .ip(n6756), .op(n6741) );
  nor2_1 U8986 ( .ip1(n6741), .ip2(n7989), .op(n6742) );
  nand2_1 U8987 ( .ip1(n8741), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[11]), .op(n6745) );
  nor2_1 U8988 ( .ip1(n6744), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[12]), .op(n6827) );
  or2_1 U8989 ( .ip1(n6745), .ip2(n6827), .op(n6746) );
  nand2_1 U8990 ( .ip1(n6747), .ip2(n6746), .op(n6750) );
  nor2_1 U8991 ( .ip1(n8730), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[13]), .op(n6749) );
  and2_1 U8992 ( .ip1(n6750), .ip2(n6828), .op(n6751) );
  nor2_1 U8993 ( .ip1(n6752), .ip2(n6751), .op(n6753) );
  or2_1 U8994 ( .ip1(n6830), .ip2(n6753), .op(n6754) );
  nand2_1 U8995 ( .ip1(n6755), .ip2(n6754), .op(n6835) );
  nand2_1 U8996 ( .ip1(n6764), .ip2(n6756), .op(n6757) );
  nand2_1 U8997 ( .ip1(n6760), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[10]), .op(n6763) );
  inv_1 U8998 ( .ip(n7979), .op(n6758) );
  nand2_1 U8999 ( .ip1(n6764), .ip2(n6758), .op(n6759) );
  inv_1 U9000 ( .ip(n9013), .op(n6772) );
  nand2_1 U9001 ( .ip1(n6772), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[9]), .op(n6761) );
  nor2_1 U9002 ( .ip1(n6760), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[10]), .op(n6773) );
  or2_1 U9003 ( .ip1(n6761), .ip2(n6773), .op(n6762) );
  nand2_1 U9004 ( .ip1(n6763), .ip2(n6762), .op(n6777) );
  nand2_1 U9005 ( .ip1(n5272), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[8]), .op(n6771) );
  inv_1 U9006 ( .ip(n6782), .op(n6765) );
  nor2_1 U9007 ( .ip1(n6765), .ip2(n7965), .op(n6767) );
  inv_1 U9008 ( .ip(n6766), .op(n6790) );
  nand2_1 U9009 ( .ip1(n6767), .ip2(n6790), .op(n6768) );
  nand2_1 U9010 ( .ip1(n8762), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[7]), .op(n6769) );
  nor2_1 U9011 ( .ip1(n5272), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[8]), 
        .op(n6779) );
  or2_1 U9012 ( .ip1(n6769), .ip2(n6779), .op(n6770) );
  nand2_1 U9013 ( .ip1(n6771), .ip2(n6770), .op(n6775) );
  nor2_1 U9014 ( .ip1(n6772), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[9]), 
        .op(n6774) );
  nor2_1 U9015 ( .ip1(n6774), .ip2(n6773), .op(n6780) );
  and2_1 U9016 ( .ip1(n6775), .ip2(n6780), .op(n6776) );
  nor2_1 U9017 ( .ip1(n6777), .ip2(n6776), .op(n6825) );
  nor2_1 U9018 ( .ip1(n8762), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[7]), 
        .op(n6778) );
  nor2_1 U9019 ( .ip1(n6779), .ip2(n6778), .op(n6781) );
  nand2_1 U9020 ( .ip1(n6781), .ip2(n6780), .op(n6823) );
  nand2_1 U9021 ( .ip1(n6790), .ip2(n6782), .op(n6783) );
  inv_1 U9022 ( .ip(n8977), .op(n6784) );
  and2_1 U9023 ( .ip1(n6784), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[6]), 
        .op(n6789) );
  nor2_1 U9024 ( .ip1(n6784), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[6]), 
        .op(n6792) );
  inv_1 U9025 ( .ip(n7958), .op(n6785) );
  nand2_1 U9026 ( .ip1(n6790), .ip2(n6785), .op(n6786) );
  inv_1 U9027 ( .ip(n8980), .op(n6791) );
  nand2_1 U9028 ( .ip1(n6791), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[5]), .op(n6787) );
  nor2_1 U9029 ( .ip1(n6792), .ip2(n6787), .op(n6788) );
  xor2_1 U9030 ( .ip1(n6790), .ip2(n7958), .op(n9001) );
  inv_1 U9031 ( .ip(n9001), .op(n6815) );
  nand2_1 U9032 ( .ip1(n6815), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[4]), .op(n6795) );
  or2_1 U9033 ( .ip1(n6791), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[5]), 
        .op(n6794) );
  inv_1 U9034 ( .ip(n6792), .op(n6793) );
  or2_1 U9035 ( .ip1(n6795), .ip2(n6817), .op(n6796) );
  inv_1 U9036 ( .ip(n6798), .op(n6801) );
  nor2_1 U9037 ( .ip1(n6801), .ip2(n7949), .op(n6799) );
  xor2_1 U9038 ( .ip1(n6799), .ip2(n7941), .op(n6800) );
  nand2_1 U9039 ( .ip1(n5262), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[3]), .op(n6814) );
  nand2_1 U9040 ( .ip1(n8781), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[2]), .op(n6810) );
  nor2_1 U9041 ( .ip1(n8781), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[2]), 
        .op(n6808) );
  and2_1 U9042 ( .ip1(n6802), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[1]), 
        .op(n6806) );
  nor2_1 U9043 ( .ip1(n6802), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[1]), 
        .op(n6804) );
  nor2_1 U9044 ( .ip1(n7943), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[0]), 
        .op(n6803) );
  or2_1 U9045 ( .ip1(n5262), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[3]), 
        .op(n6811) );
  nor2_1 U9046 ( .ip1(n6815), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[4]), 
        .op(n6816) );
  or2_1 U9047 ( .ip1(n6823), .ip2(n6822), .op(n6824) );
  nand2_1 U9048 ( .ip1(n6825), .ip2(n6824), .op(n6833) );
  nor2_1 U9049 ( .ip1(n8741), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[11]), .op(n6826) );
  nor2_1 U9050 ( .ip1(n6827), .ip2(n6826), .op(n6829) );
  nand2_1 U9051 ( .ip1(n6829), .ip2(n6828), .op(n6831) );
  nor2_1 U9052 ( .ip1(n6831), .ip2(n6830), .op(n6832) );
  and2_1 U9053 ( .ip1(n6833), .ip2(n6832), .op(n6834) );
  nor2_2 U9054 ( .ip1(n6835), .ip2(n6834), .op(n8387) );
  inv_1 U9055 ( .ip(n8387), .op(n10589) );
  or2_1 U9056 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl_lcnt_en), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_stop_scl_lcnt_en), .op(n9993) );
  nor3_1 U9057 ( .ip1(i_i2c_rx_scl_lcnt_en), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_data_scl_lcnt_en), .ip3(n9993), .op(n6836)
         );
  or2_1 U9058 ( .ip1(n6836), .ip2(n11152), .op(n10630) );
  and2_1 U9059 ( .ip1(n6838), .ip2(i_i2c_fifo_rst_n), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N48) );
  and2_1 U9060 ( .ip1(n6839), .ip2(i_i2c_fifo_rst_n), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N37) );
  inv_1 U9061 ( .ip(n6939), .op(n8215) );
  nand3_1 U9062 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_addr_2byte_sent), .ip2(n8215), 
        .ip3(i_i2c_U_DW_apb_i2c_mstfsm_N487), .op(n6840) );
  nor2_1 U9063 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv), .ip2(
        i_i2c_hs_mcode_en), .op(n8801) );
  inv_1 U9064 ( .ip(i_i2c_ic_enable_sync), .op(n10915) );
  nor3_1 U9065 ( .ip1(n11170), .ip2(n10915), .ip3(n7080), .op(
        i_i2c_U_DW_apb_i2c_toggle_N33) );
  nor3_1 U9066 ( .ip1(i_i2c_slv_tx_cmplt), .ip2(n6841), .ip3(n11293), .op(
        n5109) );
  inv_1 U9067 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[3]), .op(
        n11175) );
  nand2_1 U9068 ( .ip1(i_i2c_slv_tx_ready_unconn), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly1), .op(n6842) );
  or3_1 U9069 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[1]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[0]), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[2]), .op(n7719) );
  and3_1 U9070 ( .ip1(n11769), .ip2(n5109), .ip3(n7713), .op(n5112) );
  or2_1 U9071 ( .ip1(i_i2c_byte_wait_scl), .ip2(n6847), .op(n7069) );
  inv_1 U9072 ( .ip(i_i2c_tx_fifo_rst_n), .op(n11258) );
  inv_1 U9073 ( .ip(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[2]), .op(n6854) );
  inv_1 U9074 ( .ip(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[0]), .op(n6858) );
  inv_1 U9075 ( .ip(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_empty_n), .op(n5246) );
  xor2_1 U9076 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_tx_pop_flg_sync), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_pop_flg_sync_q), .op(i_i2c_tx_pop_sync) );
  nor2_1 U9077 ( .ip1(i_i2c_tx_pop_sync), .ip2(i_i2c_tx_full), .op(n6849) );
  nor2_1 U9078 ( .ip1(n5246), .ip2(n6849), .op(n6850) );
  inv_1 U9079 ( .ip(i_i2c_tx_push), .op(n6965) );
  nor2_1 U9080 ( .ip1(n5246), .ip2(n11261), .op(n11259) );
  inv_1 U9081 ( .ip(n11259), .op(n8213) );
  nor2_1 U9082 ( .ip1(i_i2c_tx_push), .ip2(n8213), .op(n6859) );
  nor2_1 U9083 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[0]), .ip2(n6863), 
        .op(n6864) );
  nor2_1 U9084 ( .ip1(n6860), .ip2(n6864), .op(n6852) );
  nor2_1 U9085 ( .ip1(n6859), .ip2(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[1]), 
        .op(n6851) );
  not_ab_or_c_or_d U9086 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[1]), 
        .ip2(n6858), .ip3(n6852), .ip4(n6851), .op(n6853) );
  nand2_1 U9087 ( .ip1(i_i2c_tx_push), .ip2(i_i2c_tx_full), .op(n11260) );
  nand2_1 U9088 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[0]), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[1]), .op(n6855) );
  nor3_1 U9089 ( .ip1(n6855), .ip2(n6965), .ip3(n6854), .op(n6856) );
  nor2_1 U9090 ( .ip1(i_i2c_tx_full), .ip2(n6856), .op(n6857) );
  not_ab_or_c_or_d U9091 ( .ip1(i_i2c_tx_pop_sync), .ip2(n11260), .ip3(n6857), 
        .ip4(n11258), .op(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N37) );
  inv_1 U9092 ( .ip(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[1]), .op(n6862) );
  mux2_1 U9093 ( .ip1(n6860), .ip2(n6859), .s(n6858), .op(n6861) );
  nor2_1 U9094 ( .ip1(n11258), .ip2(n7055), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N48) );
  or2_1 U9095 ( .ip1(n6863), .ip2(n6864), .op(n6866) );
  or2_1 U9096 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[0]), .ip2(n6864), 
        .op(n6865) );
  nand2_1 U9097 ( .ip1(n6866), .ip2(n6865), .op(n7054) );
  nor2_1 U9098 ( .ip1(n7054), .ip2(n11258), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N47) );
  or4_1 U9099 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N49), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N37), .ip3(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N48), .ip4(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N47), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N33) );
  nand3_1 U9100 ( .ip1(n6869), .ip2(n6868), .ip3(n6867), .op(n6872) );
  nand2_1 U9101 ( .ip1(n6870), .ip2(n6905), .op(n6871) );
  nand4_1 U9102 ( .ip1(n10413), .ip2(n8217), .ip3(n6872), .ip4(n6871), .op(
        n11306) );
  and3_1 U9103 ( .ip1(n6470), .ip2(n7361), .ip3(n11306), .op(n6960) );
  nand2_1 U9104 ( .ip1(i_i2c_scl_s_hld_cmplt), .ip2(n6954), .op(n6873) );
  inv_1 U9105 ( .ip(n7075), .op(n6875) );
  nand2_1 U9106 ( .ip1(n6875), .ip2(n6874), .op(n6876) );
  inv_1 U9107 ( .ip(i_i2c_start_en), .op(n8442) );
  nor2_1 U9108 ( .ip1(n7075), .ip2(n6877), .op(n6879) );
  inv_1 U9109 ( .ip(n6880), .op(n8428) );
  nor2_1 U9110 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_N252), .ip2(n8428), .op(n6878)
         );
  or2_1 U9111 ( .ip1(n6879), .ip2(n6878), .op(n8340) );
  inv_1 U9112 ( .ip(i_i2c_scl_s_hld_cmplt), .op(n7740) );
  nand2_1 U9113 ( .ip1(n6880), .ip2(n7740), .op(n6886) );
  nand2_1 U9114 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_10bit_mst_sync_inv), .ip2(
        n8418), .op(n6885) );
  nor3_1 U9115 ( .ip1(n6905), .ip2(n7073), .ip3(n6881), .op(n6934) );
  inv_1 U9116 ( .ip(n6941), .op(n6882) );
  nand2_1 U9117 ( .ip1(n6934), .ip2(n6882), .op(n6884) );
  nand4_1 U9118 ( .ip1(n6886), .ip2(n6885), .ip3(n6884), .ip4(n6883), .op(
        n6896) );
  nand2_1 U9119 ( .ip1(n9096), .ip2(n9735), .op(n6893) );
  inv_1 U9120 ( .ip(n6888), .op(n6889) );
  nand2_1 U9121 ( .ip1(n6890), .ip2(n6889), .op(n6891) );
  ab_or_c_or_d U9122 ( .ip1(n6897), .ip2(n8340), .ip3(n6896), .ip4(n6895), 
        .op(n6898) );
  not_ab_or_c_or_d U9123 ( .ip1(n6900), .ip2(n6616), .ip3(n6899), .ip4(n6898), 
        .op(n6924) );
  nor2_1 U9124 ( .ip1(n8339), .ip2(n6901), .op(n6920) );
  inv_1 U9125 ( .ip(n6902), .op(n6904) );
  nand4_1 U9126 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_byte_waiting_q), .ip2(n6905), 
        .ip3(n6904), .ip4(n6903), .op(n6906) );
  nand2_1 U9127 ( .ip1(n6907), .ip2(n6906), .op(n6918) );
  inv_1 U9128 ( .ip(n6908), .op(n6909) );
  nand3_1 U9129 ( .ip1(n6912), .ip2(
        i_i2c_U_DW_apb_i2c_sync_ic_rstrt_en_sync_inv), .ip3(n6911), .op(n6917)
         );
  inv_1 U9130 ( .ip(n6913), .op(n6914) );
  nand3_1 U9131 ( .ip1(n6915), .ip2(n6914), .ip3(n9997), .op(n6916) );
  nand2_1 U9132 ( .ip1(n9740), .ip2(n9667), .op(n6923) );
  nor2_1 U9133 ( .ip1(i_i2c_ic_abort_sync), .ip2(n5245), .op(n6921) );
  nand2_1 U9134 ( .ip1(n8339), .ip2(n6921), .op(n6922) );
  or2_1 U9135 ( .ip1(n6946), .ip2(n6925), .op(n11047) );
  nand2_1 U9136 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_rstrt_en_sync_inv), .ip2(
        n6927), .op(n6930) );
  not_ab_or_c_or_d U9137 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_addr_1byte_sent), 
        .ip2(n6930), .ip3(n6929), .ip4(n6928), .op(n6933) );
  inv_1 U9138 ( .ip(n6931), .op(n6932) );
  inv_1 U9139 ( .ip(n6934), .op(n6935) );
  nand2_1 U9140 ( .ip1(n6936), .ip2(n6935), .op(n6940) );
  nor3_1 U9141 ( .ip1(n6937), .ip2(n8428), .ip3(n7740), .op(n6938) );
  not_ab_or_c_or_d U9142 ( .ip1(n6941), .ip2(n6940), .ip3(n6939), .ip4(n6938), 
        .op(n6942) );
  nand2_1 U9143 ( .ip1(n9448), .ip2(i_i2c_tx_fifo_data_buf[8]), .op(n8333) );
  not_ab_or_c_or_d U9144 ( .ip1(n9723), .ip2(n9699), .ip3(n9153), .ip4(n6944), 
        .op(n6950) );
  or2_1 U9145 ( .ip1(n8266), .ip2(n6945), .op(n6949) );
  inv_1 U9146 ( .ip(n6946), .op(n6947) );
  inv_1 U9147 ( .ip(n9661), .op(n6948) );
  not_ab_or_c_or_d U9148 ( .ip1(i_i2c_ic_bus_idle), .ip2(n5232), .ip3(
        i_i2c_start_en), .ip4(n6953), .op(n6956) );
  xor2_1 U9149 ( .ip1(i_i2c_U_DW_apb_i2c_intctl_set_tx_empty_en_flg_sync_q), 
        .ip2(i_i2c_U_DW_apb_i2c_intctl_set_tx_empty_en_flg_sync), .op(n6963)
         );
  and2_1 U9150 ( .ip1(i_i2c_tx_fifo_rst_n), .ip2(n6963), .op(n9927) );
  nand2_1 U9151 ( .ip1(n6962), .ip2(n9930), .op(n6967) );
  inv_1 U9152 ( .ip(n6963), .op(n6964) );
  and3_1 U9153 ( .ip1(i_i2c_tx_fifo_rst_n), .ip2(n6965), .ip3(n6964), .op(
        n9932) );
  nand2_1 U9154 ( .ip1(n9932), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[6]), .op(n6966) );
  nand2_1 U9155 ( .ip1(n6967), .ip2(n6966), .op(n4136) );
  or2_1 U9156 ( .ip1(n9935), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[0]), 
        .op(n6968) );
  nand2_1 U9157 ( .ip1(n6969), .ip2(n6968), .op(n6970) );
  nor2_1 U9158 ( .ip1(n6971), .ip2(n9692), .op(n6975) );
  nor2_1 U9159 ( .ip1(i_ssi_tx_rd_addr[0]), .ip2(n6972), .op(n6974) );
  nand2_1 U9160 ( .ip1(n6972), .ip2(i_ssi_U_fifo_U_tx_fifo_rd_addr_at_max), 
        .op(n6973) );
  nand2_1 U9161 ( .ip1(n6973), .ip2(n11219), .op(n8576) );
  nor3_1 U9162 ( .ip1(n6975), .ip2(n6974), .ip3(n8576), .op(n11767) );
  nor2_1 U9163 ( .ip1(i_ssi_tx_rd_addr[1]), .ip2(n6975), .op(n6977) );
  nand2_1 U9164 ( .ip1(n6975), .ip2(i_ssi_tx_rd_addr[1]), .op(n8574) );
  inv_1 U9165 ( .ip(n8574), .op(n6976) );
  nor2_1 U9166 ( .ip1(n6978), .ip2(n5571), .op(n6979) );
  inv_1 U9167 ( .ip(n6980), .op(n6984) );
  nor2_1 U9168 ( .ip1(i_ssi_U_mstfsm_c_state[2]), .ip2(n9058), .op(n6981) );
  nand2_1 U9169 ( .ip1(n8381), .ip2(n6981), .op(n6983) );
  nand2_1 U9170 ( .ip1(n9684), .ip2(i_ssi_sclk_fe), .op(n6982) );
  inv_1 U9171 ( .ip(n10480), .op(n6986) );
  nand2_1 U9172 ( .ip1(n6986), .ip2(i_ssi_U_mstfsm_spi1_control), .op(n6987)
         );
  inv_1 U9173 ( .ip(i_i2c_fifo_rst_n), .op(n11207) );
  or4_1 U9174 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N47), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N37), .ip3(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N48), .ip4(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N49), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N33) );
  and3_1 U9175 ( .ip1(i_ssi_U_fifo_unconnected_tx_wrd_count[2]), .ip2(
        i_ssi_U_fifo_unconnected_tx_wrd_count[1]), .ip3(
        i_ssi_U_fifo_unconnected_tx_wrd_count[0]), .op(n6990) );
  nand2_1 U9176 ( .ip1(n6991), .ip2(n6990), .op(n6993) );
  nand2_1 U9177 ( .ip1(n9071), .ip2(i_ssi_tx_full), .op(n6992) );
  and2_1 U9178 ( .ip1(n6994), .ip2(n11219), .op(i_ssi_U_fifo_U_tx_fifo_N37) );
  nand3_1 U9179 ( .ip1(n7634), .ip2(n6470), .ip3(n7361), .op(
        i_i2c_U_DW_apb_i2c_toggle_N31) );
  nor3_1 U9180 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(i_i2c_byte_wait_scl), .ip3(
        n7361), .op(n11773) );
  inv_1 U9181 ( .ip(i_i2c_rx_scl_lcnt_en), .op(n6995) );
  inv_1 U9182 ( .ip(i_i2c_rx_scl_hcnt_en), .op(n10572) );
  inv_1 U9183 ( .ip(i_i2c_mst_rx_bit_count[3]), .op(n10569) );
  nor4_1 U9184 ( .ip1(i_i2c_mst_rx_bit_count[2]), .ip2(
        i_i2c_mst_rx_bit_count[0]), .ip3(i_i2c_mst_rx_bit_count[1]), .ip4(
        n10569), .op(n7690) );
  nand3_1 U9185 ( .ip1(n7689), .ip2(n7690), .ip3(n11152), .op(n6997) );
  nor2_1 U9186 ( .ip1(n10566), .ip2(n6997), .op(n4938) );
  inv_1 U9187 ( .ip(n11152), .op(n7420) );
  inv_1 U9188 ( .ip(i_i2c_mst_rx_bit_count[0]), .op(n8318) );
  nand2_1 U9189 ( .ip1(i_i2c_mst_rx_bit_count[0]), .ip2(n8322), .op(n6998) );
  nand2_1 U9190 ( .ip1(n9645), .ip2(n6998), .op(n5116) );
  inv_1 U9191 ( .ip(i_i2c_mst_rx_bit_count[1]), .op(n9642) );
  nand4_1 U9192 ( .ip1(i_i2c_mst_rx_bit_count[0]), .ip2(n11773), .ip3(n9612), 
        .ip4(n9642), .op(n9632) );
  inv_1 U9193 ( .ip(n8322), .op(n6999) );
  nand2_1 U9194 ( .ip1(i_i2c_mst_rx_bit_count[1]), .ip2(n11311), .op(n7000) );
  nand2_1 U9195 ( .ip1(n9632), .ip2(n7000), .op(n5115) );
  inv_1 U9196 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[5]), .op(
        n11146) );
  or2_1 U9197 ( .ip1(i_i2c_ic_sda_rx_hold_sync[4]), .ip2(n7001), .op(n7004) );
  or2_1 U9198 ( .ip1(n7002), .ip2(n7001), .op(n7003) );
  nand2_1 U9199 ( .ip1(n7004), .ip2(n7003), .op(n7015) );
  nor2_1 U9200 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[4]), 
        .ip2(n7015), .op(n7007) );
  or2_1 U9201 ( .ip1(n11146), .ip2(n7007), .op(n7009) );
  nand2_1 U9202 ( .ip1(i_i2c_ic_sda_rx_hold_sync[5]), .ip2(n7005), .op(n7006)
         );
  nand2_1 U9203 ( .ip1(n7032), .ip2(n7006), .op(n7030) );
  or2_1 U9204 ( .ip1(n7030), .ip2(n7007), .op(n7008) );
  nand2_1 U9205 ( .ip1(n7009), .ip2(n7008), .op(n7038) );
  or2_1 U9206 ( .ip1(i_i2c_ic_sda_rx_hold_sync[3]), .ip2(n7011), .op(n7014) );
  inv_1 U9207 ( .ip(i_i2c_ic_sda_rx_hold_sync[2]), .op(n7010) );
  nor2_1 U9208 ( .ip1(i_i2c_ic_sda_rx_hold_sync[1]), .ip2(
        i_i2c_ic_sda_rx_hold_sync[0]), .op(n7020) );
  nand2_1 U9209 ( .ip1(n7010), .ip2(n7020), .op(n7012) );
  or2_1 U9210 ( .ip1(n7012), .ip2(n7011), .op(n7013) );
  nand2_1 U9211 ( .ip1(n7014), .ip2(n7013), .op(n7027) );
  nand2_1 U9212 ( .ip1(n7027), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[3]), .op(n7017) );
  nand2_1 U9213 ( .ip1(n7015), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[4]), .op(n7016) );
  nand2_1 U9214 ( .ip1(n7017), .ip2(n7016), .op(n9755) );
  or2_1 U9215 ( .ip1(i_i2c_ic_sda_rx_hold_sync[0]), .ip2(n7020), .op(n7019) );
  or2_1 U9216 ( .ip1(i_i2c_ic_sda_rx_hold_sync[1]), .ip2(n7020), .op(n7018) );
  nand2_1 U9217 ( .ip1(n7019), .ip2(n7018), .op(n7024) );
  inv_1 U9218 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[2]), .op(
        n11139) );
  xor2_1 U9219 ( .ip1(i_i2c_ic_sda_rx_hold_sync[2]), .ip2(n7020), .op(n7028)
         );
  nor2_1 U9220 ( .ip1(n11139), .ip2(n7028), .op(n7021) );
  or2_1 U9221 ( .ip1(n7024), .ip2(n7021), .op(n7023) );
  or2_1 U9222 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[1]), 
        .ip2(n7021), .op(n7022) );
  nand2_1 U9223 ( .ip1(n7023), .ip2(n7022), .op(n9754) );
  nor2_1 U9224 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[1]), 
        .ip2(n7024), .op(n7026) );
  nor2_1 U9225 ( .ip1(i_i2c_ic_sda_rx_hold_sync[0]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[0]), .op(n7025) );
  or2_1 U9226 ( .ip1(n7026), .ip2(n7025), .op(n9760) );
  nor2_1 U9227 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[3]), 
        .ip2(n7027), .op(n9758) );
  nand2_1 U9228 ( .ip1(n11139), .ip2(n7028), .op(n7029) );
  nand2_1 U9229 ( .ip1(n7038), .ip2(n7029), .op(n9750) );
  not_ab_or_c_or_d U9230 ( .ip1(n9754), .ip2(n9760), .ip3(n9758), .ip4(n9750), 
        .op(n7037) );
  or2_1 U9231 ( .ip1(n7030), .ip2(n11146), .op(n7036) );
  or2_1 U9232 ( .ip1(i_i2c_ic_sda_rx_hold_sync[6]), .ip2(n7031), .op(n7034) );
  or2_1 U9233 ( .ip1(n7032), .ip2(n7031), .op(n7033) );
  nand2_1 U9234 ( .ip1(n7039), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[6]), .op(n7035) );
  not_ab_or_c_or_d U9235 ( .ip1(n7038), .ip2(n9755), .ip3(n7037), .ip4(n9751), 
        .op(n7043) );
  nor2_1 U9236 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[6]), 
        .ip2(n7039), .op(n9757) );
  or2_1 U9237 ( .ip1(i_i2c_ic_sda_rx_hold_sync[7]), .ip2(n7046), .op(n7041) );
  or2_1 U9238 ( .ip1(n7044), .ip2(n7046), .op(n7040) );
  nor2_1 U9239 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[7]), 
        .ip2(n7042), .op(n9753) );
  inv_1 U9240 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[7]), .op(
        n7506) );
  not_ab_or_c_or_d U9241 ( .ip1(i_i2c_ic_sda_rx_hold_sync[7]), .ip2(n7044), 
        .ip3(n7046), .ip4(n7506), .op(n9752) );
  nor2_1 U9242 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[0]), 
        .ip2(n7047), .op(n7050) );
  nand2_1 U9243 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[0]), 
        .ip2(n7047), .op(n11133) );
  mux2_1 U9244 ( .ip1(n9765), .ip2(n7048), .s(
        i_i2c_U_DW_apb_i2c_rx_filter_sda_post_hold_done), .op(n7049) );
  nand2_1 U9245 ( .ip1(n11776), .ip2(n7049), .op(n11144) );
  nor2_1 U9246 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[17]), .ip2(n7051), 
        .op(ex_i_ahb_AHB_Slave_RAM_hsel) );
  inv_1 U9247 ( .ip(ex_i_ahb_AHB_Slave_RAM_hsel), .op(n7052) );
  nand4_1 U9248 ( .ip1(n11355), .ip2(n9070), .ip3(n7052), .ip4(
        ex_i_ahb_AHB_MASTER_CORTEXM0_htrans[1]), .op(n11182) );
  inv_1 U9249 ( .ip(i_i2c_ic_tx_tl[2]), .op(n8461) );
  not_ab_or_c_or_d U9250 ( .ip1(i_i2c_tx_fifo_rst_n), .ip2(n8461), .ip3(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N37), .ip4(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N49), .op(n7061) );
  nor2_1 U9251 ( .ip1(n7053), .ip2(i_i2c_ic_tx_tl[2]), .op(n7059) );
  nor2_1 U9252 ( .ip1(n7055), .ip2(i_i2c_ic_tx_tl[1]), .op(n7057) );
  not_ab_or_c_or_d U9253 ( .ip1(i_i2c_ic_tx_tl[1]), .ip2(n7055), .ip3(n7054), 
        .ip4(i_i2c_ic_tx_tl[0]), .op(n7056) );
  or2_1 U9254 ( .ip1(n7057), .ip2(n7056), .op(n7058) );
  nor2_1 U9255 ( .ip1(n7061), .ip2(n7060), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N34) );
  fulladder U9256 ( .a(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[5]), .b(n9927), 
        .ci(n7062), .co(n9926), .s(n7063) );
  nand2_1 U9257 ( .ip1(n7063), .ip2(n9930), .op(n7065) );
  nand2_1 U9258 ( .ip1(n9932), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[5]), .op(n7064) );
  nand2_1 U9259 ( .ip1(n7065), .ip2(n7064), .op(n4137) );
  nor4_1 U9260 ( .ip1(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[0]), 
        .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[3]), 
        .ip3(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[2]), 
        .ip4(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[1]), 
        .op(n7066) );
  nand2_1 U9261 ( .ip1(n7066), .ip2(n8534), .op(n7077) );
  inv_1 U9262 ( .ip(i_i2c_ic_data_oe), .op(n7067) );
  xor2_1 U9263 ( .ip1(n7067), .ip2(n10579), .op(n7068) );
  nand2_1 U9264 ( .ip1(i_i2c_mst_rx_ack_vld), .ip2(n11773), .op(n7688) );
  nand2_1 U9265 ( .ip1(n7069), .ip2(n7688), .op(n7071) );
  nand2_1 U9266 ( .ip1(i_i2c_mst_tx_ack_vld), .ip2(n7688), .op(n7070) );
  nand3_1 U9267 ( .ip1(n8569), .ip2(n7071), .ip3(n7070), .op(n7076) );
  or3_1 U9268 ( .ip1(i_i2c_mst_debug_cstate[3]), .ip2(
        i_i2c_U_DW_apb_i2c_mstfsm_delay_stop_en), .ip3(n7072), .op(n7074) );
  not_ab_or_c_or_d U9269 ( .ip1(n7075), .ip2(n7074), .ip3(i_i2c_byte_wait_scl), 
        .ip4(n7073), .op(n11774) );
  not_ab_or_c_or_d U9270 ( .ip1(n7077), .ip2(n7076), .ip3(n11774), .ip4(
        i_i2c_start_en), .op(n7079) );
  and2_1 U9271 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_mst_arb_lost), .ip2(n11167), 
        .op(n7078) );
  inv_1 U9272 ( .ip(i_ssi_tx_pop_sync), .op(n7084) );
  inv_1 U9273 ( .ip(i_ssi_U_regfile_txflr[3]), .op(n11518) );
  nand2_1 U9274 ( .ip1(n11569), .ip2(n11518), .op(n7082) );
  nor2_1 U9275 ( .ip1(n7082), .ip2(n7087), .op(n7083) );
  nor2_1 U9276 ( .ip1(i_ssi_U_regfile_txflr[1]), .ip2(n9973), .op(n9971) );
  nand2_1 U9277 ( .ip1(i_ssi_U_regfile_txflr[0]), .ip2(n9971), .op(n7092) );
  nor4_1 U9278 ( .ip1(i_ssi_U_regfile_txflr[0]), .ip2(i_ssi_U_regfile_txflr[1]), .ip3(i_ssi_U_regfile_txflr[2]), .ip4(i_ssi_U_regfile_txflr[3]), .op(n7085)
         );
  nor2_1 U9279 ( .ip1(n7085), .ip2(n11148), .op(n7086) );
  and2_1 U9280 ( .ip1(n7087), .ip2(n7086), .op(n7088) );
  nand2_1 U9281 ( .ip1(i_ssi_tx_pop_sync), .ip2(n7088), .op(n9969) );
  nor2_1 U9282 ( .ip1(i_ssi_U_regfile_txflr[0]), .ip2(i_ssi_U_regfile_txflr[1]), .op(n7089) );
  nand3_1 U9283 ( .ip1(n9973), .ip2(n11569), .ip3(n9969), .op(n9946) );
  inv_1 U9284 ( .ip(i_ssi_U_regfile_txflr[0]), .op(n11581) );
  nand2_1 U9285 ( .ip1(i_ssi_U_regfile_txflr[1]), .ip2(n9970), .op(n7091) );
  inv_1 U9286 ( .ip(i_i2c_ic_clk_oe), .op(n10005) );
  or2_1 U9287 ( .ip1(n7185), .ip2(n9773), .op(n7098) );
  or2_1 U9288 ( .ip1(i_i2c_ic_sda_tx_hold_sync[7]), .ip2(n7098), .op(n7101) );
  nand2_1 U9289 ( .ip1(n7101), .ip2(i_i2c_ic_sda_tx_hold_sync[8]), .op(n7250)
         );
  inv_1 U9290 ( .ip(i_i2c_ic_sda_tx_hold_sync[10]), .op(n7094) );
  inv_1 U9291 ( .ip(i_i2c_ic_sda_tx_hold_sync[9]), .op(n7093) );
  nor2_1 U9292 ( .ip1(n7211), .ip2(i_i2c_ic_sda_tx_hold_sync[13]), .op(n7204)
         );
  inv_1 U9293 ( .ip(i_i2c_ic_sda_tx_hold_sync[14]), .op(n7096) );
  or2_1 U9294 ( .ip1(n7180), .ip2(n9773), .op(n7106) );
  or2_1 U9295 ( .ip1(i_i2c_ic_sda_tx_hold_sync[6]), .ip2(n7106), .op(n7103) );
  nor2_1 U9296 ( .ip1(n7101), .ip2(i_i2c_ic_sda_tx_hold_sync[8]), .op(n7105)
         );
  or2_1 U9297 ( .ip1(n7150), .ip2(n9773), .op(n7107) );
  inv_1 U9298 ( .ip(n7164), .op(n7146) );
  or2_1 U9299 ( .ip1(n7146), .ip2(n9773), .op(n7115) );
  or2_1 U9300 ( .ip1(i_i2c_ic_sda_tx_hold_sync[4]), .ip2(n7115), .op(n7112) );
  inv_1 U9301 ( .ip(n7145), .op(n7152) );
  or2_1 U9302 ( .ip1(n7152), .ip2(n9773), .op(n7116) );
  or2_1 U9303 ( .ip1(i_i2c_ic_sda_tx_hold_sync[3]), .ip2(n7116), .op(n7119) );
  or2_1 U9304 ( .ip1(n7160), .ip2(n9773), .op(n7122) );
  or2_1 U9305 ( .ip1(i_i2c_ic_sda_tx_hold_sync[2]), .ip2(n7122), .op(n7136) );
  nand2_1 U9306 ( .ip1(n7123), .ip2(n9773), .op(n7306) );
  nand2_1 U9307 ( .ip1(n7156), .ip2(i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv), .op(n7130) );
  nand2_1 U9308 ( .ip1(i_i2c_ic_sda_tx_hold_sync[0]), .ip2(
        i_i2c_ic_sda_tx_hold_sync[1]), .op(n7125) );
  and2_1 U9309 ( .ip1(n7200), .ip2(n7128), .op(n7827) );
  inv_1 U9310 ( .ip(n7827), .op(n7911) );
  nand2_1 U9311 ( .ip1(n9773), .ip2(n7911), .op(n7129) );
  nand2_1 U9312 ( .ip1(n7130), .ip2(n7129), .op(n7132) );
  inv_1 U9313 ( .ip(n7132), .op(n7131) );
  inv_1 U9314 ( .ip(i_i2c_ic_sda_tx_hold_sync[1]), .op(n7155) );
  and2_1 U9315 ( .ip1(n7132), .ip2(n7155), .op(n7313) );
  nand2_1 U9316 ( .ip1(n7154), .ip2(i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv), .op(n7320) );
  nor2_1 U9317 ( .ip1(i_i2c_ic_sda_tx_hold_sync[0]), .ip2(n7320), .op(n7316)
         );
  or2_1 U9318 ( .ip1(n7305), .ip2(n7308), .op(n7135) );
  and2_1 U9319 ( .ip1(n7299), .ip2(n7138), .op(n7139) );
  nand2_1 U9320 ( .ip1(n7142), .ip2(n7245), .op(n7143) );
  inv_1 U9321 ( .ip(i_i2c_ic_sda_tx_hold_sync[8]), .op(n7194) );
  nor2_1 U9322 ( .ip1(n7146), .ip2(n7163), .op(n7148) );
  nand2_1 U9323 ( .ip1(n7147), .ip2(n7148), .op(n7181) );
  inv_1 U9324 ( .ip(n7148), .op(n7149) );
  nand2_1 U9325 ( .ip1(n7150), .ip2(n7149), .op(n7151) );
  nand2_1 U9326 ( .ip1(n7181), .ip2(n7151), .op(n7175) );
  nand2_1 U9327 ( .ip1(n7152), .ip2(n7160), .op(n7153) );
  nand2_1 U9328 ( .ip1(n7163), .ip2(n7153), .op(n7162) );
  nand2_1 U9329 ( .ip1(i_i2c_ic_sda_tx_hold_sync[3]), .ip2(n7162), .op(n7168)
         );
  inv_1 U9330 ( .ip(i_i2c_ic_sda_tx_hold_sync[0]), .op(n7912) );
  not_ab_or_c_or_d U9331 ( .ip1(n7156), .ip2(n7155), .ip3(n7154), .ip4(n7912), 
        .op(n7158) );
  nor2_1 U9332 ( .ip1(n7156), .ip2(n7155), .op(n7157) );
  fulladder U9333 ( .a(n7159), .b(n7161), .ci(n7160), .co(n7167) );
  nor2_1 U9334 ( .ip1(i_i2c_ic_sda_tx_hold_sync[3]), .ip2(n7162), .op(n7166)
         );
  xor2_1 U9335 ( .ip1(n7164), .ip2(n7163), .op(n7169) );
  nor2_4 U9336 ( .ip1(i_i2c_ic_sda_tx_hold_sync[4]), .ip2(n7169), .op(n7165)
         );
  not_ab_or_c_or_d U9337 ( .ip1(n7168), .ip2(n7167), .ip3(n7166), .ip4(n7165), 
        .op(n7173) );
  inv_1 U9338 ( .ip(i_i2c_ic_sda_tx_hold_sync[4]), .op(n7170) );
  or2_1 U9339 ( .ip1(n7173), .ip2(n7172), .op(n7174) );
  fulladder U9340 ( .a(i_i2c_ic_sda_tx_hold_sync[5]), .b(n7175), .ci(n7174), 
        .co(n7187) );
  and2_1 U9341 ( .ip1(n7187), .ip2(i_i2c_ic_sda_tx_hold_sync[6]), .op(n7179)
         );
  inv_1 U9342 ( .ip(n7181), .op(n7177) );
  not_ab_or_c_or_d U9343 ( .ip1(i_i2c_ic_sda_tx_hold_sync[7]), .ip2(n7185), 
        .ip3(n7179), .ip4(n7178), .op(n7192) );
  nor2_1 U9344 ( .ip1(n7181), .ip2(n7180), .op(n7183) );
  nand2_1 U9345 ( .ip1(n7182), .ip2(n7183), .op(n7186) );
  inv_1 U9346 ( .ip(n7186), .op(n7196) );
  inv_1 U9347 ( .ip(n7183), .op(n7184) );
  nand2_1 U9348 ( .ip1(n7186), .ip2(n7189), .op(n7188) );
  not_ab_or_c_or_d U9349 ( .ip1(i_i2c_ic_sda_tx_hold_sync[7]), .ip2(n7188), 
        .ip3(i_i2c_ic_sda_tx_hold_sync[6]), .ip4(n7187), .op(n7195) );
  inv_1 U9350 ( .ip(n7189), .op(n7190) );
  nor2_1 U9351 ( .ip1(i_i2c_ic_sda_tx_hold_sync[7]), .ip2(n7190), .op(n7191)
         );
  or4_1 U9352 ( .ip1(n7192), .ip2(n7196), .ip3(n7195), .ip4(n7191), .op(n7193)
         );
  nand2_1 U9353 ( .ip1(n7194), .ip2(n7193), .op(n7198) );
  nand2_1 U9354 ( .ip1(n7196), .ip2(n7195), .op(n7197) );
  nand2_1 U9355 ( .ip1(n7198), .ip2(n7197), .op(n7199) );
  nor2_4 U9356 ( .ip1(n9773), .ip2(n7201), .op(n7321) );
  and2_1 U9357 ( .ip1(n7202), .ip2(n7248), .op(n7863) );
  inv_1 U9358 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[15]), .op(
        n7862) );
  inv_1 U9359 ( .ip(n7863), .op(n7203) );
  inv_1 U9360 ( .ip(n7204), .op(n7205) );
  nand2_1 U9361 ( .ip1(n7208), .ip2(n7245), .op(n7209) );
  and2_1 U9362 ( .ip1(n7210), .ip2(n7248), .op(n7354) );
  inv_1 U9363 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[14]), .op(
        n11102) );
  nand2_1 U9364 ( .ip1(n7214), .ip2(n7245), .op(n7215) );
  and2_1 U9365 ( .ip1(n7216), .ip2(n7248), .op(n7871) );
  inv_1 U9366 ( .ip(n7871), .op(n7353) );
  nand2_1 U9367 ( .ip1(n7221), .ip2(n7245), .op(n7222) );
  and2_1 U9368 ( .ip1(n7223), .ip2(n7248), .op(n7887) );
  inv_1 U9369 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[12]), .op(
        n11094) );
  nand2_1 U9370 ( .ip1(n7227), .ip2(n7245), .op(n7228) );
  and2_1 U9371 ( .ip1(n7229), .ip2(n7248), .op(n7858) );
  inv_1 U9372 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[11]), .op(
        n11092) );
  nand2_1 U9373 ( .ip1(n7858), .ip2(n11092), .op(n7889) );
  inv_1 U9374 ( .ip(n7889), .op(n7237) );
  nor2_1 U9375 ( .ip1(n7230), .ip2(i_i2c_ic_sda_tx_hold_sync[9]), .op(n7231)
         );
  nand2_1 U9376 ( .ip1(n7233), .ip2(n7245), .op(n7234) );
  and2_1 U9377 ( .ip1(n7235), .ip2(n7248), .op(n7892) );
  inv_1 U9378 ( .ip(n7892), .op(n7239) );
  nor2_1 U9379 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[10]), .ip2(
        n7239), .op(n7236) );
  nor2_1 U9380 ( .ip1(n7237), .ip2(n7236), .op(n7242) );
  inv_1 U9381 ( .ip(n7858), .op(n7238) );
  nand2_1 U9382 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[11]), 
        .ip2(n7238), .op(n7241) );
  nand3_1 U9383 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[10]), 
        .ip2(n7889), .ip3(n7239), .op(n7240) );
  nand2_1 U9384 ( .ip1(n7241), .ip2(n7240), .op(n7347) );
  nor2_1 U9385 ( .ip1(n7242), .ip2(n7347), .op(n7351) );
  nand2_1 U9386 ( .ip1(n7246), .ip2(n7245), .op(n7247) );
  and2_1 U9387 ( .ip1(n7249), .ip2(n7248), .op(n7893) );
  inv_1 U9388 ( .ip(n7893), .op(n7349) );
  inv_1 U9389 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[9]), .op(
        n11086) );
  or2_1 U9390 ( .ip1(n7256), .ip2(n7284), .op(n7257) );
  inv_1 U9391 ( .ip(n7880), .op(n7262) );
  nor2_1 U9392 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[8]), .ip2(
        n7262), .op(n7346) );
  inv_1 U9393 ( .ip(n7284), .op(n7275) );
  nand2_1 U9394 ( .ip1(n7275), .ip2(n7265), .op(n7266) );
  nand2_1 U9395 ( .ip1(n7267), .ip2(n7266), .op(n7268) );
  inv_1 U9396 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[7]), .op(
        n11080) );
  nand2_1 U9397 ( .ip1(n7343), .ip2(n11080), .op(n7882) );
  nand2_1 U9398 ( .ip1(n7275), .ip2(n7282), .op(n7276) );
  nand2_1 U9399 ( .ip1(n7281), .ip2(n7276), .op(n7277) );
  inv_1 U9400 ( .ip(n7828), .op(n7280) );
  nand2_1 U9401 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[6]), .ip2(
        n7280), .op(n7342) );
  inv_1 U9402 ( .ip(n7830), .op(n7287) );
  nand2_1 U9403 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[5]), .ip2(
        n7287), .op(n7339) );
  inv_1 U9404 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[5]), .op(
        n11074) );
  nand2_1 U9405 ( .ip1(n7830), .ip2(n11074), .op(n7829) );
  inv_1 U9406 ( .ip(n7288), .op(n7290) );
  inv_1 U9407 ( .ip(n7291), .op(n7298) );
  nand2_1 U9408 ( .ip1(n7299), .ip2(n7298), .op(n7292) );
  inv_1 U9409 ( .ip(n7837), .op(n7296) );
  nand2_1 U9410 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[4]), .ip2(
        n7296), .op(n7336) );
  inv_1 U9411 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[4]), .op(
        n11070) );
  nand2_1 U9412 ( .ip1(n7837), .ip2(n11070), .op(n7848) );
  nand2_1 U9413 ( .ip1(n7298), .ip2(n7297), .op(n7301) );
  inv_1 U9414 ( .ip(n7299), .op(n7300) );
  xnor2_1 U9415 ( .ip1(n7301), .ip2(n7300), .op(n7302) );
  inv_1 U9416 ( .ip(n7302), .op(n7303) );
  inv_1 U9417 ( .ip(n7831), .op(n7304) );
  nand2_1 U9418 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[3]), .ip2(
        n7304), .op(n7333) );
  inv_1 U9419 ( .ip(n7305), .op(n7307) );
  nand2_1 U9420 ( .ip1(n7307), .ip2(n7306), .op(n7309) );
  xnor2_1 U9421 ( .ip1(n7309), .ip2(n7308), .op(n7310) );
  inv_1 U9422 ( .ip(n7310), .op(n7311) );
  inv_1 U9423 ( .ip(n7832), .op(n7312) );
  nand2_1 U9424 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[2]), .ip2(
        n7312), .op(n7330) );
  inv_1 U9425 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[2]), .op(
        n11062) );
  nand2_1 U9426 ( .ip1(n7832), .ip2(n11062), .op(n7836) );
  inv_1 U9427 ( .ip(n7313), .op(n7315) );
  nand2_1 U9428 ( .ip1(n7315), .ip2(n7314), .op(n7317) );
  xor2_1 U9429 ( .ip1(n7317), .ip2(n7316), .op(n7318) );
  inv_1 U9430 ( .ip(n7324), .op(n7319) );
  nand2_1 U9431 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[1]), .ip2(
        n7319), .op(n7328) );
  xnor2_1 U9432 ( .ip1(i_i2c_ic_sda_tx_hold_sync[0]), .ip2(n7320), .op(n7322)
         );
  inv_1 U9433 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[0]), .op(
        n7358) );
  inv_1 U9434 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[1]), .op(
        n11058) );
  nand2_1 U9435 ( .ip1(n7324), .ip2(n11058), .op(n7325) );
  nand2_1 U9436 ( .ip1(n7326), .ip2(n7325), .op(n7327) );
  nand2_1 U9437 ( .ip1(n7328), .ip2(n7327), .op(n7833) );
  nand2_1 U9438 ( .ip1(n7836), .ip2(n7833), .op(n7329) );
  nand2_1 U9439 ( .ip1(n7330), .ip2(n7329), .op(n7331) );
  inv_1 U9440 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[3]), .op(
        n11067) );
  nand2_1 U9441 ( .ip1(n7831), .ip2(n11067), .op(n7842) );
  nand2_1 U9442 ( .ip1(n7331), .ip2(n7842), .op(n7332) );
  nand2_1 U9443 ( .ip1(n7333), .ip2(n7332), .op(n7334) );
  nand2_1 U9444 ( .ip1(n7848), .ip2(n7334), .op(n7335) );
  nand2_1 U9445 ( .ip1(n7336), .ip2(n7335), .op(n7337) );
  nand2_1 U9446 ( .ip1(n7829), .ip2(n7337), .op(n7338) );
  nand2_1 U9447 ( .ip1(n7339), .ip2(n7338), .op(n7340) );
  inv_1 U9448 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[6]), .op(
        n11076) );
  nand2_1 U9449 ( .ip1(n7828), .ip2(n11076), .op(n7856) );
  nand2_1 U9450 ( .ip1(n7340), .ip2(n7856), .op(n7341) );
  nand2_1 U9451 ( .ip1(n7342), .ip2(n7341), .op(n7344) );
  inv_1 U9452 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[8]), .op(
        n11082) );
  not_ab_or_c_or_d U9453 ( .ip1(n7882), .ip2(n7344), .ip3(n7881), .ip4(n7857), 
        .op(n7345) );
  not_ab_or_c_or_d U9454 ( .ip1(n7893), .ip2(n11086), .ip3(n7346), .ip4(n7345), 
        .op(n7348) );
  not_ab_or_c_or_d U9455 ( .ip1(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[9]), .ip2(n7349), .ip3(
        n7348), .ip4(n7347), .op(n7350) );
  not_ab_or_c_or_d U9456 ( .ip1(n7887), .ip2(n11094), .ip3(n7351), .ip4(n7350), 
        .op(n7352) );
  not_ab_or_c_or_d U9457 ( .ip1(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[13]), .ip2(n7353), .ip3(
        n7352), .ip4(n7888), .op(n10422) );
  nand2_1 U9458 ( .ip1(n7354), .ip2(n11102), .op(n7864) );
  inv_1 U9459 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[13]), .op(
        n11098) );
  nand2_1 U9460 ( .ip1(n7871), .ip2(n11098), .op(n7865) );
  nand2_1 U9461 ( .ip1(n7864), .ip2(n7865), .op(n10421) );
  nor2_1 U9462 ( .ip1(n10422), .ip2(n10421), .op(n7355) );
  nor2_1 U9463 ( .ip1(n10427), .ip2(n7355), .op(n7356) );
  nor2_1 U9464 ( .ip1(n10423), .ip2(n7356), .op(n7357) );
  nand3_1 U9465 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_empty_n), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_rd_addr_at_max), .ip3(
        i_i2c_tx_pop_sync), .op(n7359) );
  nand2_1 U9466 ( .ip1(i_i2c_tx_fifo_rst_n), .ip2(n7359), .op(n11249) );
  inv_1 U9467 ( .ip(i_i2c_tx_rd_addr[0]), .op(n9456) );
  nor2_1 U9468 ( .ip1(n9456), .ip2(n8213), .op(n8212) );
  nor2_1 U9469 ( .ip1(i_i2c_tx_rd_addr[1]), .ip2(n8212), .op(n8423) );
  nand2_1 U9470 ( .ip1(i_i2c_tx_rd_addr[1]), .ip2(i_i2c_tx_rd_addr[0]), .op(
        n9464) );
  nor2_1 U9471 ( .ip1(n9464), .ip2(n8213), .op(n11250) );
  nor3_1 U9472 ( .ip1(n11249), .ip2(n8423), .ip3(n11250), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N45) );
  nand3_1 U9473 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_old_is_read), .ip2(n6470), 
        .ip3(i_i2c_U_DW_apb_i2c_mstfsm_N487), .op(n7360) );
  nand2_1 U9474 ( .ip1(n7361), .ip2(n7360), .op(n5208) );
  inv_1 U9475 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[0]), .op(
        n7386) );
  nor2_1 U9476 ( .ip1(n7362), .ip2(n7386), .op(n8250) );
  inv_1 U9477 ( .ip(i_i2c_ic_hs_spklen[4]), .op(n7363) );
  nand2_1 U9478 ( .ip1(n5317), .ip2(n7363), .op(n7364) );
  nand2_1 U9479 ( .ip1(n7365), .ip2(n7364), .op(n7378) );
  nand2_1 U9480 ( .ip1(i_i2c_ic_hs_spklen[0]), .ip2(n7386), .op(n7366) );
  nand2_1 U9481 ( .ip1(n7367), .ip2(n7366), .op(n7374) );
  inv_1 U9482 ( .ip(n7368), .op(n7369) );
  nor2_1 U9483 ( .ip1(n7370), .ip2(n7369), .op(n7373) );
  nand2_1 U9484 ( .ip1(i_i2c_ic_hs_spklen[4]), .ip2(n10558), .op(n7371) );
  nand2_1 U9485 ( .ip1(n7379), .ip2(n7371), .op(n7372) );
  not_ab_or_c_or_d U9486 ( .ip1(n7375), .ip2(n7374), .ip3(n7373), .ip4(n7372), 
        .op(n7377) );
  not_ab_or_c_or_d U9487 ( .ip1(n7379), .ip2(n7378), .ip3(n7377), .ip4(n7376), 
        .op(n7383) );
  and2_1 U9488 ( .ip1(n7381), .ip2(n7380), .op(n7382) );
  nor2_1 U9489 ( .ip1(n7383), .ip2(n7382), .op(n7385) );
  nand2_1 U9490 ( .ip1(i_i2c_ic_fs_spklen[0]), .ip2(n7386), .op(n7392) );
  inv_1 U9491 ( .ip(n7387), .op(n7391) );
  inv_1 U9492 ( .ip(n7388), .op(n7390) );
  not_ab_or_c_or_d U9493 ( .ip1(n7392), .ip2(n7391), .ip3(n7390), .ip4(n7389), 
        .op(n7408) );
  inv_1 U9494 ( .ip(n7400), .op(n7397) );
  inv_1 U9495 ( .ip(n7393), .op(n7395) );
  not_ab_or_c_or_d U9496 ( .ip1(n7397), .ip2(n7396), .ip3(n7395), .ip4(n7394), 
        .op(n7407) );
  inv_1 U9497 ( .ip(n7398), .op(n7399) );
  nor2_1 U9498 ( .ip1(n7400), .ip2(n7399), .op(n7402) );
  inv_1 U9499 ( .ip(n7407), .op(n7401) );
  nor2_1 U9500 ( .ip1(n7402), .ip2(n7401), .op(n7406) );
  nor2_1 U9501 ( .ip1(n5319), .ip2(n7411), .op(n7403) );
  or2_1 U9502 ( .ip1(n7404), .ip2(n7403), .op(n7405) );
  not_ab_or_c_or_d U9503 ( .ip1(n7408), .ip2(n7407), .ip3(n7406), .ip4(n7405), 
        .op(n7409) );
  not_ab_or_c_or_d U9504 ( .ip1(n5319), .ip2(n7411), .ip3(n7410), .ip4(n7409), 
        .op(n7412) );
  xor2_1 U9505 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_scl_clk_int), .ip2(n8437), 
        .op(n7414) );
  nor3_1 U9506 ( .ip1(n7415), .ip2(n8250), .ip3(n10561), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_N83) );
  inv_1 U9507 ( .ip(i_i2c_scl_s_setup_cmplt), .op(n8310) );
  nand2_1 U9508 ( .ip1(n7740), .ip2(n8310), .op(n8306) );
  inv_1 U9509 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl), .op(n7416) );
  nor2_1 U9510 ( .ip1(n7741), .ip2(n7416), .op(n7418) );
  not_ab_or_c_or_d U9511 ( .ip1(i_i2c_scl_s_hld_cmplt), .ip2(n8310), .ip3(
        n6616), .ip4(n11119), .op(n7417) );
  inv_1 U9512 ( .ip(i_i2c_re_start_en), .op(n8443) );
  or2_1 U9513 ( .ip1(n7418), .ip2(n7743), .op(n4961) );
  inv_1 U9514 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[3]), .op(n7745)
         );
  nor3_1 U9515 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[2]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[1]), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[0]), .op(n11172) );
  nor2_1 U9516 ( .ip1(n7745), .ip2(n11172), .op(n7419) );
  inv_1 U9517 ( .ip(i_i2c_debug_wr), .op(n11156) );
  nand3_1 U9518 ( .ip1(i_i2c_scl_lcnt_cmplt), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_data_scl_lcnt_en), .ip3(i_i2c_scl_hcnt_en), 
        .op(n7428) );
  nor3_1 U9519 ( .ip1(n9096), .ip2(i_i2c_mst_rxbyte_rdy), .ip3(n8329), .op(
        n11770) );
  and3_1 U9520 ( .ip1(i_i2c_mst_rx_ack_vld), .ip2(n11770), .ip3(
        i_i2c_U_DW_apb_i2c_mstfsm_mst_gen_ack_en_r), .op(n7426) );
  inv_1 U9521 ( .ip(i_i2c_s_det), .op(n10801) );
  ab_or_c_or_d U9522 ( .ip1(n11302), .ip2(n10801), .ip3(n8551), .ip4(n11301), 
        .op(n7423) );
  nand2_1 U9523 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_ic_enable_sync_vld), .ip2(
        n7423), .op(n7918) );
  inv_1 U9524 ( .ip(i_i2c_slv_rx_ack_vld), .op(n7424) );
  nor3_1 U9525 ( .ip1(i_i2c_scl_lcnt_cmplt), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[3]), .ip3(n11152), .op(n11173) );
  inv_1 U9526 ( .ip(n11173), .op(n7427) );
  nor2_1 U9527 ( .ip1(n9999), .ip2(n7427), .op(n7430) );
  nand2_1 U9528 ( .ip1(n11152), .ip2(n7428), .op(n7695) );
  nand2_1 U9529 ( .ip1(n7429), .ip2(n7695), .op(n10583) );
  nor2_1 U9530 ( .ip1(n7430), .ip2(n10583), .op(n7431) );
  nor2_1 U9531 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_data_scl_lcnt_en), .ip2(
        n7431), .op(n7432) );
  nor2_1 U9532 ( .ip1(n8523), .ip2(n7432), .op(n4148) );
  inv_1 U9533 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[9]), .op(
        n7438) );
  nor2_1 U9534 ( .ip1(n7438), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[9]), .op(n7437) );
  not_ab_or_c_or_d U9535 ( .ip1(n7438), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[9]), .ip3(
        i_i2c_ic_tx_abrt_source[9]), .ip4(n7437), .op(n7439) );
  nor2_1 U9536 ( .ip1(n7488), .ip2(n7439), .op(n4698) );
  inv_1 U9537 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[2]), .op(
        n7441) );
  nor2_1 U9538 ( .ip1(n7441), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[2]), .op(n7440) );
  not_ab_or_c_or_d U9539 ( .ip1(n7441), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[2]), .ip3(
        i_i2c_ic_tx_abrt_source[2]), .ip4(n7440), .op(n7442) );
  nor2_1 U9540 ( .ip1(n7488), .ip2(n7442), .op(n4705) );
  inv_1 U9541 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[0]), .op(
        n7444) );
  nor2_1 U9542 ( .ip1(n7444), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[0]), .op(n7443) );
  not_ab_or_c_or_d U9543 ( .ip1(n7444), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[0]), .ip3(
        i_i2c_ic_tx_abrt_source[0]), .ip4(n7443), .op(n7445) );
  nor2_1 U9544 ( .ip1(n7488), .ip2(n7445), .op(n4707) );
  inv_1 U9545 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[12]), .op(
        n7447) );
  nor2_1 U9546 ( .ip1(n7447), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[12]), .op(n7446) );
  not_ab_or_c_or_d U9547 ( .ip1(n7447), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[12]), .ip3(
        i_i2c_ic_tx_abrt_source[12]), .ip4(n7446), .op(n7448) );
  nor2_1 U9548 ( .ip1(n7488), .ip2(n7448), .op(n4695) );
  inv_1 U9549 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[8]), .op(
        n7450) );
  nor2_1 U9550 ( .ip1(n7450), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[8]), .op(n7449) );
  not_ab_or_c_or_d U9551 ( .ip1(n7450), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[8]), .ip3(
        i_i2c_ic_tx_abrt_source[8]), .ip4(n7449), .op(n7451) );
  nor2_1 U9552 ( .ip1(n7488), .ip2(n7451), .op(n4699) );
  inv_1 U9553 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[3]), .op(
        n7453) );
  nor2_1 U9554 ( .ip1(n7453), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[3]), .op(n7452) );
  not_ab_or_c_or_d U9555 ( .ip1(n7453), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[3]), .ip3(
        i_i2c_ic_tx_abrt_source[3]), .ip4(n7452), .op(n7454) );
  nor2_1 U9556 ( .ip1(n7488), .ip2(n7454), .op(n4704) );
  inv_1 U9557 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[6]), .op(
        n7456) );
  nor2_1 U9558 ( .ip1(n7456), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[6]), .op(n7455) );
  not_ab_or_c_or_d U9559 ( .ip1(n7456), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[6]), .ip3(
        i_i2c_ic_tx_abrt_source[6]), .ip4(n7455), .op(n7457) );
  nor2_1 U9560 ( .ip1(n7488), .ip2(n7457), .op(n4701) );
  inv_1 U9561 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[14]), .op(
        n7459) );
  nor2_1 U9562 ( .ip1(n7459), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[14]), .op(n7458) );
  not_ab_or_c_or_d U9563 ( .ip1(n7459), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[14]), .ip3(
        i_i2c_ic_tx_abrt_source[14]), .ip4(n7458), .op(n7460) );
  nor2_1 U9564 ( .ip1(n7488), .ip2(n7460), .op(n4693) );
  inv_1 U9565 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[11]), .op(
        n7462) );
  nor2_1 U9566 ( .ip1(n7462), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[11]), .op(n7461) );
  not_ab_or_c_or_d U9567 ( .ip1(n7462), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[11]), .ip3(
        i_i2c_ic_tx_abrt_source[11]), .ip4(n7461), .op(n7463) );
  nor2_1 U9568 ( .ip1(n7488), .ip2(n7463), .op(n4696) );
  inv_1 U9569 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[5]), .op(
        n7465) );
  nor2_1 U9570 ( .ip1(n7465), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[5]), .op(n7464) );
  not_ab_or_c_or_d U9571 ( .ip1(n7465), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[5]), .ip3(
        i_i2c_ic_tx_abrt_source[5]), .ip4(n7464), .op(n7466) );
  nor2_1 U9572 ( .ip1(n7488), .ip2(n7466), .op(n4702) );
  inv_1 U9573 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[10]), .op(
        n7468) );
  nor2_1 U9574 ( .ip1(n7468), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[10]), .op(n7467) );
  not_ab_or_c_or_d U9575 ( .ip1(n7468), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[10]), .ip3(
        i_i2c_ic_tx_abrt_source[10]), .ip4(n7467), .op(n7469) );
  nor2_1 U9576 ( .ip1(n7488), .ip2(n7469), .op(n4697) );
  inv_1 U9577 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[4]), .op(
        n7471) );
  nor2_1 U9578 ( .ip1(n7471), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[4]), .op(n7470) );
  not_ab_or_c_or_d U9579 ( .ip1(n7471), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[4]), .ip3(
        i_i2c_ic_tx_abrt_source[4]), .ip4(n7470), .op(n7472) );
  nor2_1 U9580 ( .ip1(n7488), .ip2(n7472), .op(n4703) );
  inv_1 U9581 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[7]), .op(
        n7474) );
  nor2_1 U9582 ( .ip1(n7474), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[7]), .op(n7473) );
  not_ab_or_c_or_d U9583 ( .ip1(n7474), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[7]), .ip3(
        i_i2c_ic_tx_abrt_source[7]), .ip4(n7473), .op(n7475) );
  nor2_1 U9584 ( .ip1(n7488), .ip2(n7475), .op(n4700) );
  inv_1 U9585 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[13]), .op(
        n7477) );
  nor2_1 U9586 ( .ip1(n7477), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[13]), .op(n7476) );
  not_ab_or_c_or_d U9587 ( .ip1(n7477), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[13]), .ip3(
        i_i2c_ic_tx_abrt_source[13]), .ip4(n7476), .op(n7478) );
  nor2_1 U9588 ( .ip1(n7488), .ip2(n7478), .op(n4694) );
  inv_1 U9589 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[1]), .op(
        n7480) );
  nor2_1 U9590 ( .ip1(n7480), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[1]), .op(n7479) );
  not_ab_or_c_or_d U9591 ( .ip1(n7480), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[1]), .ip3(
        i_i2c_ic_tx_abrt_source[1]), .ip4(n7479), .op(n7481) );
  nor2_1 U9592 ( .ip1(n7488), .ip2(n7481), .op(n4706) );
  inv_1 U9593 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[15]), .op(
        n7483) );
  nor2_1 U9594 ( .ip1(n7483), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[15]), .op(n7482) );
  not_ab_or_c_or_d U9595 ( .ip1(n7483), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[15]), .ip3(
        i_i2c_ic_tx_abrt_source[15]), .ip4(n7482), .op(n7484) );
  nor2_1 U9596 ( .ip1(n7488), .ip2(n7484), .op(n4692) );
  inv_1 U9597 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[16]), .op(
        n7486) );
  nor2_1 U9598 ( .ip1(n7486), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[16]), .op(n7485) );
  not_ab_or_c_or_d U9599 ( .ip1(n7486), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[16]), .ip3(
        i_i2c_ic_tx_abrt_source[16]), .ip4(n7485), .op(n7487) );
  nor2_1 U9600 ( .ip1(n7488), .ip2(n7487), .op(n5219) );
  nand2_1 U9601 ( .ip1(i_i2c_tx_full), .ip2(n11261), .op(n7489) );
  nor2_1 U9602 ( .ip1(i_i2c_tx_wr_addr[0]), .ip2(n9766), .op(n7491) );
  nand2_1 U9603 ( .ip1(n9766), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_wr_addr_at_max), .op(n7490) );
  nand2_1 U9604 ( .ip1(i_i2c_tx_fifo_rst_n), .ip2(n7490), .op(n11254) );
  not_ab_or_c_or_d U9605 ( .ip1(i_i2c_tx_wr_addr[0]), .ip2(n9766), .ip3(n7491), 
        .ip4(n11254), .op(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N41) );
  nor2_1 U9606 ( .ip1(n11053), .ip2(n9182), .op(n7492) );
  not_ab_or_c_or_d U9607 ( .ip1(n11053), .ip2(
        i_i2c_U_DW_apb_i2c_mstfsm_abrt_in_idle), .ip3(
        i_i2c_U_DW_apb_i2c_mstfsm_mst_tx_flush), .ip4(n7492), .op(n7495) );
  inv_1 U9608 ( .ip(i_i2c_slv_ack_det), .op(n9154) );
  or2_1 U9609 ( .ip1(n8344), .ip2(n8302), .op(n7494) );
  or2_1 U9610 ( .ip1(n5245), .ip2(n8302), .op(n7493) );
  nand3_1 U9611 ( .ip1(i_i2c_ic_enable_sync), .ip2(n9732), .ip3(n8428), .op(
        n8264) );
  nor2_1 U9612 ( .ip1(n7495), .ip2(n8264), .op(n4864) );
  fulladder U9613 ( .a(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[4]), .b(n9927), 
        .ci(n7496), .co(n7062), .s(n7497) );
  nand2_1 U9614 ( .ip1(n7497), .ip2(n9930), .op(n7499) );
  nand2_1 U9615 ( .ip1(n9932), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[4]), .op(n7498) );
  nand2_1 U9616 ( .ip1(n7499), .ip2(n7498), .op(n4138) );
  nor2_1 U9617 ( .ip1(i_apb_pwdata_int[5]), .ip2(n9837), .op(n7502) );
  nor2_1 U9618 ( .ip1(i_apb_pwdata_int[4]), .ip2(n9837), .op(n7504) );
  nor2_1 U9619 ( .ip1(n7504), .ip2(i_ssi_U_regfile_ctrlr0_ir_int[5]), .op(
        n7501) );
  nor2_1 U9620 ( .ip1(n7502), .ip2(n7501), .op(n4593) );
  nor2_1 U9621 ( .ip1(n7502), .ip2(i_ssi_U_regfile_ctrlr0_ir_int[4]), .op(
        n7503) );
  nor2_1 U9622 ( .ip1(n7504), .ip2(n7503), .op(n4592) );
  inv_1 U9623 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[4]), .op(
        n11142) );
  nand2_1 U9624 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[1]), 
        .ip2(n7505), .op(n11140) );
  nand2_1 U9625 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[3]), 
        .ip2(n11138), .op(n11143) );
  nand2_1 U9626 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[6]), 
        .ip2(n11145), .op(n7507) );
  inv_1 U9627 ( .ip(i_ssi_reg_addr[5]), .op(n7509) );
  nand3_1 U9628 ( .ip1(i_ssi_reg_addr[4]), .ip2(n7509), .ip3(n7607), .op(n9909) );
  nand2_1 U9629 ( .ip1(i_ssi_reg_addr[1]), .ip2(i_ssi_reg_addr[2]), .op(n11616) );
  nand2_1 U9630 ( .ip1(n9832), .ip2(n11606), .op(n11636) );
  nor2_1 U9631 ( .ip1(i_ssi_reg_addr[0]), .ip2(n11636), .op(n7612) );
  inv_1 U9632 ( .ip(n9832), .op(n11697) );
  nand2_1 U9633 ( .ip1(i_ssi_prdata[31]), .ip2(n11697), .op(n7510) );
  nand2_1 U9634 ( .ip1(n7573), .ip2(n7510), .op(n4213) );
  nand2_1 U9635 ( .ip1(i_ssi_prdata[18]), .ip2(n11697), .op(n7511) );
  nand2_1 U9636 ( .ip1(n7573), .ip2(n7511), .op(n4226) );
  nand2_1 U9637 ( .ip1(i_ssi_prdata[16]), .ip2(n11697), .op(n7512) );
  nand2_1 U9638 ( .ip1(n7573), .ip2(n7512), .op(n4228) );
  nand2_1 U9639 ( .ip1(i_ssi_prdata[19]), .ip2(n11697), .op(n7513) );
  nand2_1 U9640 ( .ip1(n7573), .ip2(n7513), .op(n4225) );
  nand2_1 U9641 ( .ip1(i_ssi_prdata[23]), .ip2(n11697), .op(n7514) );
  nand2_1 U9642 ( .ip1(n7573), .ip2(n7514), .op(n4221) );
  nand2_1 U9643 ( .ip1(i_ssi_prdata[27]), .ip2(n11697), .op(n7515) );
  nand2_1 U9644 ( .ip1(n7573), .ip2(n7515), .op(n4217) );
  nand2_1 U9645 ( .ip1(i_ssi_prdata[22]), .ip2(n11697), .op(n7516) );
  nand2_1 U9646 ( .ip1(n7573), .ip2(n7516), .op(n4222) );
  nand2_1 U9647 ( .ip1(i_ssi_prdata[26]), .ip2(n11697), .op(n7517) );
  nand2_1 U9648 ( .ip1(n7573), .ip2(n7517), .op(n4218) );
  nand2_1 U9649 ( .ip1(i_ssi_prdata[30]), .ip2(n11697), .op(n7518) );
  nand2_1 U9650 ( .ip1(n7573), .ip2(n7518), .op(n4214) );
  nand2_1 U9651 ( .ip1(i_ssi_prdata[15]), .ip2(n11697), .op(n7538) );
  or2_1 U9652 ( .ip1(i_ssi_reg_addr[0]), .ip2(n11697), .op(n7520) );
  or2_1 U9653 ( .ip1(n11606), .ip2(n11697), .op(n7519) );
  nand2_1 U9654 ( .ip1(i_ssi_reg_addr[2]), .ip2(n9820), .op(n9785) );
  nand2_1 U9655 ( .ip1(i_ssi_baudr[15]), .ip2(n11691), .op(n7523) );
  nand2_1 U9656 ( .ip1(i_ssi_cfs[3]), .ip2(n11692), .op(n7522) );
  nand2_1 U9657 ( .ip1(n5394), .ip2(n11693), .op(n7521) );
  nand3_1 U9658 ( .ip1(n7523), .ip2(n7522), .ip3(n7521), .op(n7524) );
  nand2_1 U9659 ( .ip1(n11624), .ip2(n7524), .op(n7537) );
  inv_1 U9660 ( .ip(i_ssi_rx_rd_addr[2]), .op(n7531) );
  nor3_1 U9661 ( .ip1(i_ssi_rx_rd_addr[1]), .ip2(i_ssi_rx_rd_addr[0]), .ip3(
        n7531), .op(n11677) );
  nand2_1 U9662 ( .ip1(n11677), .ip2(i_ssi_U_dff_rx_mem[63]), .op(n7534) );
  nand2_1 U9663 ( .ip1(i_ssi_rx_rd_addr[1]), .ip2(i_ssi_rx_rd_addr[0]), .op(
        n11125) );
  nor2_1 U9664 ( .ip1(i_ssi_rx_rd_addr[2]), .ip2(n11125), .op(n11686) );
  inv_1 U9665 ( .ip(i_ssi_rx_rd_addr[1]), .op(n11126) );
  inv_1 U9666 ( .ip(i_ssi_rx_rd_addr[0]), .op(n11123) );
  and2_1 U9667 ( .ip1(n11675), .ip2(i_ssi_U_dff_rx_mem[15]), .op(n7530) );
  nor3_1 U9668 ( .ip1(i_ssi_rx_rd_addr[2]), .ip2(i_ssi_rx_rd_addr[1]), .ip3(
        i_ssi_rx_rd_addr[0]), .op(n11674) );
  nand2_1 U9669 ( .ip1(n11674), .ip2(i_ssi_U_dff_rx_mem[127]), .op(n7528) );
  nor3_1 U9670 ( .ip1(i_ssi_rx_rd_addr[2]), .ip2(i_ssi_rx_rd_addr[0]), .ip3(
        n11126), .op(n11678) );
  nand2_1 U9671 ( .ip1(n11678), .ip2(i_ssi_U_dff_rx_mem[95]), .op(n7527) );
  nor3_1 U9672 ( .ip1(i_ssi_rx_rd_addr[2]), .ip2(i_ssi_rx_rd_addr[1]), .ip3(
        n11123), .op(n11687) );
  nand2_1 U9673 ( .ip1(n11687), .ip2(i_ssi_U_dff_rx_mem[111]), .op(n7526) );
  nor3_1 U9674 ( .ip1(i_ssi_rx_rd_addr[0]), .ip2(n11126), .ip3(n7531), .op(
        n11676) );
  nand2_1 U9675 ( .ip1(n11676), .ip2(i_ssi_U_dff_rx_mem[31]), .op(n7525) );
  nand4_1 U9676 ( .ip1(n7528), .ip2(n7527), .ip3(n7526), .ip4(n7525), .op(
        n7529) );
  not_ab_or_c_or_d U9677 ( .ip1(i_ssi_U_dff_rx_mem[79]), .ip2(n11686), .ip3(
        n7530), .ip4(n7529), .op(n7533) );
  nor3_1 U9678 ( .ip1(i_ssi_rx_rd_addr[1]), .ip2(n7531), .ip3(n11123), .op(
        n11679) );
  nand2_1 U9679 ( .ip1(n11679), .ip2(i_ssi_U_dff_rx_mem[47]), .op(n7532) );
  nand3_1 U9680 ( .ip1(n7534), .ip2(n7533), .ip3(n7532), .op(n7535) );
  nand2_1 U9681 ( .ip1(n11782), .ip2(n7535), .op(n7536) );
  nand4_1 U9682 ( .ip1(n7573), .ip2(n7538), .ip3(n7537), .ip4(n7536), .op(
        n4229) );
  nand2_1 U9683 ( .ip1(i_ssi_prdata[11]), .ip2(n11697), .op(n7555) );
  nand2_1 U9684 ( .ip1(n6224), .ip2(n11691), .op(n7541) );
  nand2_1 U9685 ( .ip1(n11692), .ip2(i_ssi_ctrlr0[11]), .op(n7540) );
  nand2_1 U9686 ( .ip1(i_ssi_U_regfile_ctrlr1_int[11]), .ip2(n11693), .op(
        n7539) );
  nand3_1 U9687 ( .ip1(n7541), .ip2(n7540), .ip3(n7539), .op(n7542) );
  nand2_1 U9688 ( .ip1(n11624), .ip2(n7542), .op(n7554) );
  nand2_1 U9689 ( .ip1(n11674), .ip2(i_ssi_U_dff_rx_mem[123]), .op(n7551) );
  and2_1 U9690 ( .ip1(n11675), .ip2(i_ssi_U_dff_rx_mem[11]), .op(n7548) );
  nand2_1 U9691 ( .ip1(n11677), .ip2(i_ssi_U_dff_rx_mem[59]), .op(n7546) );
  nand2_1 U9692 ( .ip1(n11679), .ip2(i_ssi_U_dff_rx_mem[43]), .op(n7545) );
  nand2_1 U9693 ( .ip1(n11687), .ip2(i_ssi_U_dff_rx_mem[107]), .op(n7544) );
  nand2_1 U9694 ( .ip1(n11676), .ip2(i_ssi_U_dff_rx_mem[27]), .op(n7543) );
  nand4_1 U9695 ( .ip1(n7546), .ip2(n7545), .ip3(n7544), .ip4(n7543), .op(
        n7547) );
  not_ab_or_c_or_d U9696 ( .ip1(i_ssi_U_dff_rx_mem[91]), .ip2(n11678), .ip3(
        n7548), .ip4(n7547), .op(n7550) );
  nand2_1 U9697 ( .ip1(n11686), .ip2(i_ssi_U_dff_rx_mem[75]), .op(n7549) );
  nand3_1 U9698 ( .ip1(n7551), .ip2(n7550), .ip3(n7549), .op(n7552) );
  nand2_1 U9699 ( .ip1(n11782), .ip2(n7552), .op(n7553) );
  nand4_1 U9700 ( .ip1(n7573), .ip2(n7555), .ip3(n7554), .ip4(n7553), .op(
        n4233) );
  nand2_1 U9701 ( .ip1(n5257), .ip2(n11691), .op(n7558) );
  nand2_1 U9702 ( .ip1(n11692), .ip2(i_ssi_ctrlr0[10]), .op(n7557) );
  nand2_1 U9703 ( .ip1(i_ssi_U_regfile_ctrlr1_int[10]), .ip2(n11693), .op(
        n7556) );
  nand3_1 U9704 ( .ip1(n7558), .ip2(n7557), .ip3(n7556), .op(n7559) );
  nand2_1 U9705 ( .ip1(n11624), .ip2(n7559), .op(n7572) );
  nand2_1 U9706 ( .ip1(n11678), .ip2(i_ssi_U_dff_rx_mem[90]), .op(n7568) );
  and2_1 U9707 ( .ip1(n11675), .ip2(i_ssi_U_dff_rx_mem[10]), .op(n7565) );
  nand2_1 U9708 ( .ip1(n11676), .ip2(i_ssi_U_dff_rx_mem[26]), .op(n7563) );
  nand2_1 U9709 ( .ip1(n11677), .ip2(i_ssi_U_dff_rx_mem[58]), .op(n7562) );
  nand2_1 U9710 ( .ip1(n11686), .ip2(i_ssi_U_dff_rx_mem[74]), .op(n7561) );
  nand2_1 U9711 ( .ip1(n11674), .ip2(i_ssi_U_dff_rx_mem[122]), .op(n7560) );
  nand4_1 U9712 ( .ip1(n7563), .ip2(n7562), .ip3(n7561), .ip4(n7560), .op(
        n7564) );
  not_ab_or_c_or_d U9713 ( .ip1(i_ssi_U_dff_rx_mem[106]), .ip2(n11687), .ip3(
        n7565), .ip4(n7564), .op(n7567) );
  nand2_1 U9714 ( .ip1(n11679), .ip2(i_ssi_U_dff_rx_mem[42]), .op(n7566) );
  nand3_1 U9715 ( .ip1(n7568), .ip2(n7567), .ip3(n7566), .op(n7569) );
  nand2_1 U9716 ( .ip1(n11782), .ip2(n7569), .op(n7571) );
  nand2_1 U9717 ( .ip1(i_ssi_prdata[10]), .ip2(n11697), .op(n7570) );
  nand4_1 U9718 ( .ip1(n7573), .ip2(n7572), .ip3(n7571), .ip4(n7570), .op(
        n4234) );
  nand2_1 U9719 ( .ip1(n11674), .ip2(i_ssi_U_dff_rx_mem[126]), .op(n7582) );
  and2_1 U9720 ( .ip1(n11675), .ip2(i_ssi_U_dff_rx_mem[14]), .op(n7579) );
  nand2_1 U9721 ( .ip1(n11678), .ip2(i_ssi_U_dff_rx_mem[94]), .op(n7577) );
  nand2_1 U9722 ( .ip1(n11679), .ip2(i_ssi_U_dff_rx_mem[46]), .op(n7576) );
  nand2_1 U9723 ( .ip1(n11677), .ip2(i_ssi_U_dff_rx_mem[62]), .op(n7575) );
  nand2_1 U9724 ( .ip1(n11687), .ip2(i_ssi_U_dff_rx_mem[110]), .op(n7574) );
  nand4_1 U9725 ( .ip1(n7577), .ip2(n7576), .ip3(n7575), .ip4(n7574), .op(
        n7578) );
  not_ab_or_c_or_d U9726 ( .ip1(i_ssi_U_dff_rx_mem[78]), .ip2(n11686), .ip3(
        n7579), .ip4(n7578), .op(n7581) );
  nand2_1 U9727 ( .ip1(n11676), .ip2(i_ssi_U_dff_rx_mem[30]), .op(n7580) );
  nand3_1 U9728 ( .ip1(n7582), .ip2(n7581), .ip3(n7580), .op(n7588) );
  inv_1 U9729 ( .ip(n11624), .op(n7609) );
  inv_1 U9730 ( .ip(n11692), .op(n9847) );
  nor2_1 U9731 ( .ip1(n9847), .ip2(n9960), .op(n7584) );
  not_ab_or_c_or_d U9732 ( .ip1(n11693), .ip2(i_ssi_U_regfile_ctrlr1_int[14]), 
        .ip3(n7585), .ip4(n7584), .op(n7586) );
  nor2_1 U9733 ( .ip1(n7609), .ip2(n7586), .op(n7587) );
  not_ab_or_c_or_d U9734 ( .ip1(n11782), .ip2(n7588), .ip3(n7587), .ip4(n7612), 
        .op(n7590) );
  nand2_1 U9735 ( .ip1(i_ssi_prdata[14]), .ip2(n11697), .op(n7589) );
  nand2_1 U9736 ( .ip1(n7590), .ip2(n7589), .op(n4230) );
  nor2_1 U9737 ( .ip1(n7591), .ip2(n9900), .op(n7592) );
  not_ab_or_c_or_d U9738 ( .ip1(i_ssi_U_regfile_ctrlr1_int[7]), .ip2(n11693), 
        .ip3(n7592), .ip4(n11692), .op(n7593) );
  nor2_1 U9739 ( .ip1(n7609), .ip2(n7593), .op(n7594) );
  not_ab_or_c_or_d U9740 ( .ip1(i_ssi_prdata[7]), .ip2(n11697), .ip3(n7594), 
        .ip4(n7612), .op(n7606) );
  nand2_1 U9741 ( .ip1(n11678), .ip2(i_ssi_U_dff_rx_mem[87]), .op(n7603) );
  and2_1 U9742 ( .ip1(n11675), .ip2(i_ssi_U_dff_rx_mem[7]), .op(n7600) );
  nand2_1 U9743 ( .ip1(n11687), .ip2(i_ssi_U_dff_rx_mem[103]), .op(n7598) );
  nand2_1 U9744 ( .ip1(n11679), .ip2(i_ssi_U_dff_rx_mem[39]), .op(n7597) );
  nand2_1 U9745 ( .ip1(n11686), .ip2(i_ssi_U_dff_rx_mem[71]), .op(n7596) );
  nand2_1 U9746 ( .ip1(n11674), .ip2(i_ssi_U_dff_rx_mem[119]), .op(n7595) );
  nand4_1 U9747 ( .ip1(n7598), .ip2(n7597), .ip3(n7596), .ip4(n7595), .op(
        n7599) );
  not_ab_or_c_or_d U9748 ( .ip1(i_ssi_U_dff_rx_mem[23]), .ip2(n11676), .ip3(
        n7600), .ip4(n7599), .op(n7602) );
  nand2_1 U9749 ( .ip1(n11677), .ip2(i_ssi_U_dff_rx_mem[55]), .op(n7601) );
  nand3_1 U9750 ( .ip1(n7603), .ip2(n7602), .ip3(n7601), .op(n7604) );
  nand2_1 U9751 ( .ip1(n11782), .ip2(n7604), .op(n7605) );
  nand2_1 U9752 ( .ip1(n7606), .ip2(n7605), .op(n4237) );
  or4_1 U9753 ( .ip1(i_ssi_reg_addr[0]), .ip2(i_ssi_reg_addr[5]), .ip3(
        i_ssi_reg_addr[4]), .ip4(n7607), .op(n9829) );
  not_ab_or_c_or_d U9754 ( .ip1(n5392), .ip2(n11693), .ip3(n11576), .ip4(
        n11692), .op(n7611) );
  nand2_1 U9755 ( .ip1(i_ssi_baudr[6]), .ip2(n11691), .op(n7610) );
  inv_1 U9756 ( .ip(n11576), .op(n9855) );
  nor2_1 U9757 ( .ip1(i_ssi_U_regfile_sr_6_), .ip2(n9855), .op(n7608) );
  not_ab_or_c_or_d U9758 ( .ip1(n7611), .ip2(n7610), .ip3(n7609), .ip4(n7608), 
        .op(n7613) );
  not_ab_or_c_or_d U9759 ( .ip1(i_ssi_prdata[6]), .ip2(n11697), .ip3(n7613), 
        .ip4(n7612), .op(n7625) );
  nand2_1 U9760 ( .ip1(n11687), .ip2(i_ssi_U_dff_rx_mem[102]), .op(n7622) );
  and2_1 U9761 ( .ip1(n11675), .ip2(i_ssi_U_dff_rx_mem[6]), .op(n7619) );
  nand2_1 U9762 ( .ip1(n11679), .ip2(i_ssi_U_dff_rx_mem[38]), .op(n7617) );
  nand2_1 U9763 ( .ip1(n11677), .ip2(i_ssi_U_dff_rx_mem[54]), .op(n7616) );
  nand2_1 U9764 ( .ip1(n11676), .ip2(i_ssi_U_dff_rx_mem[22]), .op(n7615) );
  nand2_1 U9765 ( .ip1(n11674), .ip2(i_ssi_U_dff_rx_mem[118]), .op(n7614) );
  nand4_1 U9766 ( .ip1(n7617), .ip2(n7616), .ip3(n7615), .ip4(n7614), .op(
        n7618) );
  not_ab_or_c_or_d U9767 ( .ip1(i_ssi_U_dff_rx_mem[70]), .ip2(n11686), .ip3(
        n7619), .ip4(n7618), .op(n7621) );
  nand2_1 U9768 ( .ip1(n11678), .ip2(i_ssi_U_dff_rx_mem[86]), .op(n7620) );
  nand3_1 U9769 ( .ip1(n7622), .ip2(n7621), .ip3(n7620), .op(n7623) );
  nand2_1 U9770 ( .ip1(n11782), .ip2(n7623), .op(n7624) );
  nand2_1 U9771 ( .ip1(n7625), .ip2(n7624), .op(n4238) );
  nand2_1 U9772 ( .ip1(i_ssi_U_mstfsm_c_state[1]), .ip2(n5281), .op(n7627) );
  nor4_1 U9773 ( .ip1(i_ssi_tmod[0]), .ip2(n7627), .ip3(n7629), .ip4(n7626), 
        .op(n7632) );
  nor2_1 U9774 ( .ip1(i_ssi_U_mstfsm_tx_load_en_int), .ip2(n7630), .op(n7631)
         );
  nor2_1 U9775 ( .ip1(n7632), .ip2(n7631), .op(n4586) );
  nand2_1 U9776 ( .ip1(i_ssi_risr[3]), .ip2(i_ssi_imr[3]), .op(
        i_ssi_ssi_rxo_intr_n) );
  inv_1 U9777 ( .ip(n8525), .op(n8528) );
  nand3_1 U9778 ( .ip1(n8528), .ip2(n7922), .ip3(n8527), .op(
        i_i2c_U_DW_apb_i2c_slvfsm_N284) );
  inv_1 U9779 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[0]), .op(
        n11713) );
  inv_1 U9780 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[3]), .op(n8448) );
  inv_1 U9781 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[1]), .op(
        n11715) );
  inv_1 U9782 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[2]), .op(
        n11718) );
  nand3_1 U9783 ( .ip1(n8448), .ip2(n11715), .ip3(n11718), .op(n7633) );
  inv_1 U9784 ( .ip(i_i2c_slv_rxbyte_rdy), .op(n11114) );
  inv_1 U9785 ( .ip(n11301), .op(n8290) );
  nor2_1 U9786 ( .ip1(n7634), .ip2(i_i2c_slv_debug_cstate[1]), .op(n11320) );
  inv_1 U9787 ( .ip(n11320), .op(n8529) );
  not_ab_or_c_or_d U9788 ( .ip1(n8290), .ip2(n8529), .ip3(i_i2c_slv_rxbyte_rdy), .ip4(n8534), .op(n7677) );
  nand2_1 U9789 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[0]), .ip2(
        n7677), .op(n7635) );
  nand2_1 U9790 ( .ip1(n8278), .ip2(n7635), .op(n5084) );
  inv_1 U9791 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_data_d_int_0_), 
        .op(n9408) );
  mux2_1 U9792 ( .ip1(n9408), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_data_d_int_0_), .s(
        i_i2c_U_DW_apb_i2c_rx_filter_sda_data_int), .op(n7673) );
  inv_1 U9793 ( .ip(n7636), .op(n7637) );
  nor2_1 U9794 ( .ip1(n7638), .ip2(n7637), .op(n7639) );
  or2_1 U9795 ( .ip1(n7640), .ip2(n7639), .op(n7641) );
  nand2_1 U9796 ( .ip1(n7642), .ip2(n7641), .op(n7652) );
  or2_1 U9797 ( .ip1(n7643), .ip2(n7646), .op(n7649) );
  or2_1 U9798 ( .ip1(n7645), .ip2(n7644), .op(n7647) );
  or2_1 U9799 ( .ip1(n7647), .ip2(n7646), .op(n7648) );
  nand2_1 U9800 ( .ip1(n7649), .ip2(n7648), .op(n7651) );
  not_ab_or_c_or_d U9801 ( .ip1(n7653), .ip2(n7652), .ip3(n7651), .ip4(n7650), 
        .op(n7670) );
  inv_1 U9802 ( .ip(n7654), .op(n7656) );
  nand2_1 U9803 ( .ip1(n7656), .ip2(n7655), .op(n7662) );
  inv_1 U9804 ( .ip(n7657), .op(n7658) );
  nand2_1 U9805 ( .ip1(n7659), .ip2(n7658), .op(n7660) );
  nand3_1 U9806 ( .ip1(n7662), .ip2(n7661), .ip3(n7660), .op(n7663) );
  nand2_1 U9807 ( .ip1(n7664), .ip2(n7663), .op(n7667) );
  not_ab_or_c_or_d U9808 ( .ip1(n7668), .ip2(n7667), .ip3(n7666), .ip4(n7665), 
        .op(n7669) );
  ab_or_c_or_d U9809 ( .ip1(n7672), .ip2(n7671), .ip3(n7670), .ip4(n7669), 
        .op(n9405) );
  nand3_1 U9810 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[0]), 
        .ip2(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[2]), .ip3(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[1]), .op(n11268) );
  inv_1 U9811 ( .ip(n11268), .op(n11264) );
  nand3_1 U9812 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[3]), 
        .ip2(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[4]), .ip3(n11264), 
        .op(n11275) );
  nor3_1 U9813 ( .ip1(n11280), .ip2(n11276), .ip3(n11275), .op(n11278) );
  nor2_1 U9814 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[7]), 
        .ip2(n11278), .op(n7674) );
  nor2_1 U9815 ( .ip1(n11277), .ip2(n7674), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_N130) );
  nor2_1 U9816 ( .ip1(i_i2c_slv_tx_ack_vld), .ip2(n7713), .op(n7675) );
  nor2_1 U9817 ( .ip1(n11316), .ip2(n7675), .op(n5111) );
  nand2_1 U9818 ( .ip1(n6616), .ip2(i_i2c_U_DW_apb_i2c_tx_shift_stop_sda), 
        .op(n7676) );
  nand2_1 U9819 ( .ip1(i_i2c_scl_p_setup_cmplt), .ip2(n8266), .op(n7685) );
  nand3_1 U9820 ( .ip1(n11774), .ip2(n7676), .ip3(n7685), .op(n5049) );
  inv_1 U9821 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_3_), .op(
        n11115) );
  nor4_1 U9822 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[2]), 
        .ip2(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[0]), .ip3(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[1]), .ip4(n11115), 
        .op(n9600) );
  nand2_1 U9823 ( .ip1(i_i2c_sda_vld), .ip2(n11115), .op(n9569) );
  nand3_1 U9824 ( .ip1(n9608), .ip2(i_i2c_rx_slv_read), .ip3(n9569), .op(n7679) );
  nand2_1 U9825 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[0]), .ip2(
        n9638), .op(n7678) );
  nand2_1 U9826 ( .ip1(n7679), .ip2(n7678), .op(n9577) );
  and2_1 U9827 ( .ip1(n9566), .ip2(n9577), .op(
        i_i2c_U_DW_apb_i2c_rx_shift_rx_slv_read_s) );
  nor2_1 U9828 ( .ip1(i_i2c_scl_lcnt_cmplt), .ip2(i_i2c_scl_p_setup_cmplt), 
        .op(n7681) );
  nor2_1 U9829 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_stop_scl), .ip2(n8266), .op(
        n7680) );
  or2_1 U9830 ( .ip1(n7681), .ip2(n7680), .op(n7682) );
  nand2_1 U9831 ( .ip1(n11774), .ip2(n7682), .op(n5050) );
  inv_1 U9832 ( .ip(i_i2c_scl_p_setup_en), .op(n10677) );
  nand2_1 U9833 ( .ip1(n11776), .ip2(n8266), .op(n7683) );
  nand2_1 U9834 ( .ip1(n10677), .ip2(n7683), .op(n7684) );
  nand2_1 U9835 ( .ip1(i_i2c_scl_lcnt_cmplt), .ip2(n7684), .op(n7686) );
  nand2_1 U9836 ( .ip1(n7686), .ip2(n7685), .op(n7687) );
  and2_1 U9837 ( .ip1(n11774), .ip2(n7687), .op(n5068) );
  nor2_1 U9838 ( .ip1(i_i2c_scl_lcnt_cmplt), .ip2(i_i2c_mst_rx_bit_count[3]), 
        .op(n10571) );
  nor2_1 U9839 ( .ip1(n10571), .ip2(n7688), .op(n7694) );
  inv_1 U9840 ( .ip(n7689), .op(n7692) );
  inv_1 U9841 ( .ip(n7690), .op(n7691) );
  not_ab_or_c_or_d U9842 ( .ip1(n11152), .ip2(n7692), .ip3(n10566), .ip4(n7691), .op(n7693) );
  or2_1 U9843 ( .ip1(n7694), .ip2(n7693), .op(n4959) );
  inv_1 U9844 ( .ip(n11172), .op(n11168) );
  nor2_1 U9845 ( .ip1(n11168), .ip2(n7745), .op(n10574) );
  and2_1 U9846 ( .ip1(n10574), .ip2(n7695), .op(n11154) );
  nand2_1 U9847 ( .ip1(n7746), .ip2(n11154), .op(n7711) );
  nand2_1 U9848 ( .ip1(i_i2c_mst_tx_ack_vld), .ip2(n11772), .op(n7696) );
  nand2_1 U9849 ( .ip1(n7711), .ip2(n7696), .op(n4179) );
  xor2_1 U9850 ( .ip1(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_flg_sync), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_flg_sync_q), .op(
        i_i2c_tx_abrt_flg_edg) );
  inv_1 U9851 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[1]), .op(n7702)
         );
  inv_1 U9852 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[0]), .op(n8522)
         );
  nand2_1 U9853 ( .ip1(n7753), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[0]), .op(n7700) );
  mux2_1 U9854 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[1]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[3]), .s(n7702), .op(n7697) );
  nand2_1 U9855 ( .ip1(n7697), .ip2(n8522), .op(n7699) );
  nand3_1 U9856 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[0]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[2]), .ip3(n7702), .op(n7698)
         );
  nand3_1 U9857 ( .ip1(n7700), .ip2(n7699), .ip3(n7698), .op(n7701) );
  nand2_1 U9858 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[2]), .ip2(
        n7701), .op(n7707) );
  inv_1 U9859 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[2]), .op(n9629)
         );
  nand4_1 U9860 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[0]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[6]), .ip3(n9629), .ip4(n7702), 
        .op(n7706) );
  mux2_1 U9861 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[5]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[7]), .s(n7702), .op(n7703) );
  nand3_1 U9862 ( .ip1(n7703), .ip2(n9629), .ip3(n8522), .op(n7705) );
  nand3_1 U9863 ( .ip1(n7753), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[4]), .ip3(n9629), .op(n7704)
         );
  and4_1 U9864 ( .ip1(n7707), .ip2(n7706), .ip3(n7705), .ip4(n7704), .op(n7710) );
  nor2_1 U9865 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_data_sda), .ip2(n11160), 
        .op(n7709) );
  nand2_1 U9866 ( .ip1(n11173), .ip2(n7746), .op(n7708) );
  mux2_1 U9867 ( .ip1(n7710), .ip2(n7709), .s(n7708), .op(n7712) );
  nand2_1 U9868 ( .ip1(n7712), .ip2(n7711), .op(n4123) );
  inv_1 U9869 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly1), .op(n7714)
         );
  not_ab_or_c_or_d U9870 ( .ip1(i_i2c_tx_fifo_data_buf[7]), .ip2(n7714), .ip3(
        n7713), .ip4(n11316), .op(n7739) );
  nor2_1 U9871 ( .ip1(n11316), .ip2(n7714), .op(
        i_i2c_U_DW_apb_i2c_tx_shift_N403) );
  inv_1 U9872 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_q), .op(n7715) );
  nor2_1 U9873 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_qq), .ip2(n7715), 
        .op(n7718) );
  nand2_1 U9874 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv), .ip2(n7716), 
        .op(n7717) );
  inv_1 U9875 ( .ip(n11174), .op(n7720) );
  nand4_1 U9876 ( .ip1(n7720), .ip2(i_i2c_slv_tx_ready_unconn), .ip3(n11175), 
        .ip4(n7719), .op(n7721) );
  nand3_1 U9877 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_N403), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_data_sda), .ip3(n7721), .op(n7738) );
  nand3_1 U9878 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[1]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[0]), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[2]), .op(n7751) );
  inv_1 U9879 ( .ip(n7751), .op(n7724) );
  inv_1 U9880 ( .ip(i_i2c_tx_fifo_data_buf[0]), .op(n9734) );
  nor3_1 U9881 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[1]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[2]), .ip3(
        i_i2c_tx_fifo_data_buf[6]), .op(n7723) );
  nand3_1 U9882 ( .ip1(i_i2c_slv_tx_ready_unconn), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly1), .ip3(n11175), .op(
        n7722) );
  not_ab_or_c_or_d U9883 ( .ip1(n7724), .ip2(n9734), .ip3(n7723), .ip4(n7722), 
        .op(n7736) );
  nand2_1 U9884 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[1]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[0]), .op(n7725) );
  nor2_1 U9885 ( .ip1(i_i2c_tx_fifo_data_buf[4]), .ip2(n7725), .op(n7731) );
  inv_1 U9886 ( .ip(i_i2c_tx_fifo_data_buf[1]), .op(n9428) );
  nand2_1 U9887 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[1]), .ip2(
        n9428), .op(n7726) );
  inv_1 U9888 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[2]), .op(
        n11319) );
  or2_1 U9889 ( .ip1(n7726), .ip2(n11319), .op(n7729) );
  inv_1 U9890 ( .ip(i_i2c_tx_fifo_data_buf[2]), .op(n9416) );
  nand2_1 U9891 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[0]), .ip2(
        n9416), .op(n7727) );
  or2_1 U9892 ( .ip1(n7727), .ip2(n11319), .op(n7728) );
  nand2_1 U9893 ( .ip1(n7729), .ip2(n7728), .op(n7730) );
  or2_1 U9894 ( .ip1(n7731), .ip2(n7730), .op(n7734) );
  not_ab_or_c_or_d U9895 ( .ip1(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[2]), .ip2(
        i_i2c_tx_fifo_data_buf[3]), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[1]), .ip4(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[0]), .op(n7733) );
  nor3_1 U9896 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[0]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[2]), .ip3(
        i_i2c_tx_fifo_data_buf[5]), .op(n7732) );
  not_ab_or_c_or_d U9897 ( .ip1(n7751), .ip2(n7734), .ip3(n7733), .ip4(n7732), 
        .op(n7735) );
  nand3_1 U9898 ( .ip1(n7736), .ip2(n7735), .ip3(n7750), .op(n7737) );
  nand3_1 U9899 ( .ip1(n7739), .ip2(n7738), .ip3(n7737), .op(n5110) );
  nand4_1 U9900 ( .ip1(i_i2c_scl_lcnt_cmplt), .ip2(i_i2c_re_start_en), .ip3(
        n7740), .ip4(n8266), .op(n8347) );
  inv_1 U9901 ( .ip(n8348), .op(n8354) );
  nor2_1 U9902 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl_lcnt_en), .ip2(
        n8354), .op(n7742) );
  or2_1 U9903 ( .ip1(n7743), .ip2(n7742), .op(n7744) );
  nand2_1 U9904 ( .ip1(n8347), .ip2(n7744), .op(n4962) );
  nand3_1 U9905 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[2]), .ip2(
        n8563), .ip3(n7753), .op(n7749) );
  inv_1 U9906 ( .ip(n7753), .op(n9628) );
  nand2_1 U9907 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[3]), .ip2(
        n9631), .op(n7748) );
  nand2_1 U9908 ( .ip1(n7749), .ip2(n7748), .op(n4144) );
  nand2_1 U9909 ( .ip1(n5109), .ip2(n7758), .op(n7757) );
  nand4_1 U9910 ( .ip1(i_i2c_mst_rx_bit_count[0]), .ip2(
        i_i2c_mst_rx_bit_count[2]), .ip3(i_i2c_mst_rx_bit_count[1]), .ip4(
        n9612), .op(n9183) );
  nand2_1 U9911 ( .ip1(i_i2c_tx_fifo_data_buf[8]), .ip2(n9639), .op(n7756) );
  nor2_1 U9912 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[3]), .ip2(n9629), .op(n7752) );
  nand4_1 U9913 ( .ip1(n9449), .ip2(n7754), .ip3(n7753), .ip4(n7752), .op(
        n7755) );
  nand3_1 U9914 ( .ip1(n7757), .ip2(n7756), .ip3(n7755), .op(
        i_i2c_U_DW_apb_i2c_tx_shift_N74) );
  and3_1 U9915 ( .ip1(n7758), .ip2(i_i2c_slv_tx_ready_unconn), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly1), .op(n11317) );
  nor2_1 U9916 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[3]), .ip2(
        n11317), .op(n7759) );
  nor2_1 U9917 ( .ip1(n11316), .ip2(n7759), .op(n5105) );
  nor2_1 U9918 ( .ip1(n7760), .ip2(n8372), .op(i_i2c_U_DW_apb_i2c_mstfsm_N72)
         );
  not_ab_or_c_or_d U9919 ( .ip1(i_apb_pwdata_int[1]), .ip2(i_apb_pwdata_int[0]), .ip3(i_apb_pwdata_int[2]), .ip4(i_apb_pwdata_int[3]), .op(n7761) );
  inv_1 U9920 ( .ip(n9844), .op(n7764) );
  nand2_1 U9921 ( .ip1(n7764), .ip2(n5358), .op(n7763) );
  inv_1 U9922 ( .ip(n9837), .op(n7765) );
  nand2_1 U9923 ( .ip1(n7765), .ip2(i_apb_pwdata_int[3]), .op(n7762) );
  nand2_1 U9924 ( .ip1(n7763), .ip2(n7762), .op(n4591) );
  nand2_1 U9925 ( .ip1(n7764), .ip2(n5356), .op(n7767) );
  nand2_1 U9926 ( .ip1(n7765), .ip2(i_apb_pwdata_int[2]), .op(n7766) );
  nand2_1 U9927 ( .ip1(n7767), .ip2(n7766), .op(n4590) );
  nand2_1 U9928 ( .ip1(n11676), .ip2(i_ssi_U_dff_rx_mem[20]), .op(n7776) );
  and2_1 U9929 ( .ip1(n11675), .ip2(i_ssi_U_dff_rx_mem[4]), .op(n7773) );
  nand2_1 U9930 ( .ip1(n11687), .ip2(i_ssi_U_dff_rx_mem[100]), .op(n7771) );
  nand2_1 U9931 ( .ip1(n11679), .ip2(i_ssi_U_dff_rx_mem[36]), .op(n7770) );
  nand2_1 U9932 ( .ip1(n11686), .ip2(i_ssi_U_dff_rx_mem[68]), .op(n7769) );
  nand2_1 U9933 ( .ip1(n11674), .ip2(i_ssi_U_dff_rx_mem[116]), .op(n7768) );
  nand4_1 U9934 ( .ip1(n7771), .ip2(n7770), .ip3(n7769), .ip4(n7768), .op(
        n7772) );
  not_ab_or_c_or_d U9935 ( .ip1(i_ssi_U_dff_rx_mem[84]), .ip2(n11678), .ip3(
        n7773), .ip4(n7772), .op(n7775) );
  nand2_1 U9936 ( .ip1(n11677), .ip2(i_ssi_U_dff_rx_mem[52]), .op(n7774) );
  nand3_1 U9937 ( .ip1(n7776), .ip2(n7775), .ip3(n7774), .op(n7777) );
  nand2_1 U9938 ( .ip1(n11598), .ip2(n7777), .op(n7787) );
  nand3_1 U9939 ( .ip1(i_ssi_reg_addr[0]), .ip2(i_ssi_reg_addr[3]), .ip3(n7778), .op(n11615) );
  nand2_1 U9940 ( .ip1(i_ssi_baudr[4]), .ip2(n11691), .op(n7780) );
  nand2_1 U9941 ( .ip1(i_ssi_U_regfile_ctrlr1_int[4]), .ip2(n11693), .op(n7779) );
  nand2_1 U9942 ( .ip1(n7780), .ip2(n7779), .op(n7782) );
  nor2_1 U9943 ( .ip1(n9829), .ip2(n9785), .op(n7807) );
  inv_1 U9944 ( .ip(n7807), .op(n11584) );
  nand2_1 U9945 ( .ip1(i_ssi_risr[4]), .ip2(i_ssi_imr[4]), .op(
        i_ssi_ssi_rxf_intr_n) );
  nor2_1 U9946 ( .ip1(n11584), .ip2(i_ssi_ssi_rxf_intr_n), .op(n7781) );
  not_ab_or_c_or_d U9947 ( .ip1(n11587), .ip2(i_ssi_risr[4]), .ip3(n7782), 
        .ip4(n7781), .op(n7786) );
  inv_1 U9948 ( .ip(i_ssi_rx_full), .op(n11151) );
  nor2_1 U9949 ( .ip1(n9855), .ip2(n11151), .op(n7784) );
  not_ab_or_c_or_d U9950 ( .ip1(n11600), .ip2(i_ssi_imr[4]), .ip3(n11606), 
        .ip4(n7784), .op(n7785) );
  nand3_1 U9951 ( .ip1(n7787), .ip2(n7786), .ip3(n7785), .op(n7788) );
  nand2_1 U9952 ( .ip1(n11624), .ip2(n7788), .op(n7790) );
  nand2_1 U9953 ( .ip1(i_ssi_prdata[4]), .ip2(n11697), .op(n7789) );
  nand2_1 U9954 ( .ip1(n7790), .ip2(n7789), .op(n4240) );
  nand2_1 U9955 ( .ip1(n11697), .ip2(i_ssi_prdata[2]), .op(n7826) );
  nor2_1 U9956 ( .ip1(n9908), .ip2(n11615), .op(n11599) );
  nand2_1 U9957 ( .ip1(i_ssi_U_regfile_rxflr[2]), .ip2(n11599), .op(n7812) );
  inv_1 U9958 ( .ip(n11579), .op(n9846) );
  nor2_1 U9959 ( .ip1(i_ssi_U_regfile_txflr[2]), .ip2(n9846), .op(n7791) );
  or2_1 U9960 ( .ip1(n9846), .ip2(n7791), .op(n7806) );
  inv_1 U9961 ( .ip(n10384), .op(n7792) );
  nor2_1 U9962 ( .ip1(n9900), .ip2(n7792), .op(n7793) );
  not_ab_or_c_or_d U9963 ( .ip1(n5356), .ip2(n11692), .ip3(n11568), .ip4(n7793), .op(n7796) );
  inv_1 U9964 ( .ip(n11568), .op(n7794) );
  nor2_1 U9965 ( .ip1(i_ssi_mwcr[2]), .ip2(n7794), .op(n7795) );
  or2_1 U9966 ( .ip1(n7796), .ip2(n7795), .op(n7798) );
  nand2_1 U9967 ( .ip1(i_ssi_U_regfile_ctrlr1_int[2]), .ip2(n11693), .op(n7797) );
  nand2_1 U9968 ( .ip1(n7798), .ip2(n7797), .op(n7799) );
  or2_1 U9969 ( .ip1(n9852), .ip2(n7799), .op(n7801) );
  or2_1 U9970 ( .ip1(i_ssi_txftlr[2]), .ip2(n7799), .op(n7800) );
  nand2_1 U9971 ( .ip1(n7801), .ip2(n7800), .op(n7803) );
  inv_1 U9972 ( .ip(i_ssi_rxftlr[2]), .op(n11229) );
  mux2_1 U9973 ( .ip1(n7803), .ip2(n11229), .s(n11573), .op(n7804) );
  mux2_1 U9974 ( .ip1(i_ssi_U_fifo_U_tx_fifo_empty_n), .ip2(n7804), .s(n9855), 
        .op(n7805) );
  nand2_1 U9975 ( .ip1(n7806), .ip2(n7805), .op(n7810) );
  inv_1 U9976 ( .ip(i_ssi_imr[2]), .op(n8386) );
  nor2_1 U9977 ( .ip1(n11587), .ip2(n7807), .op(n7808) );
  inv_1 U9978 ( .ip(i_ssi_risr[2]), .op(n8385) );
  not_ab_or_c_or_d U9979 ( .ip1(n11615), .ip2(n8386), .ip3(n7808), .ip4(n8385), 
        .op(n7809) );
  not_ab_or_c_or_d U9980 ( .ip1(i_ssi_imr[2]), .ip2(n11600), .ip3(n7810), 
        .ip4(n7809), .op(n7811) );
  inv_1 U9981 ( .ip(n11606), .op(n9814) );
  nand3_1 U9982 ( .ip1(n7812), .ip2(n7811), .ip3(n9814), .op(n7813) );
  nand2_1 U9983 ( .ip1(n11624), .ip2(n7813), .op(n7825) );
  nand2_1 U9984 ( .ip1(i_ssi_U_dff_rx_mem[98]), .ip2(n11687), .op(n7822) );
  and2_1 U9985 ( .ip1(n11675), .ip2(i_ssi_U_dff_rx_mem[2]), .op(n7819) );
  nand2_1 U9986 ( .ip1(n11677), .ip2(i_ssi_U_dff_rx_mem[50]), .op(n7817) );
  nand2_1 U9987 ( .ip1(n11676), .ip2(i_ssi_U_dff_rx_mem[18]), .op(n7816) );
  nand2_1 U9988 ( .ip1(n11674), .ip2(i_ssi_U_dff_rx_mem[114]), .op(n7815) );
  nand2_1 U9989 ( .ip1(n11678), .ip2(i_ssi_U_dff_rx_mem[82]), .op(n7814) );
  nand4_1 U9990 ( .ip1(n7817), .ip2(n7816), .ip3(n7815), .ip4(n7814), .op(
        n7818) );
  not_ab_or_c_or_d U9991 ( .ip1(n11686), .ip2(i_ssi_U_dff_rx_mem[66]), .ip3(
        n7819), .ip4(n7818), .op(n7821) );
  nand2_1 U9992 ( .ip1(n11679), .ip2(i_ssi_U_dff_rx_mem[34]), .op(n7820) );
  nand3_1 U9993 ( .ip1(n7822), .ip2(n7821), .ip3(n7820), .op(n7823) );
  nand2_1 U9994 ( .ip1(n11782), .ip2(n7823), .op(n7824) );
  nand3_1 U9995 ( .ip1(n7826), .ip2(n7825), .ip3(n7824), .op(n4242) );
  nand2_1 U9996 ( .ip1(i_i2c_ic_sda_tx_hold_sync[1]), .ip2(n7827), .op(n7916)
         );
  nor2_1 U9997 ( .ip1(n7828), .ip2(n11076), .op(n7854) );
  inv_1 U9998 ( .ip(n7829), .op(n7852) );
  nor2_1 U9999 ( .ip1(n7830), .ip2(n11074), .op(n7850) );
  nor2_1 U10000 ( .ip1(n7831), .ip2(n11067), .op(n7840) );
  nor2_1 U10001 ( .ip1(n7832), .ip2(n11062), .op(n7834) );
  or2_1 U10002 ( .ip1(n7834), .ip2(n7833), .op(n7835) );
  and2_1 U10003 ( .ip1(n7836), .ip2(n7835), .op(n7838) );
  nor2_1 U10004 ( .ip1(n7837), .ip2(n11070), .op(n7841) );
  or2_1 U10005 ( .ip1(n7838), .ip2(n7841), .op(n7839) );
  inv_1 U10006 ( .ip(n7841), .op(n7844) );
  inv_1 U10007 ( .ip(n7842), .op(n7843) );
  nor2_1 U10008 ( .ip1(n7850), .ip2(n7849), .op(n7851) );
  nor2_1 U10009 ( .ip1(n7852), .ip2(n7851), .op(n7853) );
  or2_1 U10010 ( .ip1(n7854), .ip2(n7853), .op(n7855) );
  nand2_1 U10011 ( .ip1(n7856), .ip2(n7855), .op(n7879) );
  nor2_1 U10012 ( .ip1(n7857), .ip2(n7881), .op(n7877) );
  nor2_1 U10013 ( .ip1(n7858), .ip2(n11092), .op(n7859) );
  nor2_1 U10014 ( .ip1(n7859), .ip2(n7888), .op(n7898) );
  nor2_1 U10015 ( .ip1(n7893), .ip2(n11086), .op(n7860) );
  inv_1 U10016 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[10]), .op(
        n11089) );
  nor2_1 U10017 ( .ip1(n7892), .ip2(n11089), .op(n7894) );
  nor2_1 U10018 ( .ip1(n7860), .ip2(n7894), .op(n7861) );
  nand2_1 U10019 ( .ip1(n7898), .ip2(n7861), .op(n7876) );
  nand2_1 U10020 ( .ip1(n7863), .ip2(n7862), .op(n7870) );
  inv_1 U10021 ( .ip(n7864), .op(n7867) );
  nor2_1 U10022 ( .ip1(n10427), .ip2(n7865), .op(n7866) );
  nor2_1 U10023 ( .ip1(n7867), .ip2(n7866), .op(n7868) );
  or2_1 U10024 ( .ip1(n10425), .ip2(n7868), .op(n7869) );
  or2_1 U10025 ( .ip1(n7871), .ip2(n11098), .op(n7873) );
  inv_1 U10026 ( .ip(n10427), .op(n7872) );
  nand2_1 U10027 ( .ip1(n7873), .ip2(n7872), .op(n7874) );
  nor2_1 U10028 ( .ip1(n7874), .ip2(n10425), .op(n7875) );
  and2_1 U10029 ( .ip1(n7877), .ip2(n7886), .op(n7878) );
  nand2_1 U10030 ( .ip1(n7879), .ip2(n7878), .op(n7910) );
  nand2_1 U10031 ( .ip1(n7880), .ip2(n11082), .op(n7884) );
  or2_1 U10032 ( .ip1(n7882), .ip2(n7881), .op(n7883) );
  and2_1 U10033 ( .ip1(n7886), .ip2(n7885), .op(n7908) );
  nand2_1 U10034 ( .ip1(n7887), .ip2(n11094), .op(n7891) );
  or2_1 U10035 ( .ip1(n7889), .ip2(n7888), .op(n7890) );
  nand2_1 U10036 ( .ip1(n7892), .ip2(n11089), .op(n7897) );
  nand2_1 U10037 ( .ip1(n7893), .ip2(n11086), .op(n7895) );
  or2_1 U10038 ( .ip1(n7895), .ip2(n7894), .op(n7896) );
  and2_1 U10039 ( .ip1(n7899), .ip2(n7898), .op(n7900) );
  inv_1 U10040 ( .ip(n7902), .op(n7903) );
  and2_1 U10041 ( .ip1(n7904), .ip2(n7903), .op(n7905) );
  nor2_1 U10042 ( .ip1(n7906), .ip2(n7905), .op(n7907) );
  nor2_1 U10043 ( .ip1(n7908), .ip2(n7907), .op(n7909) );
  and2_1 U10044 ( .ip1(n7910), .ip2(n7909), .op(n7915) );
  nor2_1 U10045 ( .ip1(n7912), .ip2(n7911), .op(n7914) );
  not_ab_or_c_or_d U10046 ( .ip1(n7916), .ip2(n7915), .ip3(n7914), .ip4(n7913), 
        .op(n10061) );
  inv_1 U10047 ( .ip(n10061), .op(n7919) );
  nand2_1 U10048 ( .ip1(n11770), .ip2(
        i_i2c_U_DW_apb_i2c_mstfsm_mst_gen_ack_en_r), .op(n7917) );
  nor3_1 U10049 ( .ip1(i_i2c_slv_debug_cstate[3]), .ip2(n7921), .ip3(n8527), 
        .op(n8219) );
  and3_1 U10050 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[0]), .ip2(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[1]), .ip3(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[2]), .op(n8260) );
  nand2_1 U10051 ( .ip1(n8260), .ip2(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[3]), .op(n8244) );
  inv_1 U10052 ( .ip(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[4]), .op(
        n8231) );
  nor2_1 U10053 ( .ip1(n8244), .ip2(n8231), .op(n8253) );
  nand2_1 U10054 ( .ip1(n8253), .ip2(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[5]), .op(n11297) );
  inv_1 U10055 ( .ip(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[6]), .op(
        n11296) );
  nor2_1 U10056 ( .ip1(n11297), .ip2(n11296), .op(n11290) );
  nand2_1 U10057 ( .ip1(n11290), .ip2(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[7]), .op(n7923) );
  nand2_1 U10058 ( .ip1(n8259), .ip2(n7923), .op(n11295) );
  nand3_1 U10059 ( .ip1(n7924), .ip2(n8330), .ip3(n11295), .op(
        i_i2c_scl_hld_low_en) );
  or4_1 U10060 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv), .ip2(
        i_i2c_sda_int), .ip3(i_i2c_p_det), .ip4(n10915), .op(n10955) );
  and3_1 U10061 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[1]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[0]), .ip3(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[2]), .op(n8209) );
  inv_1 U10062 ( .ip(n7925), .op(n7926) );
  inv_1 U10063 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[12]), .op(n7976)
         );
  nor2_1 U10064 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[13]), .ip2(
        n7926), .op(n7974) );
  nor3_1 U10065 ( .ip1(n7976), .ip2(n7974), .ip3(n7977), .op(n7927) );
  nor2_1 U10066 ( .ip1(n7926), .ip2(n7927), .op(n7929) );
  nor2_1 U10067 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[13]), .ip2(
        n7927), .op(n7928) );
  or2_1 U10068 ( .ip1(n7929), .ip2(n7928), .op(n7931) );
  inv_1 U10069 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[14]), .op(n7935)
         );
  nand2_1 U10070 ( .ip1(n7934), .ip2(n7935), .op(n7930) );
  inv_1 U10071 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[15]), .op(n7936)
         );
  nand2_1 U10072 ( .ip1(n7937), .ip2(n7936), .op(n7932) );
  inv_1 U10073 ( .ip(n7932), .op(n7933) );
  nor3_1 U10074 ( .ip1(n7935), .ip2(n7934), .ip3(n7933), .op(n8000) );
  nor2_1 U10075 ( .ip1(n7937), .ip2(n7936), .op(n7999) );
  inv_1 U10076 ( .ip(n7938), .op(n7982) );
  nor2_1 U10077 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[9]), .ip2(n7982), .op(n7980) );
  inv_1 U10078 ( .ip(n7939), .op(n7968) );
  inv_1 U10079 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[6]), .op(n7964)
         );
  nor2_1 U10080 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[7]), .ip2(n7968), .op(n7962) );
  nor3_1 U10081 ( .ip1(n7964), .ip2(n7965), .ip3(n7962), .op(n7967) );
  inv_1 U10082 ( .ip(n7940), .op(n7961) );
  inv_1 U10083 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[4]), .op(n7957)
         );
  nor2_1 U10084 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[5]), .ip2(n7961), .op(n7956) );
  nor3_1 U10085 ( .ip1(n7957), .ip2(n7956), .ip3(n7958), .op(n7960) );
  inv_1 U10086 ( .ip(n7941), .op(n7954) );
  inv_1 U10087 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[2]), .op(n7951)
         );
  and2_1 U10088 ( .ip1(n7949), .ip2(n7951), .op(n7948) );
  nor2_1 U10089 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[3]), .ip2(n7954), .op(n7950) );
  inv_1 U10090 ( .ip(n7942), .op(n7945) );
  inv_1 U10091 ( .ip(n7943), .op(n7944) );
  not_ab_or_c_or_d U10092 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[1]), 
        .ip2(n7945), .ip3(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[0]), .ip4(
        n7944), .op(n7947) );
  nor2_1 U10093 ( .ip1(n7945), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[1]), .op(n7946) );
  nor3_1 U10094 ( .ip1(n7951), .ip2(n7950), .ip3(n7949), .op(n7952) );
  not_ab_or_c_or_d U10095 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[3]), 
        .ip2(n7954), .ip3(n7953), .ip4(n7952), .op(n7955) );
  not_ab_or_c_or_d U10096 ( .ip1(n7958), .ip2(n7957), .ip3(n7956), .ip4(n7955), 
        .op(n7959) );
  not_ab_or_c_or_d U10097 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[5]), 
        .ip2(n7961), .ip3(n7960), .ip4(n7959), .op(n7963) );
  not_ab_or_c_or_d U10098 ( .ip1(n7965), .ip2(n7964), .ip3(n7963), .ip4(n7962), 
        .op(n7966) );
  not_ab_or_c_or_d U10099 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[7]), 
        .ip2(n7968), .ip3(n7967), .ip4(n7966), .op(n7973) );
  inv_1 U10100 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[8]), .op(n7981)
         );
  and2_1 U10101 ( .ip1(n7979), .ip2(n7981), .op(n7972) );
  inv_1 U10102 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[10]), .op(n7990)
         );
  nand2_1 U10103 ( .ip1(n7989), .ip2(n7990), .op(n7971) );
  inv_1 U10104 ( .ip(n7969), .op(n7993) );
  nor2_1 U10105 ( .ip1(n7993), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[11]), .op(n7988) );
  inv_1 U10106 ( .ip(n7988), .op(n7970) );
  or4_1 U10107 ( .ip1(n7980), .ip2(n7973), .ip3(n7972), .ip4(n7986), .op(n7978) );
  ab_or_c_or_d U10108 ( .ip1(n7977), .ip2(n7976), .ip3(n7975), .ip4(n7974), 
        .op(n7994) );
  nor2_1 U10109 ( .ip1(n7978), .ip2(n7994), .op(n7997) );
  nor3_1 U10110 ( .ip1(n7981), .ip2(n7980), .ip3(n7979), .op(n7983) );
  nor2_1 U10111 ( .ip1(n7982), .ip2(n7983), .op(n7985) );
  nor2_1 U10112 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[9]), .ip2(n7983), .op(n7984) );
  or2_1 U10113 ( .ip1(n7985), .ip2(n7984), .op(n7987) );
  nor3_1 U10114 ( .ip1(n7990), .ip2(n7989), .ip3(n7988), .op(n7991) );
  not_ab_or_c_or_d U10115 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[11]), 
        .ip2(n7993), .ip3(n7992), .ip4(n7991), .op(n7995) );
  nor2_1 U10116 ( .ip1(n7995), .ip2(n7994), .op(n7996) );
  or2_1 U10117 ( .ip1(n7997), .ip2(n7996), .op(n7998) );
  nand2_1 U10118 ( .ip1(n8801), .ip2(n8002), .op(n8208) );
  or2_1 U10119 ( .ip1(i_i2c_ic_fs_spklen[1]), .ip2(i_i2c_ic_fs_spklen[2]), 
        .op(n8007) );
  and2_1 U10120 ( .ip1(i_i2c_ic_fs_spklen[3]), .ip2(n8007), .op(n8015) );
  and2_1 U10121 ( .ip1(i_i2c_ic_fs_spklen[4]), .ip2(n8015), .op(n8016) );
  and2_1 U10122 ( .ip1(i_i2c_ic_fs_spklen[5]), .ip2(n8016), .op(n8018) );
  and2_1 U10123 ( .ip1(i_i2c_ic_fs_spklen[6]), .ip2(n8018), .op(n8017) );
  and2_1 U10124 ( .ip1(i_i2c_ic_fs_spklen[7]), .ip2(n8017), .op(n8038) );
  nand2_1 U10125 ( .ip1(n8041), .ip2(n8090), .op(n8047) );
  nor2_1 U10126 ( .ip1(n8047), .ip2(n8051), .op(n8044) );
  nand2_1 U10127 ( .ip1(n8005), .ip2(n8004), .op(n8178) );
  nor2_2 U10128 ( .ip1(n8005), .ip2(n8004), .op(n8177) );
  or2_1 U10129 ( .ip1(n8182), .ip2(n8177), .op(n8006) );
  xor2_1 U10130 ( .ip1(i_i2c_ic_fs_spklen[3]), .ip2(n8007), .op(n8009) );
  nor2_1 U10131 ( .ip1(n8012), .ip2(n8011), .op(n8165) );
  nor2_1 U10132 ( .ip1(n8162), .ip2(n8165), .op(n8008) );
  nand2_1 U10133 ( .ip1(n8010), .ip2(n8009), .op(n8163) );
  or2_1 U10134 ( .ip1(n8169), .ip2(n8162), .op(n8013) );
  xor2_1 U10135 ( .ip1(i_i2c_ic_fs_spklen[4]), .ip2(n8015), .op(n8028) );
  xor2_1 U10136 ( .ip1(i_i2c_ic_fs_spklen[5]), .ip2(n8016), .op(n8030) );
  nor2_2 U10137 ( .ip1(n8031), .ip2(n8030), .op(n8027) );
  xor2_1 U10138 ( .ip1(i_i2c_ic_fs_spklen[7]), .ip2(n8017), .op(n8020) );
  xor2_1 U10139 ( .ip1(i_i2c_ic_fs_spklen[6]), .ip2(n8018), .op(n8022) );
  nor2_2 U10140 ( .ip1(n8023), .ip2(n8022), .op(n8125) );
  nand2_2 U10141 ( .ip1(n8129), .ip2(n5273), .op(n8033) );
  nor2_2 U10142 ( .ip1(n5452), .ip2(n8033), .op(n8019) );
  nand2_2 U10143 ( .ip1(n8154), .ip2(n8019), .op(n8037) );
  nand2_1 U10144 ( .ip1(n8021), .ip2(n8020), .op(n8130) );
  nand2_1 U10145 ( .ip1(n8023), .ip2(n8022), .op(n8136) );
  and2_1 U10146 ( .ip1(n8129), .ip2(n8024), .op(n8025) );
  nor2_2 U10147 ( .ip1(n8026), .ip2(n8025), .op(n8036) );
  inv_1 U10148 ( .ip(n8027), .op(n8148) );
  nand2_1 U10149 ( .ip1(n8029), .ip2(n8028), .op(n8152) );
  inv_1 U10150 ( .ip(n8152), .op(n8146) );
  nand2_1 U10151 ( .ip1(n8148), .ip2(n8146), .op(n8032) );
  nand3_4 U10152 ( .ip1(n8037), .ip2(n8036), .ip3(n8035), .op(n8097) );
  nand2_1 U10153 ( .ip1(n8058), .ip2(n8041), .op(n8048) );
  nor2_1 U10154 ( .ip1(n8048), .ip2(n8051), .op(n8042) );
  and2_1 U10155 ( .ip1(n8097), .ip2(n8042), .op(n8043) );
  or2_1 U10156 ( .ip1(n8044), .ip2(n8043), .op(n8045) );
  nand2_1 U10157 ( .ip1(n8880), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[15]), .op(n8055) );
  inv_1 U10158 ( .ip(n8047), .op(n8050) );
  inv_1 U10159 ( .ip(n8097), .op(n8087) );
  nor2_1 U10160 ( .ip1(n8048), .ip2(n8087), .op(n8049) );
  nand2_1 U10161 ( .ip1(n8881), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[14]), .op(n8053) );
  or2_1 U10162 ( .ip1(n8056), .ip2(n8053), .op(n8054) );
  nand2_1 U10163 ( .ip1(n8055), .ip2(n8054), .op(n8078) );
  inv_1 U10164 ( .ip(n8090), .op(n8066) );
  nor2_1 U10165 ( .ip1(n8066), .ip2(n8059), .op(n8062) );
  inv_1 U10166 ( .ip(n8058), .op(n8088) );
  nor2_1 U10167 ( .ip1(n8088), .ip2(n8059), .op(n8060) );
  and2_1 U10168 ( .ip1(n8097), .ip2(n8060), .op(n8061) );
  nand2_1 U10169 ( .ip1(n8887), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[13]), .op(n8075) );
  nor2_1 U10170 ( .ip1(n8066), .ip2(n8091), .op(n8069) );
  nor2_1 U10171 ( .ip1(n8088), .ip2(n8091), .op(n8067) );
  and2_1 U10172 ( .ip1(n8097), .ip2(n8067), .op(n8068) );
  inv_1 U10173 ( .ip(n8070), .op(n8071) );
  nand2_1 U10174 ( .ip1(n8888), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[12]), .op(n8073) );
  or2_1 U10175 ( .ip1(n8110), .ip2(n8073), .op(n8074) );
  nand2_1 U10176 ( .ip1(n8075), .ip2(n8074), .op(n8076) );
  and2_1 U10177 ( .ip1(n8112), .ip2(n8076), .op(n8077) );
  nor2_1 U10178 ( .ip1(n8078), .ip2(n8077), .op(n8117) );
  inv_1 U10179 ( .ip(n8095), .op(n8082) );
  nand2_1 U10180 ( .ip1(n8082), .ip2(n8093), .op(n8083) );
  nand2_1 U10181 ( .ip1(n5461), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[8]), .op(n8084) );
  or2_1 U10182 ( .ip1(n8118), .ip2(n8084), .op(n8086) );
  nand2_1 U10183 ( .ip1(n8897), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[9]), .op(n8085) );
  nor2_1 U10184 ( .ip1(n8093), .ip2(n8094), .op(n8099) );
  nor2_1 U10185 ( .ip1(n8095), .ip2(n8094), .op(n8096) );
  and2_1 U10186 ( .ip1(n8097), .ip2(n8096), .op(n8098) );
  inv_1 U10187 ( .ip(n8100), .op(n8101) );
  nand2_1 U10188 ( .ip1(n8817), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[11]), .op(n8108) );
  nand2_1 U10189 ( .ip1(n8895), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[10]), .op(n8105) );
  or2_1 U10190 ( .ip1(n8106), .ip2(n8105), .op(n8107) );
  nor2_1 U10191 ( .ip1(n8888), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[12]), .op(n8111) );
  nor2_1 U10192 ( .ip1(n8111), .ip2(n8110), .op(n8113) );
  nand2_1 U10193 ( .ip1(n8113), .ip2(n8112), .op(n8122) );
  nand2_1 U10194 ( .ip1(n8117), .ip2(n8116), .op(n8205) );
  nor2_1 U10195 ( .ip1(n5461), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[8]), .op(n8119) );
  nor2_1 U10196 ( .ip1(n8119), .ip2(n8118), .op(n8121) );
  nand2_1 U10197 ( .ip1(n8121), .ip2(n8120), .op(n8123) );
  nor2_1 U10198 ( .ip1(n8123), .ip2(n8122), .op(n8203) );
  nand2_1 U10199 ( .ip1(n8135), .ip2(n5273), .op(n8124) );
  nand2_1 U10200 ( .ip1(n8136), .ip2(n8124), .op(n8128) );
  nor2_1 U10201 ( .ip1(n5452), .ip2(n8125), .op(n8126) );
  and2_1 U10202 ( .ip1(n8126), .ip2(n8154), .op(n8127) );
  nand2_1 U10203 ( .ip1(n8129), .ip2(n8130), .op(n8131) );
  inv_1 U10204 ( .ip(n8921), .op(n8133) );
  nand2_1 U10205 ( .ip1(n8133), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[7]), .op(n8141) );
  nand2_1 U10206 ( .ip1(n5273), .ip2(n8136), .op(n8137) );
  nand2_1 U10207 ( .ip1(n8922), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[6]), .op(n8139) );
  or2_1 U10208 ( .ip1(n8142), .ip2(n8139), .op(n8140) );
  nand2_1 U10209 ( .ip1(n8141), .ip2(n8140), .op(n8161) );
  nor2_1 U10210 ( .ip1(n8922), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[6]), .op(n8143) );
  nor2_1 U10211 ( .ip1(n8144), .ip2(n8151), .op(n8145) );
  nand2_1 U10212 ( .ip1(n8148), .ip2(n8147), .op(n8149) );
  nand2_1 U10213 ( .ip1(n8928), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[5]), .op(n8158) );
  nor2_1 U10214 ( .ip1(n8928), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[5]), .op(n8194) );
  inv_1 U10215 ( .ip(n8151), .op(n8153) );
  nand2_1 U10216 ( .ip1(n8153), .ip2(n8152), .op(n8155) );
  nand2_1 U10217 ( .ip1(n5467), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[4]), .op(n8156) );
  or2_1 U10218 ( .ip1(n8194), .ip2(n8156), .op(n8157) );
  nand2_1 U10219 ( .ip1(n8158), .ip2(n8157), .op(n8159) );
  and2_1 U10220 ( .ip1(n8196), .ip2(n8159), .op(n8160) );
  nor2_1 U10221 ( .ip1(n8161), .ip2(n8160), .op(n8201) );
  inv_1 U10222 ( .ip(n8162), .op(n8164) );
  nand2_1 U10223 ( .ip1(n8164), .ip2(n8163), .op(n8168) );
  inv_1 U10224 ( .ip(n8165), .op(n8170) );
  nand2_1 U10225 ( .ip1(n8171), .ip2(n8170), .op(n8166) );
  nand2_1 U10226 ( .ip1(n8169), .ip2(n8166), .op(n8167) );
  nand2_1 U10227 ( .ip1(n5465), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[3]), .op(n8176) );
  nor2_1 U10228 ( .ip1(n5465), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[3]), .op(n8188) );
  nand2_1 U10229 ( .ip1(n8170), .ip2(n8169), .op(n8173) );
  inv_1 U10230 ( .ip(n8171), .op(n8172) );
  nand2_1 U10231 ( .ip1(n8935), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[2]), .op(n8174) );
  or2_1 U10232 ( .ip1(n8188), .ip2(n8174), .op(n8175) );
  nand2_1 U10233 ( .ip1(n8176), .ip2(n8175), .op(n8193) );
  inv_1 U10234 ( .ip(n8177), .op(n8179) );
  nand2_1 U10235 ( .ip1(n8179), .ip2(n8178), .op(n8180) );
  nand2_1 U10236 ( .ip1(n8939), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[1]), .op(n8187) );
  or2_1 U10237 ( .ip1(n8181), .ip2(i_i2c_ic_fs_spklen[0]), .op(n8183) );
  nand2_1 U10238 ( .ip1(n8183), .ip2(n8182), .op(n8940) );
  nor2_1 U10239 ( .ip1(n8940), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[0]), .op(n8185) );
  nor2_1 U10240 ( .ip1(n8939), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[1]), .op(n8184) );
  or2_1 U10241 ( .ip1(n8185), .ip2(n8184), .op(n8186) );
  nand2_1 U10242 ( .ip1(n8187), .ip2(n8186), .op(n8191) );
  nor2_1 U10243 ( .ip1(n8935), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[2]), .op(n8189) );
  nor2_1 U10244 ( .ip1(n8189), .ip2(n8188), .op(n8190) );
  and2_1 U10245 ( .ip1(n8191), .ip2(n8190), .op(n8192) );
  nor2_1 U10246 ( .ip1(n8193), .ip2(n8192), .op(n8199) );
  nor2_1 U10247 ( .ip1(n5467), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[4]), .op(n8195) );
  nor2_1 U10248 ( .ip1(n8195), .ip2(n8194), .op(n8197) );
  nand2_1 U10249 ( .ip1(n8197), .ip2(n8196), .op(n8198) );
  or2_1 U10250 ( .ip1(n8199), .ip2(n8198), .op(n8200) );
  nand2_1 U10251 ( .ip1(n8201), .ip2(n8200), .op(n8202) );
  and2_1 U10252 ( .ip1(n8203), .ip2(n8202), .op(n8204) );
  nor2_1 U10253 ( .ip1(n8205), .ip2(n8204), .op(n8206) );
  nor2_1 U10254 ( .ip1(i_i2c_ic_fs_sync), .ip2(i_i2c_hs_mcode_en), .op(n8962)
         );
  nand2_1 U10255 ( .ip1(n8962), .ip2(n10719), .op(n8874) );
  nand2_1 U10256 ( .ip1(n8206), .ip2(n8874), .op(n8207) );
  and2_2 U10257 ( .ip1(n8209), .ip2(n10918), .op(n10926) );
  nor2_4 U10258 ( .ip1(n10930), .ip2(n7957), .op(n10931) );
  nand2_4 U10259 ( .ip1(n10931), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[5]), .op(n10935) );
  nor2_2 U10260 ( .ip1(n10957), .ip2(n7935), .op(n10956) );
  nand2_1 U10261 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_ic_enable_sync_vld), .ip2(
        i_i2c_slv_rx_ack_vld), .op(n8211) );
  nand2_1 U10262 ( .ip1(n10915), .ip2(n8211), .op(n5088) );
  not_ab_or_c_or_d U10263 ( .ip1(n9456), .ip2(n8213), .ip3(n8212), .ip4(n11249), .op(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N44) );
  nand2_1 U10264 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_abrt_in_idle), .ip2(n8428), 
        .op(n8214) );
  nand2_1 U10265 ( .ip1(n9400), .ip2(n8214), .op(n5204) );
  nand3_1 U10266 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_addr_1byte_sent), .ip2(n8215), .ip3(i_i2c_U_DW_apb_i2c_mstfsm_N487), .op(n8216) );
  nand2_1 U10267 ( .ip1(n8217), .ip2(n8216), .op(n5207) );
  inv_1 U10268 ( .ip(n5232), .op(n8218) );
  nor2_1 U10269 ( .ip1(n8218), .ip2(n8372), .op(i_i2c_U_DW_apb_i2c_mstfsm_N76)
         );
  inv_1 U10270 ( .ip(n8286), .op(n8220) );
  nor2_1 U10271 ( .ip1(n8253), .ip2(n11293), .op(n8221) );
  nor2_1 U10272 ( .ip1(n11292), .ip2(n8221), .op(n8254) );
  nor2_1 U10273 ( .ip1(n8254), .ip2(n8231), .op(n8249) );
  inv_1 U10274 ( .ip(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[7]), .op(
        n8241) );
  nor2_1 U10275 ( .ip1(n8241), .ip2(i_i2c_ic_sda_setup[7]), .op(n8243) );
  inv_1 U10276 ( .ip(i_i2c_ic_sda_setup[5]), .op(n8238) );
  nor2_1 U10277 ( .ip1(i_i2c_ic_sda_setup[6]), .ip2(n11296), .op(n8237) );
  inv_1 U10278 ( .ip(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[3]), .op(
        n8258) );
  and2_1 U10279 ( .ip1(n8258), .ip2(i_i2c_ic_sda_setup[3]), .op(n8230) );
  inv_1 U10280 ( .ip(i_i2c_ic_sda_setup[2]), .op(n8228) );
  inv_1 U10281 ( .ip(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[1]), .op(
        n11286) );
  nor2_1 U10282 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[2]), .ip2(
        n8228), .op(n8225) );
  inv_1 U10283 ( .ip(i_i2c_ic_sda_setup[1]), .op(n8223) );
  inv_1 U10284 ( .ip(i_i2c_ic_sda_setup[0]), .op(n8222) );
  not_ab_or_c_or_d U10285 ( .ip1(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[1]), .ip2(n8223), .ip3(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[0]), .ip4(n8222), .op(
        n8224) );
  not_ab_or_c_or_d U10286 ( .ip1(i_i2c_ic_sda_setup[1]), .ip2(n11286), .ip3(
        n8225), .ip4(n8224), .op(n8227) );
  nor2_1 U10287 ( .ip1(i_i2c_ic_sda_setup[3]), .ip2(n8258), .op(n8226) );
  not_ab_or_c_or_d U10288 ( .ip1(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[2]), .ip2(n8228), .ip3(
        n8227), .ip4(n8226), .op(n8229) );
  not_ab_or_c_or_d U10289 ( .ip1(i_i2c_ic_sda_setup[4]), .ip2(n8231), .ip3(
        n8230), .ip4(n8229), .op(n8233) );
  nor2_1 U10290 ( .ip1(n8231), .ip2(i_i2c_ic_sda_setup[4]), .op(n8232) );
  nor2_1 U10291 ( .ip1(n8233), .ip2(n8232), .op(n8235) );
  nor2_1 U10292 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[5]), .ip2(
        n8238), .op(n8234) );
  nor2_1 U10293 ( .ip1(n8235), .ip2(n8234), .op(n8236) );
  not_ab_or_c_or_d U10294 ( .ip1(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[5]), .ip2(n8238), .ip3(
        n8237), .ip4(n8236), .op(n8240) );
  and2_1 U10295 ( .ip1(n11296), .ip2(i_i2c_ic_sda_setup[6]), .op(n8239) );
  not_ab_or_c_or_d U10296 ( .ip1(i_i2c_ic_sda_setup[7]), .ip2(n8241), .ip3(
        n8240), .ip4(n8239), .op(n8242) );
  inv_1 U10297 ( .ip(n8269), .op(n8246) );
  nor2_1 U10298 ( .ip1(n8244), .ip2(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[4]), .op(n8245) );
  nor2_1 U10299 ( .ip1(n8246), .ip2(n8245), .op(n8247) );
  nor2_1 U10300 ( .ip1(n8247), .ip2(n11293), .op(n8248) );
  or2_1 U10301 ( .ip1(n8249), .ip2(n8248), .op(n5214) );
  inv_1 U10302 ( .ip(n8250), .op(n10551) );
  inv_1 U10303 ( .ip(n10550), .op(n10553) );
  and2_1 U10304 ( .ip1(n5317), .ip2(n10555), .op(n10556) );
  inv_1 U10305 ( .ip(n10556), .op(n10559) );
  nor2_1 U10306 ( .ip1(n8251), .ip2(n10559), .op(n10560) );
  and2_1 U10307 ( .ip1(n5316), .ip2(n10560), .op(n10562) );
  nor2_1 U10308 ( .ip1(n5319), .ip2(n10562), .op(n8252) );
  nor2_1 U10309 ( .ip1(n8252), .ip2(n10561), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_N89) );
  nand2_1 U10310 ( .ip1(n8259), .ip2(n8253), .op(n8255) );
  mux2_1 U10311 ( .ip1(n8255), .ip2(n8254), .s(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[5]), .op(n8256) );
  inv_1 U10312 ( .ip(n11299), .op(n8273) );
  nand2_1 U10313 ( .ip1(n8256), .ip2(n8273), .op(n5213) );
  nor2_1 U10314 ( .ip1(n8260), .ip2(n11293), .op(n8257) );
  or2_1 U10315 ( .ip1(n11292), .ip2(n8257), .op(n11289) );
  nand2_1 U10316 ( .ip1(n11289), .ip2(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[3]), .op(n8262) );
  nand3_1 U10317 ( .ip1(n8260), .ip2(n8259), .ip3(n8258), .op(n8261) );
  nand3_1 U10318 ( .ip1(n8262), .ip2(n8261), .ip3(n8273), .op(n5215) );
  inv_1 U10319 ( .ip(i_i2c_U_DW_apb_i2c_sync_tx_empty_sync_r), .op(n8331) );
  nor3_1 U10320 ( .ip1(n5245), .ip2(n8331), .ip3(
        i_i2c_U_DW_apb_i2c_mstfsm_N487), .op(n8263) );
  nor2_1 U10321 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_tx_empty_hld), .ip2(n8263), 
        .op(n8265) );
  nor2_1 U10322 ( .ip1(n8265), .ip2(n8264), .op(n5036) );
  nor2_1 U10323 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_stop_scl_lcnt_en), .ip2(
        n8266), .op(n8268) );
  inv_1 U10324 ( .ip(n11774), .op(n8267) );
  nor2_1 U10325 ( .ip1(n8268), .ip2(n8267), .op(n5048) );
  inv_1 U10326 ( .ip(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[0]), .op(
        n11287) );
  nor3_1 U10327 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[1]), .ip2(
        n11293), .ip3(n11287), .op(n8276) );
  or2_1 U10328 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[0]), .ip2(
        n11293), .op(n8271) );
  or2_1 U10329 ( .ip1(n8269), .ip2(n11293), .op(n8270) );
  nand2_1 U10330 ( .ip1(n8271), .ip2(n8270), .op(n8272) );
  or2_1 U10331 ( .ip1(n11286), .ip2(n8444), .op(n8274) );
  nand2_1 U10332 ( .ip1(n8274), .ip2(n8273), .op(n8275) );
  or2_1 U10333 ( .ip1(n8276), .ip2(n8275), .op(n5217) );
  nand2_1 U10334 ( .ip1(n8447), .ip2(n11713), .op(n8277) );
  nand3_1 U10335 ( .ip1(n9566), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[1]), .ip3(n8277), .op(
        n8279) );
  or2_1 U10336 ( .ip1(n8278), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[1]), .op(n9065) );
  nand2_1 U10337 ( .ip1(n8279), .ip2(n9065), .op(n5083) );
  inv_1 U10338 ( .ip(n11167), .op(n8281) );
  nor2_1 U10339 ( .ip1(n11769), .ip2(i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_q), .op(n8280) );
  nor2_1 U10340 ( .ip1(n8281), .ip2(n8280), .op(n4177) );
  nor2_1 U10341 ( .ip1(n8551), .ip2(n11301), .op(n9721) );
  or2_1 U10342 ( .ip1(n9721), .ip2(n8282), .op(n8285) );
  inv_1 U10343 ( .ip(n8296), .op(n8283) );
  or2_1 U10344 ( .ip1(n8283), .ip2(n8282), .op(n8284) );
  nand2_1 U10345 ( .ip1(n8285), .ip2(n8284), .op(n8288) );
  and4_1 U10346 ( .ip1(n11293), .ip2(n8286), .ip3(n9721), .ip4(
        i_i2c_U_DW_apb_i2c_slvfsm_slv_tx_flush), .op(n8287) );
  or2_1 U10347 ( .ip1(n8288), .ip2(n8287), .op(n5230) );
  or2_1 U10348 ( .ip1(i_i2c_mst_activity_sync), .ip2(i_i2c_slv_activity_sync), 
        .op(i_i2c_activity) );
  inv_1 U10349 ( .ip(i_i2c_rx_addr_match), .op(n8289) );
  nor2_1 U10350 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_10bit_slv_sync_inv), .ip2(
        n8289), .op(n8432) );
  nor3_1 U10351 ( .ip1(i_i2c_slv_rxbyte_rdy), .ip2(n8534), .ip3(n8290), .op(
        n8303) );
  or2_1 U10352 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_slv_tx_flush), .ip2(n5245), 
        .op(n8292) );
  or2_1 U10353 ( .ip1(n8331), .ip2(n5245), .op(n8291) );
  nand2_1 U10354 ( .ip1(n8292), .ip2(n8291), .op(n8293) );
  nor2_1 U10355 ( .ip1(n8293), .ip2(n8330), .op(n8301) );
  nand2_1 U10356 ( .ip1(n8294), .ip2(n8296), .op(n8295) );
  or2_1 U10357 ( .ip1(i_i2c_tx_fifo_data_buf[8]), .ip2(n8531), .op(n8298) );
  or2_1 U10358 ( .ip1(n8296), .ip2(n8531), .op(n8297) );
  nand2_1 U10359 ( .ip1(n8298), .ip2(n8297), .op(n8299) );
  not_ab_or_c_or_d U10360 ( .ip1(n8539), .ip2(n8432), .ip3(n8303), .ip4(n8549), 
        .op(n8305) );
  inv_1 U10361 ( .ip(i_i2c_slv_activity), .op(n8573) );
  nand2_1 U10362 ( .ip1(n10915), .ip2(n8573), .op(n8304) );
  nand2_1 U10363 ( .ip1(i_i2c_ic_slave_en_sync), .ip2(n8304), .op(n8555) );
  nor2_1 U10364 ( .ip1(n8305), .ip2(n8555), .op(i_i2c_U_DW_apb_i2c_slvfsm_N37)
         );
  nor2_1 U10365 ( .ip1(n6616), .ip2(n8306), .op(n8307) );
  nor2_1 U10366 ( .ip1(n8307), .ip2(n8443), .op(n8309) );
  nand2_1 U10367 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda), .ip2(n8348), 
        .op(n8308) );
  nand2_1 U10368 ( .ip1(n8309), .ip2(n8308), .op(n4960) );
  nand2_1 U10369 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_re_scl_s_hld_en), .ip2(
        n8348), .op(n8312) );
  nor2_1 U10370 ( .ip1(n8310), .ip2(n8347), .op(n8353) );
  inv_1 U10371 ( .ip(n8353), .op(n8311) );
  nand2_1 U10372 ( .ip1(n8312), .ip2(n8311), .op(n5196) );
  nand2_1 U10373 ( .ip1(n9930), .ip2(n8452), .op(n8314) );
  nand2_1 U10374 ( .ip1(n9932), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[0]), .op(n8313) );
  nand2_1 U10375 ( .ip1(n8314), .ip2(n8313), .op(n4142) );
  fulladder U10376 ( .a(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[1]), .b(n9927), .ci(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[0]), .co(n8362), .s(n8315) );
  nand2_1 U10377 ( .ip1(n9930), .ip2(n8315), .op(n8317) );
  nand2_1 U10378 ( .ip1(n9932), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[1]), .op(n8316) );
  nand2_1 U10379 ( .ip1(n8317), .ip2(n8316), .op(n4141) );
  inv_1 U10380 ( .ip(i_i2c_mst_rx_bit_count[2]), .op(n9643) );
  inv_1 U10381 ( .ip(n11116), .op(n8319) );
  nor2_1 U10382 ( .ip1(n10569), .ip2(n8319), .op(n8320) );
  nor2_1 U10383 ( .ip1(n8320), .ip2(n11152), .op(n8321) );
  nand2_1 U10384 ( .ip1(i_i2c_rx_scl_lcnt_en), .ip2(n8357), .op(n8325) );
  or2_1 U10385 ( .ip1(n8323), .ip2(n10566), .op(n8324) );
  nand2_1 U10386 ( .ip1(n8325), .ip2(n8324), .op(n5201) );
  or2_1 U10387 ( .ip1(n10569), .ip2(n8359), .op(n8327) );
  or2_1 U10388 ( .ip1(n9183), .ip2(n8359), .op(n8326) );
  nand2_1 U10389 ( .ip1(n8327), .ip2(n8326), .op(n5113) );
  nand2_1 U10390 ( .ip1(i_i2c_tx_wr_addr[2]), .ip2(i_i2c_tx_wr_addr[1]), .op(
        n9782) );
  inv_1 U10391 ( .ip(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N41), .op(n8328) );
  nor2_1 U10392 ( .ip1(n9782), .ip2(n8328), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N40) );
  nand2_1 U10393 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(n11050), .op(n8346) );
  not_ab_or_c_or_d U10394 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_slv_tx_flush), 
        .ip2(n8331), .ip3(n8330), .ip4(n5245), .op(n8421) );
  and2_1 U10395 ( .ip1(n8334), .ip2(n8333), .op(n9742) );
  nand3_1 U10396 ( .ip1(i_i2c_scl_s_hld_cmplt), .ip2(
        i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv), .ip3(n8340), .op(n8341) );
  nand2_1 U10397 ( .ip1(i_i2c_U_DW_apb_i2c_sync_tx_empty_int_inv), .ip2(n8344), 
        .op(n8546) );
  nor2_1 U10398 ( .ip1(n11776), .ip2(i_i2c_scl_s_setup_en), .op(n8351) );
  inv_1 U10399 ( .ip(n8347), .op(n8349) );
  nor2_1 U10400 ( .ip1(n8349), .ip2(n8348), .op(n8350) );
  nor2_1 U10401 ( .ip1(n8351), .ip2(n8350), .op(n8352) );
  nor2_1 U10402 ( .ip1(n8353), .ip2(n8352), .op(n8356) );
  nor2_1 U10403 ( .ip1(i_i2c_scl_s_setup_en), .ip2(n8354), .op(n8355) );
  nor2_1 U10404 ( .ip1(n8356), .ip2(n8355), .op(n5198) );
  nor2_1 U10405 ( .ip1(n11119), .ip2(n11152), .op(n10575) );
  nor2_1 U10406 ( .ip1(i_i2c_mst_rx_data_scl), .ip2(n10565), .op(n8358) );
  or2_1 U10407 ( .ip1(n10567), .ip2(n8358), .op(n8361) );
  inv_1 U10408 ( .ip(n8359), .op(n8360) );
  nand2_1 U10409 ( .ip1(n8361), .ip2(n8360), .op(n4937) );
  inv_1 U10410 ( .ip(i_i2c_ic_10bit_slv), .op(
        i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_slv_1_sync_N2) );
  fulladder U10411 ( .a(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[2]), .b(n9927), .ci(n8362), .co(n8368), .s(n8363) );
  nand2_1 U10412 ( .ip1(n8363), .ip2(n9930), .op(n8365) );
  nand2_1 U10413 ( .ip1(n9932), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[2]), .op(n8364) );
  nand2_1 U10414 ( .ip1(n8365), .ip2(n8364), .op(n4140) );
  inv_1 U10415 ( .ip(i_i2c_slv_addressed), .op(n8366) );
  and3_1 U10416 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv), .ip2(
        i_i2c_p_det_ifaddr_sync), .ip3(n8366), .op(n8367) );
  nor2_1 U10417 ( .ip1(n8367), .ip2(n9777), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_N241) );
  fulladder U10418 ( .a(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[3]), .b(n9927), .ci(n8368), .co(n7496), .s(n8369) );
  nand2_1 U10419 ( .ip1(n8369), .ip2(n9930), .op(n8371) );
  nand2_1 U10420 ( .ip1(n9932), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[3]), .op(n8370) );
  nand2_1 U10421 ( .ip1(n8371), .ip2(n8370), .op(n4139) );
  nand2_1 U10422 ( .ip1(i_ssi_risr[5]), .ip2(i_ssi_imr[5]), .op(
        i_ssi_ssi_mst_intr_n) );
  nand2_1 U10423 ( .ip1(n11576), .ip2(n9832), .op(n8374) );
  nand2_1 U10424 ( .ip1(n8374), .ip2(i_ssi_U_regfile_sr_6_), .op(n8377) );
  inv_1 U10425 ( .ip(i_ssi_U_regfile_multi_mst_edge), .op(n8376) );
  inv_1 U10426 ( .ip(i_ssi_fsm_multi_mst), .op(n8375) );
  and2_1 U10427 ( .ip1(n11600), .ip2(n9838), .op(n9917) );
  inv_1 U10428 ( .ip(n8378), .op(n8379) );
  nor2_1 U10429 ( .ip1(n5571), .ip2(n8379), .op(n8380) );
  nor2_1 U10430 ( .ip1(i_ssi_U_mstfsm_last_frame), .ip2(n8380), .op(n8384) );
  nor3_1 U10431 ( .ip1(n8381), .ip2(n5574), .ip3(n9684), .op(n8382) );
  nor2_1 U10432 ( .ip1(n8384), .ip2(n8383), .op(n4429) );
  nand2_1 U10433 ( .ip1(i_ssi_imr[1]), .ip2(i_ssi_risr[1]), .op(
        i_ssi_ssi_txo_intr_n) );
  nand2_1 U10434 ( .ip1(i_ssi_imr[0]), .ip2(i_ssi_risr[0]), .op(
        i_ssi_ssi_txe_intr_n) );
  nor2_1 U10435 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_st_scl_s_hld_en), .ip2(
        i_i2c_start_en), .op(n11771) );
  and2_2 U10436 ( .ip1(n10593), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[2]), .op(n10596) );
  and2_2 U10437 ( .ip1(n10596), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[3]), .op(n10599) );
  and2_2 U10438 ( .ip1(n10599), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[4]), .op(n10602) );
  and2_2 U10439 ( .ip1(n10602), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[5]), .op(n10605) );
  and2_2 U10440 ( .ip1(n10605), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[6]), .op(n10608) );
  and2_2 U10441 ( .ip1(n10608), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[7]), .op(n10611) );
  and2_2 U10442 ( .ip1(n10611), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[8]), .op(n10614) );
  and2_2 U10443 ( .ip1(n10614), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[9]), .op(n10617) );
  and2_2 U10444 ( .ip1(n10617), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[10]), .op(n10620) );
  and2_2 U10445 ( .ip1(n10620), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[11]), .op(n10623) );
  and2_1 U10446 ( .ip1(n10626), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[13]), .op(n10629) );
  and2_1 U10447 ( .ip1(n10629), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[14]), .op(n10631) );
  nand3_1 U10448 ( .ip1(i_apb_penable), .ip2(i_apb_psel_en), .ip3(i_apb_pwrite), .op(n8389) );
  nand2_1 U10449 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[6]), .op(n8393) );
  nor2_1 U10450 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(n11114), .op(n8412) );
  nand2_1 U10451 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[6]), 
        .ip2(n8412), .op(n8392) );
  nor2_1 U10452 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(i_i2c_slv_rxbyte_rdy), .op(
        n8413) );
  nand2_1 U10453 ( .ip1(i_i2c_rx_push_data[6]), .ip2(n8413), .op(n8391) );
  nand3_1 U10454 ( .ip1(n8393), .ip2(n8392), .ip3(n8391), .op(n4127) );
  nand2_1 U10455 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[5]), .op(n8396) );
  nand2_1 U10456 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[5]), 
        .ip2(n8412), .op(n8395) );
  nand2_1 U10457 ( .ip1(i_i2c_rx_push_data[5]), .ip2(n8413), .op(n8394) );
  nand3_1 U10458 ( .ip1(n8396), .ip2(n8395), .ip3(n8394), .op(n4128) );
  nand2_1 U10459 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[4]), .op(n8399) );
  nand2_1 U10460 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[4]), 
        .ip2(n8412), .op(n8398) );
  nand2_1 U10461 ( .ip1(i_i2c_rx_push_data[4]), .ip2(n8413), .op(n8397) );
  nand3_1 U10462 ( .ip1(n8399), .ip2(n8398), .ip3(n8397), .op(n4129) );
  nand2_1 U10463 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[2]), .op(n8402) );
  nand2_1 U10464 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[2]), 
        .ip2(n8412), .op(n8401) );
  nand2_1 U10465 ( .ip1(i_i2c_rx_push_data[2]), .ip2(n8413), .op(n8400) );
  nand3_1 U10466 ( .ip1(n8402), .ip2(n8401), .ip3(n8400), .op(n4131) );
  nand2_1 U10467 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[3]), .op(n8405) );
  nand2_1 U10468 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[3]), 
        .ip2(n8412), .op(n8404) );
  nand2_1 U10469 ( .ip1(i_i2c_rx_push_data[3]), .ip2(n8413), .op(n8403) );
  nand3_1 U10470 ( .ip1(n8405), .ip2(n8404), .ip3(n8403), .op(n4130) );
  nand2_1 U10471 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[1]), .op(n8408) );
  nand2_1 U10472 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[1]), 
        .ip2(n8412), .op(n8407) );
  nand2_1 U10473 ( .ip1(i_i2c_rx_push_data[1]), .ip2(n8413), .op(n8406) );
  nand3_1 U10474 ( .ip1(n8408), .ip2(n8407), .ip3(n8406), .op(n4132) );
  nand2_1 U10475 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[7]), .op(n8411) );
  nand2_1 U10476 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[7]), 
        .ip2(n8412), .op(n8410) );
  nand2_1 U10477 ( .ip1(i_i2c_rx_push_data[7]), .ip2(n8413), .op(n8409) );
  nand3_1 U10478 ( .ip1(n8411), .ip2(n8410), .ip3(n8409), .op(n4126) );
  nand2_1 U10479 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[0]), 
        .ip2(n8412), .op(n8416) );
  nand2_1 U10480 ( .ip1(i_i2c_rx_push_data[0]), .ip2(n8413), .op(n8415) );
  nand2_1 U10481 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[0]), .op(n8414) );
  nand3_1 U10482 ( .ip1(n8416), .ip2(n8415), .ip3(n8414), .op(n4133) );
  nand2_1 U10483 ( .ip1(n11320), .ip2(n8417), .op(n8420) );
  nand2_1 U10484 ( .ip1(n8418), .ip2(i_i2c_mst_rxbyte_rdy), .op(n8419) );
  nand2_1 U10485 ( .ip1(n8420), .ip2(n8419), .op(
        i_i2c_U_DW_apb_i2c_rx_shift_N30) );
  inv_1 U10486 ( .ip(n8421), .op(n8422) );
  nor2_1 U10487 ( .ip1(n8422), .ip2(n8555), .op(i_i2c_U_DW_apb_i2c_slvfsm_N39)
         );
  inv_1 U10488 ( .ip(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N44), .op(n8424) );
  inv_1 U10489 ( .ip(i_i2c_tx_rd_addr[2]), .op(n9457) );
  nor3_1 U10490 ( .ip1(n8424), .ip2(n8423), .ip3(n9457), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N39) );
  inv_1 U10491 ( .ip(n8425), .op(n8426) );
  nand2_1 U10492 ( .ip1(n8427), .ip2(n8426), .op(n8430) );
  nand2_1 U10493 ( .ip1(i_i2c_abrt_in_rcve_trns), .ip2(n8428), .op(n8429) );
  nand2_1 U10494 ( .ip1(n8430), .ip2(n8429), .op(n5190) );
  inv_1 U10495 ( .ip(i_i2c_slv_rx_2addr), .op(n9576) );
  inv_1 U10496 ( .ip(i_i2c_rx_slv_read), .op(n8538) );
  nor3_1 U10497 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_10bit_slv_sync_inv), .ip2(
        n9576), .ip3(n8538), .op(n8431) );
  not_ab_or_c_or_d U10498 ( .ip1(n11301), .ip2(n8432), .ip3(
        i_i2c_slv_addressed), .ip4(n8431), .op(n8433) );
  or2_1 U10499 ( .ip1(n8433), .ip2(n8534), .op(n8436) );
  nand3_1 U10500 ( .ip1(i_i2c_rx_addr_match), .ip2(n8447), .ip3(
        i_i2c_U_DW_apb_i2c_sync_ic_10bit_slv_sync_inv), .op(n8434) );
  or2_1 U10501 ( .ip1(n8434), .ip2(n8534), .op(n8435) );
  nand2_1 U10502 ( .ip1(n8436), .ip2(n8435), .op(n5085) );
  inv_1 U10503 ( .ip(n8439), .op(n8438) );
  nand2_1 U10504 ( .ip1(n8438), .ip2(n8437), .op(n8441) );
  nand2_1 U10505 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_scl_clk_int), .ip2(n8439), 
        .op(n8440) );
  nand2_1 U10506 ( .ip1(n8441), .ip2(n8440), .op(n5137) );
  nand2_1 U10507 ( .ip1(n8443), .ip2(n8442), .op(i_i2c_U_DW_apb_i2c_toggle_N30) );
  or2_1 U10508 ( .ip1(n11293), .ip2(n8444), .op(n8446) );
  or2_1 U10509 ( .ip1(n11287), .ip2(n8444), .op(n8445) );
  nand2_1 U10510 ( .ip1(n8446), .ip2(n8445), .op(n5218) );
  nand2_1 U10511 ( .ip1(n9566), .ip2(n9065), .op(n9066) );
  or2_1 U10512 ( .ip1(n9066), .ip2(n8448), .op(n8451) );
  nand2_1 U10513 ( .ip1(n8447), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[2]), .op(n8449) );
  or2_1 U10514 ( .ip1(n8449), .ip2(n8448), .op(n8450) );
  nand2_1 U10515 ( .ip1(n8451), .ip2(n8450), .op(n5081) );
  inv_1 U10516 ( .ip(i_i2c_ic_en), .op(n11178) );
  inv_1 U10517 ( .ip(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[1]), .op(n8459)
         );
  inv_1 U10518 ( .ip(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[0]), .op(n8452)
         );
  nor2_1 U10519 ( .ip1(i_i2c_ic_tx_tl[0]), .ip2(n8452), .op(n8453) );
  or2_1 U10520 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[1]), .ip2(n8453), .op(n8456) );
  inv_1 U10521 ( .ip(i_i2c_ic_tx_tl[1]), .op(n8454) );
  or2_1 U10522 ( .ip1(n8454), .ip2(n8453), .op(n8455) );
  nand2_1 U10523 ( .ip1(n8456), .ip2(n8455), .op(n8458) );
  nor2_1 U10524 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[2]), .ip2(
        n8461), .op(n8457) );
  not_ab_or_c_or_d U10525 ( .ip1(i_i2c_ic_tx_tl[1]), .ip2(n8459), .ip3(n8458), 
        .ip4(n8457), .op(n8460) );
  not_ab_or_c_or_d U10526 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[2]), 
        .ip2(n8461), .ip3(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[3]), .ip4(
        n8460), .op(n8463) );
  nand2_1 U10527 ( .ip1(n8463), .ip2(n8462), .op(n8464) );
  mux2_1 U10528 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_almost_empty_n), 
        .ip2(n8464), .s(i_i2c_tx_empty_ctrl), .op(n8465) );
  nor2_1 U10529 ( .ip1(n11178), .ip2(n8465), .op(i_i2c_ic_raw_intr_stat[4]) );
  nand2_1 U10530 ( .ip1(i_i2c_ic_clr_rx_over_en), .ip2(n7435), .op(n8466) );
  nand2_1 U10531 ( .ip1(i_i2c_ic_clr_intr_en), .ip2(n7435), .op(n8472) );
  nand3_1 U10532 ( .ip1(n8466), .ip2(n8472), .ip3(i_i2c_ic_raw_intr_stat[1]), 
        .op(n8467) );
  or2_1 U10533 ( .ip1(n8467), .ip2(n11178), .op(n8471) );
  inv_1 U10534 ( .ip(i_i2c_U_DW_apb_i2c_fifo_rx_pop_dly), .op(n8468) );
  nand3_1 U10535 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_rx_error_ir), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_rx_push_sync_dly), .ip3(n8468), .op(n8469) );
  or2_1 U10536 ( .ip1(n8469), .ip2(n11178), .op(n8470) );
  nand2_1 U10537 ( .ip1(n8471), .ip2(n8470), .op(n4652) );
  nand2_1 U10538 ( .ip1(i_i2c_ic_clr_rx_under_en), .ip2(n7435), .op(n8473) );
  nand3_1 U10539 ( .ip1(n8473), .ip2(n8472), .ip3(i_i2c_ic_raw_intr_stat[0]), 
        .op(n8474) );
  or2_1 U10540 ( .ip1(n8474), .ip2(n11178), .op(n8477) );
  nand3_1 U10541 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_rx_error_ir), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_rx_pop_dly), .ip3(n5247), .op(n8475) );
  or2_1 U10542 ( .ip1(n8475), .ip2(n11178), .op(n8476) );
  nand2_1 U10543 ( .ip1(n8477), .ip2(n8476), .op(n4653) );
  nand2_1 U10544 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_tx_error_ir), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_push_dly), .op(n8478) );
  nor2_1 U10545 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_tx_pop_sync_dly), .ip2(n8478), 
        .op(n8480) );
  or2_1 U10546 ( .ip1(i_i2c_ic_raw_intr_stat[3]), .ip2(n8480), .op(n8483) );
  or2_1 U10547 ( .ip1(i_i2c_ic_clr_intr_en), .ip2(i_i2c_ic_clr_tx_over_en), 
        .op(n8479) );
  nand2_1 U10548 ( .ip1(n7435), .ip2(n8479), .op(n8481) );
  or2_1 U10549 ( .ip1(n8481), .ip2(n8480), .op(n8482) );
  nand2_1 U10550 ( .ip1(n8483), .ip2(n8482), .op(n8484) );
  nor2_1 U10551 ( .ip1(n8484), .ip2(n11178), .op(n4651) );
  nor2_1 U10552 ( .ip1(i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync_q), .op(n8486) );
  inv_1 U10553 ( .ip(i_i2c_ic_ack_general_call), .op(n8485) );
  not_ab_or_c_or_d U10554 ( .ip1(
        i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync_q), .ip3(n8486), .ip4(
        n8485), .op(n8488) );
  or2_1 U10555 ( .ip1(i_i2c_ic_raw_intr_stat[11]), .ip2(n8488), .op(n8491) );
  or2_1 U10556 ( .ip1(i_i2c_ic_clr_intr_en), .ip2(i_i2c_ic_clr_gen_call_en), 
        .op(n8487) );
  nand2_1 U10557 ( .ip1(n7435), .ip2(n8487), .op(n8489) );
  or2_1 U10558 ( .ip1(n8489), .ip2(n8488), .op(n8490) );
  nand2_1 U10559 ( .ip1(n8491), .ip2(n8490), .op(n8492) );
  nor2_1 U10560 ( .ip1(n8492), .ip2(n11178), .op(n4660) );
  or2_1 U10561 ( .ip1(i_i2c_ic_raw_intr_stat[8]), .ip2(i_i2c_activity), .op(
        n8496) );
  or2_1 U10562 ( .ip1(i_i2c_ic_clr_intr_en), .ip2(i_i2c_ic_clr_activity_en), 
        .op(n8493) );
  nand2_1 U10563 ( .ip1(n7435), .ip2(n8493), .op(n8494) );
  or2_1 U10564 ( .ip1(n8494), .ip2(i_i2c_activity), .op(n8495) );
  nand2_1 U10565 ( .ip1(n8496), .ip2(n8495), .op(n8497) );
  nor2_1 U10566 ( .ip1(n8497), .ip2(n11178), .op(n4657) );
  xor2_1 U10567 ( .ip1(i_i2c_U_DW_apb_i2c_intctl_ic_rd_req_flg_sync), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_ic_rd_req_flg_sync_q), .op(n8499) );
  or2_1 U10568 ( .ip1(i_i2c_ic_raw_intr_stat[5]), .ip2(n8499), .op(n8502) );
  or2_1 U10569 ( .ip1(i_i2c_ic_clr_intr_en), .ip2(i_i2c_ic_clr_rd_req_en), 
        .op(n8498) );
  nand2_1 U10570 ( .ip1(n7435), .ip2(n8498), .op(n8500) );
  nand2_1 U10571 ( .ip1(n8502), .ip2(n8501), .op(n8503) );
  nor2_1 U10572 ( .ip1(n8503), .ip2(n11178), .op(n4654) );
  xor2_1 U10573 ( .ip1(i_i2c_U_DW_apb_i2c_intctl_rx_done_flg_sync), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_rx_done_flg_sync_q), .op(n8505) );
  or2_1 U10574 ( .ip1(i_i2c_ic_raw_intr_stat[7]), .ip2(n8505), .op(n8508) );
  or2_1 U10575 ( .ip1(i_i2c_ic_clr_intr_en), .ip2(i_i2c_ic_clr_rx_done_en), 
        .op(n8504) );
  nand2_1 U10576 ( .ip1(n7435), .ip2(n8504), .op(n8506) );
  nand2_1 U10577 ( .ip1(n8508), .ip2(n8507), .op(n8509) );
  nor2_1 U10578 ( .ip1(n8509), .ip2(n11178), .op(n4656) );
  xor2_1 U10579 ( .ip1(i_i2c_U_DW_apb_i2c_intctl_p_det_flg_sync), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_p_det_flg_sync_q), .op(n8511) );
  or2_1 U10580 ( .ip1(i_i2c_ic_raw_intr_stat[9]), .ip2(n8511), .op(n8514) );
  or2_1 U10581 ( .ip1(i_i2c_ic_clr_intr_en), .ip2(i_i2c_ic_clr_stop_det_en), 
        .op(n8510) );
  nand2_1 U10582 ( .ip1(n7435), .ip2(n8510), .op(n8512) );
  nand2_1 U10583 ( .ip1(n8514), .ip2(n8513), .op(n8515) );
  nor2_1 U10584 ( .ip1(n8515), .ip2(n11178), .op(n4659) );
  xor2_1 U10585 ( .ip1(i_i2c_U_DW_apb_i2c_intctl_s_det_flg_sync), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_s_det_flg_sync_q), .op(n8517) );
  or2_1 U10586 ( .ip1(i_i2c_ic_raw_intr_stat[10]), .ip2(n8517), .op(n8520) );
  or2_1 U10587 ( .ip1(i_i2c_ic_clr_intr_en), .ip2(i_i2c_ic_clr_start_det_en), 
        .op(n8516) );
  nand2_1 U10588 ( .ip1(n7435), .ip2(n8516), .op(n8518) );
  nand2_1 U10589 ( .ip1(n8520), .ip2(n8519), .op(n8521) );
  nor2_1 U10590 ( .ip1(n8521), .ip2(n11178), .op(n4658) );
  mux2_1 U10591 ( .ip1(n8523), .ip2(n9627), .s(n8522), .op(n8524) );
  inv_1 U10592 ( .ip(n8524), .op(n4147) );
  nand2_1 U10593 ( .ip1(i_i2c_ic_enable_sync), .ip2(i_i2c_s_det), .op(n8526)
         );
  not_ab_or_c_or_d U10594 ( .ip1(n8527), .ip2(n8526), .ip3(
        i_i2c_slv_debug_cstate[0]), .ip4(n8525), .op(n8544) );
  not_ab_or_c_or_d U10595 ( .ip1(n11292), .ip2(n9399), .ip3(n8528), .ip4(
        n10801), .op(n8532) );
  nand3_1 U10596 ( .ip1(i_i2c_slv_rxbyte_rdy), .ip2(n11301), .ip3(
        i_i2c_rx_addr_match), .op(n8530) );
  nand2_1 U10597 ( .ip1(n8530), .ip2(n8529), .op(n8553) );
  nor3_1 U10598 ( .ip1(n8532), .ip2(n8531), .ip3(n8553), .op(n8533) );
  nor2_1 U10599 ( .ip1(i_i2c_p_det), .ip2(n8533), .op(n8543) );
  nor3_1 U10600 ( .ip1(i_i2c_slv_rxbyte_rdy), .ip2(n8535), .ip3(n8534), .op(
        n8542) );
  inv_1 U10601 ( .ip(n8536), .op(n8537) );
  nand3_1 U10602 ( .ip1(i_i2c_rx_gen_call), .ip2(
        i_i2c_ic_ack_general_call_sync), .ip3(n8537), .op(n8541) );
  nand4_1 U10603 ( .ip1(i_i2c_rx_addr_match), .ip2(n8539), .ip3(
        i_i2c_U_DW_apb_i2c_sync_ic_10bit_slv_sync_inv), .ip4(n8538), .op(n8540) );
  nand2_1 U10604 ( .ip1(n8541), .ip2(n8540), .op(n8550) );
  or2_1 U10605 ( .ip1(n8545), .ip2(n8555), .op(n8548) );
  or2_1 U10606 ( .ip1(n8546), .ip2(n8555), .op(n8547) );
  nand2_1 U10607 ( .ip1(n8548), .ip2(n8547), .op(i_i2c_U_DW_apb_i2c_slvfsm_N36) );
  not_ab_or_c_or_d U10608 ( .ip1(i_i2c_s_det), .ip2(n8551), .ip3(n8550), .ip4(
        n8549), .op(n8552) );
  or2_1 U10609 ( .ip1(n8552), .ip2(n8555), .op(n8558) );
  nand2_1 U10610 ( .ip1(n8554), .ip2(n8553), .op(n8556) );
  or2_1 U10611 ( .ip1(n8556), .ip2(n8555), .op(n8557) );
  nand2_1 U10612 ( .ip1(n8558), .ip2(n8557), .op(i_i2c_U_DW_apb_i2c_slvfsm_N38) );
  or2_1 U10613 ( .ip1(i_i2c_ic_raw_intr_stat[6]), .ip2(i_i2c_tx_abrt_flg_edg), 
        .op(n8561) );
  or2_1 U10614 ( .ip1(n8559), .ip2(i_i2c_tx_abrt_flg_edg), .op(n8560) );
  nand2_1 U10615 ( .ip1(n8561), .ip2(n8560), .op(n8562) );
  nor2_1 U10616 ( .ip1(n8562), .ip2(n11178), .op(n4655) );
  inv_1 U10617 ( .ip(n9631), .op(n8567) );
  or2_1 U10618 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[0]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[1]), .op(n8565) );
  or2_1 U10619 ( .ip1(n8563), .ip2(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[1]), .op(n8564) );
  nand2_1 U10620 ( .ip1(n8565), .ip2(n8564), .op(n8566) );
  nor2_1 U10621 ( .ip1(n8567), .ip2(n8566), .op(n4146) );
  inv_1 U10622 ( .ip(i_i2c_slv_tx_ack_vld), .op(n8568) );
  nand3_1 U10623 ( .ip1(n5109), .ip2(n8569), .ip3(n8568), .op(n8571) );
  nand2_1 U10624 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_slv_arb_lost), .ip2(
        n11167), .op(n8570) );
  xor2_1 U10625 ( .ip1(i_ssi_tx_rd_addr[2]), .ip2(n8574), .op(n8575) );
  nor2_2 U10626 ( .ip1(n8576), .ip2(n8575), .op(i_ssi_U_fifo_U_tx_fifo_N46) );
  and3_1 U10627 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[2]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[0]), .ip3(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[1]), .op(n8723) );
  nand2_1 U10628 ( .ip1(n6727), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[15]), .op(n8579) );
  nor2_1 U10629 ( .ip1(n6727), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[15]), .op(n8580) );
  nand2_1 U10630 ( .ip1(n6734), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[14]), .op(n8577) );
  or2_1 U10631 ( .ip1(n8580), .ip2(n8577), .op(n8578) );
  nand2_1 U10632 ( .ip1(n8579), .ip2(n8578), .op(n8587) );
  nor2_1 U10633 ( .ip1(n6734), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[14]), .op(n8581) );
  nor2_1 U10634 ( .ip1(n8581), .ip2(n8580), .op(n8590) );
  nand2_1 U10635 ( .ip1(n8730), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[13]), .op(n8584) );
  nor2_1 U10636 ( .ip1(n8730), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[13]), .op(n8588) );
  nand2_1 U10637 ( .ip1(n6744), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[12]), .op(n8582) );
  or2_1 U10638 ( .ip1(n8588), .ip2(n8582), .op(n8583) );
  and2_1 U10639 ( .ip1(n8590), .ip2(n8585), .op(n8586) );
  nor2_1 U10640 ( .ip1(n6744), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[12]), .op(n8589) );
  nor2_1 U10641 ( .ip1(n8589), .ip2(n8588), .op(n8591) );
  nand2_1 U10642 ( .ip1(n8591), .ip2(n8590), .op(n8610) );
  nand2_1 U10643 ( .ip1(n8741), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[11]), .op(n8594) );
  nor2_1 U10644 ( .ip1(n8741), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[11]), .op(n8595) );
  nand2_1 U10645 ( .ip1(n6760), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[10]), .op(n8592) );
  or2_1 U10646 ( .ip1(n8595), .ip2(n8592), .op(n8593) );
  nand2_1 U10647 ( .ip1(n8594), .ip2(n8593), .op(n8602) );
  nor2_1 U10648 ( .ip1(n6760), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[10]), .op(n8596) );
  nor2_1 U10649 ( .ip1(n8596), .ip2(n8595), .op(n8608) );
  nand2_1 U10650 ( .ip1(n6772), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[9]), .op(n8599) );
  nor2_1 U10651 ( .ip1(n6772), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[9]), .op(n8606) );
  nand2_1 U10652 ( .ip1(n5272), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[8]), .op(n8597) );
  or2_1 U10653 ( .ip1(n8606), .ip2(n8597), .op(n8598) );
  and2_1 U10654 ( .ip1(n8608), .ip2(n8600), .op(n8601) );
  or2_1 U10655 ( .ip1(n8610), .ip2(n8603), .op(n8604) );
  nand2_1 U10656 ( .ip1(n8605), .ip2(n8604), .op(n8647) );
  nor2_1 U10657 ( .ip1(n5272), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[8]), .op(n8607) );
  nor2_1 U10658 ( .ip1(n8607), .ip2(n8606), .op(n8609) );
  nand2_1 U10659 ( .ip1(n8609), .ip2(n8608), .op(n8611) );
  nor2_1 U10660 ( .ip1(n8611), .ip2(n8610), .op(n8645) );
  nand2_1 U10661 ( .ip1(n8762), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[7]), .op(n8614) );
  nor2_1 U10662 ( .ip1(n8762), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[7]), .op(n8615) );
  nand2_1 U10663 ( .ip1(n6784), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[6]), .op(n8612) );
  or2_1 U10664 ( .ip1(n8615), .ip2(n8612), .op(n8613) );
  nor2_1 U10665 ( .ip1(n6784), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[6]), .op(n8616) );
  nand2_1 U10666 ( .ip1(n6791), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[5]), .op(n8619) );
  nor2_1 U10667 ( .ip1(n6791), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[5]), .op(n8636) );
  nand2_1 U10668 ( .ip1(n6815), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[4]), .op(n8617) );
  or2_1 U10669 ( .ip1(n8636), .ip2(n8617), .op(n8618) );
  nand2_1 U10670 ( .ip1(n5262), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[3]), .op(n8625) );
  nor2_1 U10671 ( .ip1(n5262), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[3]), .op(n8630) );
  nand2_1 U10672 ( .ip1(n8781), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[2]), .op(n8623) );
  or2_1 U10673 ( .ip1(n8630), .ip2(n8623), .op(n8624) );
  nand2_1 U10674 ( .ip1(n6802), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[1]), .op(n8629) );
  nor2_1 U10675 ( .ip1(n7943), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[0]), .op(n8627) );
  nor2_1 U10676 ( .ip1(n6802), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[1]), .op(n8626) );
  nor2_1 U10677 ( .ip1(n8781), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[2]), .op(n8631) );
  nor2_1 U10678 ( .ip1(n8631), .ip2(n8630), .op(n8632) );
  nor2_1 U10679 ( .ip1(n6815), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[4]), .op(n8637) );
  nor2_1 U10680 ( .ip1(n8637), .ip2(n8636), .op(n8639) );
  nand2_1 U10681 ( .ip1(n8639), .ip2(n8638), .op(n8640) );
  or2_1 U10682 ( .ip1(n8641), .ip2(n8640), .op(n8642) );
  nand2_1 U10683 ( .ip1(n8643), .ip2(n8642), .op(n8644) );
  and2_1 U10684 ( .ip1(n8645), .ip2(n8644), .op(n8646) );
  nor2_1 U10685 ( .ip1(n8647), .ip2(n8646), .op(n8648) );
  nand2_1 U10686 ( .ip1(n8801), .ip2(n8648), .op(n8722) );
  nand2_1 U10687 ( .ip1(n8880), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[15]), .op(n8651) );
  nand2_1 U10688 ( .ip1(n8881), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[14]), .op(n8649) );
  or2_1 U10689 ( .ip1(n8652), .ip2(n8649), .op(n8650) );
  nand2_1 U10690 ( .ip1(n8651), .ip2(n8650), .op(n8659) );
  nand2_1 U10691 ( .ip1(n8887), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[13]), .op(n8656) );
  nand2_1 U10692 ( .ip1(n8888), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[12]), .op(n8654) );
  or2_1 U10693 ( .ip1(n8660), .ip2(n8654), .op(n8655) );
  nand2_1 U10694 ( .ip1(n8656), .ip2(n8655), .op(n8657) );
  and2_1 U10695 ( .ip1(n8662), .ip2(n8657), .op(n8658) );
  nor2_1 U10696 ( .ip1(n8659), .ip2(n8658), .op(n8677) );
  nor2_1 U10697 ( .ip1(n8888), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[12]), .op(n8661) );
  nor2_1 U10698 ( .ip1(n8661), .ip2(n8660), .op(n8663) );
  nand2_1 U10699 ( .ip1(n8663), .ip2(n8662), .op(n8682) );
  nand2_1 U10700 ( .ip1(n8817), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[11]), .op(n8666) );
  nand2_1 U10701 ( .ip1(n8895), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[10]), .op(n8664) );
  or2_1 U10702 ( .ip1(n8667), .ip2(n8664), .op(n8665) );
  nand2_1 U10703 ( .ip1(n8666), .ip2(n8665), .op(n8674) );
  nand2_1 U10704 ( .ip1(n8897), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[9]), .op(n8671) );
  nand2_1 U10705 ( .ip1(n5461), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[8]), .op(n8669) );
  or2_1 U10706 ( .ip1(n8678), .ip2(n8669), .op(n8670) );
  nand2_1 U10707 ( .ip1(n8671), .ip2(n8670), .op(n8672) );
  and2_1 U10708 ( .ip1(n8680), .ip2(n8672), .op(n8673) );
  nor2_1 U10709 ( .ip1(n8674), .ip2(n8673), .op(n8675) );
  or2_1 U10710 ( .ip1(n8682), .ip2(n8675), .op(n8676) );
  nand2_1 U10711 ( .ip1(n8677), .ip2(n8676), .op(n8719) );
  nor2_1 U10712 ( .ip1(n5461), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[8]), .op(n8679) );
  nor2_1 U10713 ( .ip1(n8679), .ip2(n8678), .op(n8681) );
  nand2_1 U10714 ( .ip1(n8681), .ip2(n8680), .op(n8683) );
  nor2_1 U10715 ( .ip1(n8683), .ip2(n8682), .op(n8717) );
  nand2_1 U10716 ( .ip1(n8133), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[7]), .op(n8686) );
  nand2_1 U10717 ( .ip1(n8922), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[6]), .op(n8684) );
  or2_1 U10718 ( .ip1(n8687), .ip2(n8684), .op(n8685) );
  nand2_1 U10719 ( .ip1(n8686), .ip2(n8685), .op(n8694) );
  nor2_1 U10720 ( .ip1(n8922), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[6]), .op(n8688) );
  nand2_1 U10721 ( .ip1(n8928), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[5]), .op(n8691) );
  nor2_1 U10722 ( .ip1(n8928), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[5]), .op(n8708) );
  nand2_1 U10723 ( .ip1(n5467), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[4]), .op(n8689) );
  or2_1 U10724 ( .ip1(n8708), .ip2(n8689), .op(n8690) );
  nand2_1 U10725 ( .ip1(n8691), .ip2(n8690), .op(n8692) );
  and2_1 U10726 ( .ip1(n8710), .ip2(n8692), .op(n8693) );
  nor2_1 U10727 ( .ip1(n8694), .ip2(n8693), .op(n8715) );
  nand2_1 U10728 ( .ip1(n5465), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[3]), .op(n8697) );
  nor2_1 U10729 ( .ip1(n5465), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[3]), .op(n8702) );
  nand2_1 U10730 ( .ip1(n8935), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[2]), .op(n8695) );
  or2_1 U10731 ( .ip1(n8702), .ip2(n8695), .op(n8696) );
  nand2_1 U10732 ( .ip1(n8697), .ip2(n8696), .op(n8707) );
  nand2_1 U10733 ( .ip1(n8939), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[1]), .op(n8701) );
  nor2_1 U10734 ( .ip1(n8940), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[0]), .op(n8699) );
  nor2_1 U10735 ( .ip1(n8939), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[1]), .op(n8698) );
  or2_1 U10736 ( .ip1(n8699), .ip2(n8698), .op(n8700) );
  nand2_1 U10737 ( .ip1(n8701), .ip2(n8700), .op(n8705) );
  nor2_1 U10738 ( .ip1(n8935), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[2]), .op(n8703) );
  nor2_1 U10739 ( .ip1(n8703), .ip2(n8702), .op(n8704) );
  and2_1 U10740 ( .ip1(n8705), .ip2(n8704), .op(n8706) );
  nor2_1 U10741 ( .ip1(n8707), .ip2(n8706), .op(n8713) );
  nor2_1 U10742 ( .ip1(n5467), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[4]), .op(n8709) );
  nor2_1 U10743 ( .ip1(n8709), .ip2(n8708), .op(n8711) );
  nand2_1 U10744 ( .ip1(n8711), .ip2(n8710), .op(n8712) );
  or2_1 U10745 ( .ip1(n8713), .ip2(n8712), .op(n8714) );
  nand2_1 U10746 ( .ip1(n8715), .ip2(n8714), .op(n8716) );
  and2_1 U10747 ( .ip1(n8717), .ip2(n8716), .op(n8718) );
  nor2_1 U10748 ( .ip1(n8719), .ip2(n8718), .op(n8720) );
  nand2_1 U10749 ( .ip1(n8720), .ip2(n8874), .op(n8721) );
  inv_1 U10750 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[4]), .op(
        n10647) );
  inv_1 U10751 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[6]), .op(
        n10653) );
  inv_1 U10752 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[8]), .op(
        n10659) );
  inv_1 U10753 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[10]), .op(
        n10665) );
  inv_1 U10754 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[12]), .op(
        n10671) );
  inv_1 U10755 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[14]), .op(
        n10679) );
  nor2_1 U10756 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_re_scl_s_hld_en), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_st_scl_s_hld_en), .op(n11041) );
  and3_1 U10757 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[2]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[0]), .ip3(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[1]), .op(n8878) );
  nand2_1 U10758 ( .ip1(n6727), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[15]), .op(n8727) );
  nor2_1 U10759 ( .ip1(n6727), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[15]), .op(n8728) );
  nand2_1 U10760 ( .ip1(n6734), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[14]), .op(n8725) );
  or2_1 U10761 ( .ip1(n8728), .ip2(n8725), .op(n8726) );
  nand2_1 U10762 ( .ip1(n8727), .ip2(n8726), .op(n8736) );
  nor2_1 U10763 ( .ip1(n6734), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[14]), .op(n8729) );
  nor2_1 U10764 ( .ip1(n8729), .ip2(n8728), .op(n8739) );
  nand2_1 U10765 ( .ip1(n8730), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[13]), .op(n8733) );
  nor2_1 U10766 ( .ip1(n8730), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[13]), .op(n8737) );
  nand2_1 U10767 ( .ip1(n6744), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[12]), .op(n8731) );
  or2_1 U10768 ( .ip1(n8737), .ip2(n8731), .op(n8732) );
  nand2_1 U10769 ( .ip1(n8733), .ip2(n8732), .op(n8734) );
  and2_1 U10770 ( .ip1(n8739), .ip2(n8734), .op(n8735) );
  nor2_1 U10771 ( .ip1(n6744), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[12]), .op(n8738) );
  nor2_1 U10772 ( .ip1(n8738), .ip2(n8737), .op(n8740) );
  nand2_1 U10773 ( .ip1(n8740), .ip2(n8739), .op(n8760) );
  nand2_1 U10774 ( .ip1(n8741), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[11]), .op(n8744) );
  nor2_1 U10775 ( .ip1(n8741), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[11]), .op(n8745) );
  nand2_1 U10776 ( .ip1(n6760), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[10]), .op(n8742) );
  or2_1 U10777 ( .ip1(n8745), .ip2(n8742), .op(n8743) );
  nand2_1 U10778 ( .ip1(n8744), .ip2(n8743), .op(n8752) );
  nor2_1 U10779 ( .ip1(n6760), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[10]), .op(n8746) );
  nor2_1 U10780 ( .ip1(n8746), .ip2(n8745), .op(n8758) );
  nand2_1 U10781 ( .ip1(n6772), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[9]), .op(n8749) );
  nor2_1 U10782 ( .ip1(n6772), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[9]), .op(n8756) );
  nand2_1 U10783 ( .ip1(n5272), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[8]), .op(n8747) );
  or2_1 U10784 ( .ip1(n8756), .ip2(n8747), .op(n8748) );
  and2_1 U10785 ( .ip1(n8758), .ip2(n8750), .op(n8751) );
  nor2_1 U10786 ( .ip1(n8752), .ip2(n8751), .op(n8753) );
  or2_1 U10787 ( .ip1(n8760), .ip2(n8753), .op(n8754) );
  nand2_1 U10788 ( .ip1(n8755), .ip2(n8754), .op(n8799) );
  nor2_1 U10789 ( .ip1(n5272), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[8]), .op(n8757) );
  nor2_1 U10790 ( .ip1(n8757), .ip2(n8756), .op(n8759) );
  nand2_1 U10791 ( .ip1(n8759), .ip2(n8758), .op(n8761) );
  nor2_1 U10792 ( .ip1(n8761), .ip2(n8760), .op(n8797) );
  nand2_1 U10793 ( .ip1(n8762), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[7]), .op(n8765) );
  nor2_1 U10794 ( .ip1(n8762), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[7]), .op(n8766) );
  nand2_1 U10795 ( .ip1(n6784), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[6]), .op(n8763) );
  or2_1 U10796 ( .ip1(n8766), .ip2(n8763), .op(n8764) );
  nor2_1 U10797 ( .ip1(n6784), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[6]), .op(n8767) );
  nand2_1 U10798 ( .ip1(n6791), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[5]), .op(n8770) );
  nor2_1 U10799 ( .ip1(n6791), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[5]), .op(n8788) );
  nand2_1 U10800 ( .ip1(n6815), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[4]), .op(n8768) );
  or2_1 U10801 ( .ip1(n8788), .ip2(n8768), .op(n8769) );
  nand2_1 U10802 ( .ip1(n5262), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[3]), .op(n8776) );
  nor2_1 U10803 ( .ip1(n5262), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[3]), .op(n8782) );
  nand2_1 U10804 ( .ip1(n8781), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[2]), .op(n8774) );
  or2_1 U10805 ( .ip1(n8782), .ip2(n8774), .op(n8775) );
  nand2_1 U10806 ( .ip1(n6802), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[1]), .op(n8780) );
  nor2_1 U10807 ( .ip1(n7943), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[0]), .op(n8778) );
  nor2_1 U10808 ( .ip1(n6802), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[1]), .op(n8777) );
  nor2_1 U10809 ( .ip1(n8781), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[2]), .op(n8783) );
  nor2_1 U10810 ( .ip1(n8783), .ip2(n8782), .op(n8784) );
  nor2_1 U10811 ( .ip1(n6815), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[4]), .op(n8789) );
  nor2_1 U10812 ( .ip1(n8789), .ip2(n8788), .op(n8791) );
  nand2_1 U10813 ( .ip1(n8791), .ip2(n8790), .op(n8792) );
  or2_1 U10814 ( .ip1(n8793), .ip2(n8792), .op(n8794) );
  nand2_1 U10815 ( .ip1(n8795), .ip2(n8794), .op(n8796) );
  and2_1 U10816 ( .ip1(n8797), .ip2(n8796), .op(n8798) );
  nor2_1 U10817 ( .ip1(n8799), .ip2(n8798), .op(n8800) );
  nand2_1 U10818 ( .ip1(n8801), .ip2(n8800), .op(n8877) );
  nand2_1 U10819 ( .ip1(n8880), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[15]), .op(n8804) );
  nand2_1 U10820 ( .ip1(n8881), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[14]), .op(n8802) );
  or2_1 U10821 ( .ip1(n8805), .ip2(n8802), .op(n8803) );
  nand2_1 U10822 ( .ip1(n8804), .ip2(n8803), .op(n8812) );
  nand2_1 U10823 ( .ip1(n8887), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[13]), .op(n8809) );
  nand2_1 U10824 ( .ip1(n8888), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[12]), .op(n8807) );
  or2_1 U10825 ( .ip1(n8813), .ip2(n8807), .op(n8808) );
  nand2_1 U10826 ( .ip1(n8809), .ip2(n8808), .op(n8810) );
  and2_1 U10827 ( .ip1(n8815), .ip2(n8810), .op(n8811) );
  nor2_1 U10828 ( .ip1(n8812), .ip2(n8811), .op(n8831) );
  nor2_1 U10829 ( .ip1(n8888), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[12]), .op(n8814) );
  nor2_1 U10830 ( .ip1(n8814), .ip2(n8813), .op(n8816) );
  nand2_1 U10831 ( .ip1(n8816), .ip2(n8815), .op(n8836) );
  nand2_1 U10832 ( .ip1(n8817), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[11]), .op(n8820) );
  nand2_1 U10833 ( .ip1(n8895), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[10]), .op(n8818) );
  or2_1 U10834 ( .ip1(n8821), .ip2(n8818), .op(n8819) );
  nand2_1 U10835 ( .ip1(n8820), .ip2(n8819), .op(n8828) );
  nand2_1 U10836 ( .ip1(n8897), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[9]), .op(n8825) );
  nand2_1 U10837 ( .ip1(n5461), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[8]), .op(n8823) );
  or2_1 U10838 ( .ip1(n8832), .ip2(n8823), .op(n8824) );
  nand2_1 U10839 ( .ip1(n8825), .ip2(n8824), .op(n8826) );
  and2_1 U10840 ( .ip1(n8834), .ip2(n8826), .op(n8827) );
  nor2_1 U10841 ( .ip1(n8828), .ip2(n8827), .op(n8829) );
  or2_1 U10842 ( .ip1(n8836), .ip2(n8829), .op(n8830) );
  nand2_1 U10843 ( .ip1(n8831), .ip2(n8830), .op(n8873) );
  nor2_1 U10844 ( .ip1(n5461), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[8]), .op(n8833) );
  nor2_1 U10845 ( .ip1(n8833), .ip2(n8832), .op(n8835) );
  nand2_1 U10846 ( .ip1(n8835), .ip2(n8834), .op(n8837) );
  nor2_1 U10847 ( .ip1(n8837), .ip2(n8836), .op(n8871) );
  nand2_1 U10848 ( .ip1(n8133), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[7]), .op(n8840) );
  nand2_1 U10849 ( .ip1(n8922), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[6]), .op(n8838) );
  or2_1 U10850 ( .ip1(n8841), .ip2(n8838), .op(n8839) );
  nand2_1 U10851 ( .ip1(n8840), .ip2(n8839), .op(n8848) );
  nor2_1 U10852 ( .ip1(n8922), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[6]), .op(n8842) );
  nand2_1 U10853 ( .ip1(n8928), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[5]), .op(n8845) );
  nor2_1 U10854 ( .ip1(n8928), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[5]), .op(n8862) );
  nand2_1 U10855 ( .ip1(n5467), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[4]), .op(n8843) );
  or2_1 U10856 ( .ip1(n8862), .ip2(n8843), .op(n8844) );
  nand2_1 U10857 ( .ip1(n8845), .ip2(n8844), .op(n8846) );
  and2_1 U10858 ( .ip1(n8864), .ip2(n8846), .op(n8847) );
  nor2_1 U10859 ( .ip1(n8848), .ip2(n8847), .op(n8869) );
  nand2_1 U10860 ( .ip1(n5465), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[3]), .op(n8851) );
  nor2_1 U10861 ( .ip1(n5465), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[3]), .op(n8856) );
  nand2_1 U10862 ( .ip1(n8935), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[2]), .op(n8849) );
  or2_1 U10863 ( .ip1(n8856), .ip2(n8849), .op(n8850) );
  nand2_1 U10864 ( .ip1(n8851), .ip2(n8850), .op(n8861) );
  nand2_1 U10865 ( .ip1(n8939), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[1]), .op(n8855) );
  nor2_1 U10866 ( .ip1(n8940), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[0]), .op(n8853) );
  nor2_1 U10867 ( .ip1(n8939), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[1]), .op(n8852) );
  or2_1 U10868 ( .ip1(n8853), .ip2(n8852), .op(n8854) );
  nand2_1 U10869 ( .ip1(n8855), .ip2(n8854), .op(n8859) );
  nor2_1 U10870 ( .ip1(n8935), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[2]), .op(n8857) );
  nor2_1 U10871 ( .ip1(n8857), .ip2(n8856), .op(n8858) );
  and2_1 U10872 ( .ip1(n8859), .ip2(n8858), .op(n8860) );
  nor2_1 U10873 ( .ip1(n8861), .ip2(n8860), .op(n8867) );
  nor2_1 U10874 ( .ip1(n5467), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[4]), .op(n8863) );
  nor2_1 U10875 ( .ip1(n8863), .ip2(n8862), .op(n8865) );
  nand2_1 U10876 ( .ip1(n8865), .ip2(n8864), .op(n8866) );
  or2_1 U10877 ( .ip1(n8867), .ip2(n8866), .op(n8868) );
  nand2_1 U10878 ( .ip1(n8869), .ip2(n8868), .op(n8870) );
  and2_1 U10879 ( .ip1(n8871), .ip2(n8870), .op(n8872) );
  nor2_1 U10880 ( .ip1(n8873), .ip2(n8872), .op(n8875) );
  nand2_1 U10881 ( .ip1(n8875), .ip2(n8874), .op(n8876) );
  inv_1 U10882 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[4]), .op(n11010) );
  inv_1 U10883 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[6]), .op(n11016) );
  inv_1 U10884 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[8]), .op(n11022) );
  inv_1 U10885 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[10]), .op(
        n11028) );
  inv_1 U10886 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[12]), .op(
        n11034) );
  inv_1 U10887 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[14]), .op(
        n11042) );
  inv_1 U10888 ( .ip(i_i2c_scl_s_setup_en), .op(n10994) );
  nand2_1 U10889 ( .ip1(n8880), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[15]), .op(n8884) );
  nand2_1 U10890 ( .ip1(n8881), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[14]), .op(n8882) );
  or2_1 U10891 ( .ip1(n8885), .ip2(n8882), .op(n8883) );
  nand2_1 U10892 ( .ip1(n8884), .ip2(n8883), .op(n8894) );
  nand2_1 U10893 ( .ip1(n8887), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[13]), .op(n8891) );
  nand2_1 U10894 ( .ip1(n8888), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[12]), .op(n8889) );
  or2_1 U10895 ( .ip1(n8907), .ip2(n8889), .op(n8890) );
  nand2_1 U10896 ( .ip1(n8891), .ip2(n8890), .op(n8892) );
  and2_1 U10897 ( .ip1(n8909), .ip2(n8892), .op(n8893) );
  nor2_1 U10898 ( .ip1(n8894), .ip2(n8893), .op(n8914) );
  nor2_1 U10899 ( .ip1(n8817), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[11]), .op(n8903) );
  nor2_1 U10900 ( .ip1(n8895), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[10]), .op(n8896) );
  nand2_1 U10901 ( .ip1(n8897), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[9]), .op(n8900) );
  nand2_1 U10902 ( .ip1(n5461), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[8]), .op(n8898) );
  or2_1 U10903 ( .ip1(n8915), .ip2(n8898), .op(n8899) );
  nand2_1 U10904 ( .ip1(n8900), .ip2(n8899), .op(n8901) );
  nand2_1 U10905 ( .ip1(n8817), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[11]), .op(n8905) );
  nand2_1 U10906 ( .ip1(n8895), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[10]), .op(n8902) );
  or2_1 U10907 ( .ip1(n8903), .ip2(n8902), .op(n8904) );
  nor2_1 U10908 ( .ip1(n8888), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[12]), .op(n8908) );
  nor2_1 U10909 ( .ip1(n8908), .ip2(n8907), .op(n8910) );
  nand2_1 U10910 ( .ip1(n8910), .ip2(n8909), .op(n8919) );
  nand2_1 U10911 ( .ip1(n8914), .ip2(n8913), .op(n8961) );
  nor2_1 U10912 ( .ip1(n5461), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[8]), .op(n8916) );
  nor2_1 U10913 ( .ip1(n8916), .ip2(n8915), .op(n8918) );
  nand2_1 U10914 ( .ip1(n8918), .ip2(n8917), .op(n8920) );
  nor2_1 U10915 ( .ip1(n8920), .ip2(n8919), .op(n8959) );
  nand2_1 U10916 ( .ip1(n8133), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[7]), .op(n8925) );
  nor2_1 U10917 ( .ip1(n8133), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[7]), .op(n8926) );
  nand2_1 U10918 ( .ip1(n8922), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[6]), .op(n8923) );
  or2_1 U10919 ( .ip1(n8926), .ip2(n8923), .op(n8924) );
  nand2_1 U10920 ( .ip1(n8925), .ip2(n8924), .op(n8934) );
  nor2_1 U10921 ( .ip1(n8922), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[6]), .op(n8927) );
  nor2_1 U10922 ( .ip1(n8927), .ip2(n8926), .op(n8952) );
  nand2_1 U10923 ( .ip1(n8928), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[5]), .op(n8931) );
  nor2_1 U10924 ( .ip1(n8928), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[5]), .op(n8950) );
  nand2_1 U10925 ( .ip1(n5467), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[4]), .op(n8929) );
  or2_1 U10926 ( .ip1(n8950), .ip2(n8929), .op(n8930) );
  nand2_1 U10927 ( .ip1(n8931), .ip2(n8930), .op(n8932) );
  and2_1 U10928 ( .ip1(n8952), .ip2(n8932), .op(n8933) );
  nor2_1 U10929 ( .ip1(n8934), .ip2(n8933), .op(n8957) );
  nand2_1 U10930 ( .ip1(n5465), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[3]), .op(n8938) );
  nor2_1 U10931 ( .ip1(n5465), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[3]), .op(n8944) );
  nand2_1 U10932 ( .ip1(n8935), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[2]), .op(n8936) );
  or2_1 U10933 ( .ip1(n8944), .ip2(n8936), .op(n8937) );
  nand2_1 U10934 ( .ip1(n8939), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[1]), .op(n8943) );
  nor2_1 U10935 ( .ip1(n8939), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[1]), .op(n8941) );
  nor2_1 U10936 ( .ip1(n8935), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[2]), .op(n8945) );
  nor2_1 U10937 ( .ip1(n8945), .ip2(n8944), .op(n8946) );
  and2_1 U10938 ( .ip1(n8947), .ip2(n8946), .op(n8948) );
  nor2_1 U10939 ( .ip1(n5467), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[4]), .op(n8951) );
  nor2_1 U10940 ( .ip1(n8951), .ip2(n8950), .op(n8953) );
  nand2_1 U10941 ( .ip1(n8953), .ip2(n8952), .op(n8954) );
  or2_1 U10942 ( .ip1(n8955), .ip2(n8954), .op(n8956) );
  nand2_1 U10943 ( .ip1(n8957), .ip2(n8956), .op(n8958) );
  and2_1 U10944 ( .ip1(n8959), .ip2(n8958), .op(n8960) );
  nor2_1 U10945 ( .ip1(n8961), .ip2(n8960), .op(n8964) );
  nand2_1 U10946 ( .ip1(n8964), .ip2(n8963), .op(n9052) );
  inv_1 U10947 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[15]), .op(
        n8965) );
  nand2_1 U10948 ( .ip1(n8966), .ip2(n8965), .op(n9048) );
  nor2_1 U10949 ( .ip1(n8966), .ip2(n8965), .op(n9046) );
  inv_1 U10950 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[14]), .op(
        n9054) );
  and2_1 U10951 ( .ip1(n8967), .ip2(n9054), .op(n9044) );
  nor2_1 U10952 ( .ip1(n8967), .ip2(n9054), .op(n9042) );
  inv_1 U10953 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[13]), .op(
        n8968) );
  nand2_1 U10954 ( .ip1(n8969), .ip2(n8968), .op(n9040) );
  nor2_1 U10955 ( .ip1(n8969), .ip2(n8968), .op(n9038) );
  inv_1 U10956 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[12]), .op(
        n10991) );
  nand2_1 U10957 ( .ip1(n8970), .ip2(n10991), .op(n8973) );
  inv_1 U10958 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[11]), .op(
        n9029) );
  nand2_1 U10959 ( .ip1(n9030), .ip2(n9029), .op(n8971) );
  nor2_1 U10960 ( .ip1(n8970), .ip2(n10991), .op(n9032) );
  or2_1 U10961 ( .ip1(n8971), .ip2(n9032), .op(n8972) );
  nand2_1 U10962 ( .ip1(n8973), .ip2(n8972), .op(n9036) );
  inv_1 U10963 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[8]), .op(
        n9021) );
  inv_1 U10964 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[7]), .op(
        n10979) );
  nor2_1 U10965 ( .ip1(n9018), .ip2(n10979), .op(n8974) );
  nor2_1 U10966 ( .ip1(n9019), .ip2(n8974), .op(n8976) );
  inv_1 U10967 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[9]), .op(
        n9012) );
  nor2_1 U10968 ( .ip1(n9013), .ip2(n9012), .op(n8975) );
  inv_1 U10969 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[10]), .op(
        n9010) );
  nor2_1 U10970 ( .ip1(n9011), .ip2(n9010), .op(n9014) );
  nor2_1 U10971 ( .ip1(n8975), .ip2(n9014), .op(n9025) );
  nand2_1 U10972 ( .ip1(n8976), .ip2(n9025), .op(n9009) );
  inv_1 U10973 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[6]), .op(
        n10977) );
  nor2_1 U10974 ( .ip1(n8977), .ip2(n10977), .op(n8981) );
  inv_1 U10975 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[5]), .op(
        n10973) );
  nand2_1 U10976 ( .ip1(n8980), .ip2(n10973), .op(n8978) );
  nor2_1 U10977 ( .ip1(n8981), .ip2(n8978), .op(n8979) );
  inv_1 U10978 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[4]), .op(
        n10971) );
  nand2_1 U10979 ( .ip1(n9001), .ip2(n10971), .op(n8984) );
  or2_1 U10980 ( .ip1(n8980), .ip2(n10973), .op(n8983) );
  inv_1 U10981 ( .ip(n8981), .op(n8982) );
  or2_1 U10982 ( .ip1(n8984), .ip2(n9003), .op(n8985) );
  inv_1 U10983 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[3]), .op(
        n9950) );
  nand2_1 U10984 ( .ip1(n6800), .ip2(n9950), .op(n9000) );
  inv_1 U10985 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[2]), .op(
        n10968) );
  inv_1 U10986 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[1]), .op(
        n10964) );
  inv_1 U10987 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[0]), .op(
        n10959) );
  or2_1 U10988 ( .ip1(n6800), .ip2(n9950), .op(n8997) );
  nor2_1 U10989 ( .ip1(n9001), .ip2(n10971), .op(n9002) );
  or2_1 U10990 ( .ip1(n9009), .ip2(n9008), .op(n9028) );
  nand2_1 U10991 ( .ip1(n9011), .ip2(n9010), .op(n9017) );
  nand2_1 U10992 ( .ip1(n9013), .ip2(n9012), .op(n9015) );
  or2_1 U10993 ( .ip1(n9015), .ip2(n9014), .op(n9016) );
  nand2_1 U10994 ( .ip1(n9018), .ip2(n10979), .op(n9020) );
  or2_1 U10995 ( .ip1(n9020), .ip2(n9019), .op(n9024) );
  nand2_1 U10996 ( .ip1(n9022), .ip2(n9021), .op(n9023) );
  nor2_1 U10997 ( .ip1(n9030), .ip2(n9029), .op(n9031) );
  nor2_1 U10998 ( .ip1(n9032), .ip2(n9031), .op(n9033) );
  and2_1 U10999 ( .ip1(n9034), .ip2(n9033), .op(n9035) );
  nor2_1 U11000 ( .ip1(n9036), .ip2(n9035), .op(n9037) );
  or2_1 U11001 ( .ip1(n9038), .ip2(n9037), .op(n9039) );
  nor2_1 U11002 ( .ip1(n9042), .ip2(n9041), .op(n9043) );
  nor2_1 U11003 ( .ip1(n9044), .ip2(n9043), .op(n9045) );
  or2_1 U11004 ( .ip1(n9046), .ip2(n9045), .op(n9047) );
  nand2_1 U11005 ( .ip1(n9048), .ip2(n9047), .op(n9050) );
  nand2_1 U11006 ( .ip1(n11170), .ip2(n10719), .op(n9049) );
  nand2_1 U11007 ( .ip1(n9050), .ip2(n9049), .op(n9051) );
  and3_1 U11008 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[2]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[0]), .ip3(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[1]), .op(n9949) );
  and2_1 U11009 ( .ip1(n10990), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[12]), .op(n10993) );
  inv_1 U11010 ( .ip(i_ssi_ssi_rst_n), .op(n11764) );
  inv_1 U11011 ( .ip(i_i2c_ic_hs), .op(n11763) );
  nor2_1 U11012 ( .ip1(n11702), .ip2(i_ssi_U_mstfsm_ctrl_cnt[0]), .op(n9064)
         );
  nand2_1 U11013 ( .ip1(n11702), .ip2(i_ssi_U_mstfsm_ctrl_cnt[0]), .op(n11705)
         );
  inv_1 U11014 ( .ip(n11705), .op(n9063) );
  nor2_1 U11015 ( .ip1(n5481), .ip2(n9056), .op(n9687) );
  nand2_1 U11016 ( .ip1(n9687), .ip2(n9057), .op(n9062) );
  nor3_1 U11017 ( .ip1(i_ssi_U_mstfsm_c_state[3]), .ip2(
        i_ssi_U_mstfsm_c_state[1]), .ip3(n9058), .op(n9060) );
  nand2_1 U11018 ( .ip1(n9060), .ip2(n9059), .op(n9061) );
  nand2_1 U11019 ( .ip1(n9062), .ip2(n9061), .op(n11708) );
  nor3_1 U11020 ( .ip1(n9064), .ip2(n9063), .ip3(n11708), .op(n4205) );
  mux2_1 U11021 ( .ip1(n9066), .ip2(n9065), .s(n11718), .op(n9067) );
  inv_1 U11022 ( .ip(n9067), .op(n5082) );
  inv_1 U11023 ( .ip(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[13]), .op(n9069) );
  inv_1 U11024 ( .ip(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[12]), .op(n9068) );
  nor3_1 U11025 ( .ip1(n9069), .ip2(n9070), .ip3(n9068), .op(
        ex_i_ahb_AHB_Slave_PID_hsel) );
  nor3_1 U11026 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[12]), .ip2(n9070), 
        .ip3(n9069), .op(ex_i_ahb_AHB_Slave_PWM_hsel) );
  inv_1 U11027 ( .ip(n9071), .op(n9072) );
  nand2_1 U11028 ( .ip1(n9074), .ip2(n9073), .op(n9075) );
  xor2_1 U11029 ( .ip1(i_ssi_U_fifo_unconnected_tx_wrd_count[2]), .ip2(n9075), 
        .op(n9076) );
  nor2_4 U11030 ( .ip1(n11227), .ip2(n9076), .op(n11779) );
  nand4_1 U11031 ( .ip1(i_ssi_U_fifo_unconnected_rx_wrd_count[2]), .ip2(n11760), .ip3(i_ssi_U_fifo_unconnected_rx_wrd_count[0]), .ip4(
        i_ssi_U_fifo_unconnected_rx_wrd_count[1]), .op(n9077) );
  nand2_1 U11032 ( .ip1(n11165), .ip2(n9078), .op(n9079) );
  nand2_1 U11033 ( .ip1(n11760), .ip2(i_ssi_rx_full), .op(n11166) );
  nor2_1 U11034 ( .ip1(n9080), .ip2(n11227), .op(n11777) );
  xor2_1 U11035 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[13]), .ip2(
        n10244), .op(n9081) );
  nor2_4 U11036 ( .ip1(n10275), .ip2(n9081), .op(n4152) );
  and2_1 U11037 ( .ip1(i_ssi_U_mstfsm_frame_cnt[15]), .ip2(
        i_ssi_U_mstfsm_frame_cnt[14]), .op(n10541) );
  nand3_1 U11038 ( .ip1(n9086), .ip2(n5480), .ip3(n9085), .op(n9087) );
  inv_1 U11039 ( .ip(n10385), .op(n10293) );
  nor4_1 U11040 ( .ip1(i_ssi_baudr[12]), .ip2(n5257), .ip3(n10384), .ip4(
        i_ssi_baudr[15]), .op(n9090) );
  nand3_1 U11041 ( .ip1(n9090), .ip2(n9089), .ip3(n9088), .op(n9091) );
  inv_1 U11042 ( .ip(n10294), .op(n9094) );
  nor2_1 U11043 ( .ip1(n10293), .ip2(n9094), .op(n5241) );
  inv_1 U11044 ( .ip(n9095), .op(n11282) );
  nor2_1 U11045 ( .ip1(n11282), .ip2(n9096), .op(n9097) );
  xor2_1 U11046 ( .ip1(i_i2c_tx_abrt_source[15]), .ip2(n9097), .op(n5118) );
  inv_1 U11047 ( .ip(i_i2c_rx_rd_addr[1]), .op(n11186) );
  nor3_1 U11048 ( .ip1(i_i2c_rx_rd_addr[2]), .ip2(i_i2c_rx_rd_addr[0]), .ip3(
        n11186), .op(n9167) );
  nand2_1 U11049 ( .ip1(n9167), .ip2(i_i2c_U_dff_rx_mem[40]), .op(n9107) );
  nand2_1 U11050 ( .ip1(i_i2c_rx_rd_addr[0]), .ip2(i_i2c_rx_rd_addr[1]), .op(
        n11183) );
  nor2_1 U11051 ( .ip1(i_i2c_rx_rd_addr[2]), .ip2(n11183), .op(n9169) );
  inv_1 U11052 ( .ip(i_i2c_rx_rd_addr[2]), .op(n9098) );
  inv_1 U11053 ( .ip(i_i2c_rx_rd_addr[0]), .op(n11203) );
  nor3_1 U11054 ( .ip1(n9098), .ip2(n11203), .ip3(n11186), .op(n11190) );
  and2_1 U11055 ( .ip1(i_i2c_U_dff_rx_mem[0]), .ip2(n11190), .op(n9104) );
  nor3_1 U11056 ( .ip1(i_i2c_rx_rd_addr[0]), .ip2(n9098), .ip3(n11186), .op(
        n9177) );
  nand2_1 U11057 ( .ip1(i_i2c_U_dff_rx_mem[8]), .ip2(n9177), .op(n9102) );
  nor3_1 U11058 ( .ip1(i_i2c_rx_rd_addr[0]), .ip2(i_i2c_rx_rd_addr[1]), .ip3(
        n9098), .op(n9166) );
  nand2_1 U11059 ( .ip1(i_i2c_U_dff_rx_mem[24]), .ip2(n9166), .op(n9101) );
  nor3_1 U11060 ( .ip1(i_i2c_rx_rd_addr[2]), .ip2(i_i2c_rx_rd_addr[0]), .ip3(
        i_i2c_rx_rd_addr[1]), .op(n9168) );
  nand2_1 U11061 ( .ip1(i_i2c_U_dff_rx_mem[56]), .ip2(n9168), .op(n9100) );
  nor3_1 U11062 ( .ip1(i_i2c_rx_rd_addr[1]), .ip2(n11203), .ip3(n9098), .op(
        n9170) );
  nand2_1 U11063 ( .ip1(i_i2c_U_dff_rx_mem[16]), .ip2(n9170), .op(n9099) );
  nand4_1 U11064 ( .ip1(n9102), .ip2(n9101), .ip3(n9100), .ip4(n9099), .op(
        n9103) );
  not_ab_or_c_or_d U11065 ( .ip1(i_i2c_U_dff_rx_mem[32]), .ip2(n9169), .ip3(
        n9104), .ip4(n9103), .op(n9106) );
  nor3_1 U11066 ( .ip1(i_i2c_rx_rd_addr[2]), .ip2(i_i2c_rx_rd_addr[1]), .ip3(
        n11203), .op(n9178) );
  nand2_1 U11067 ( .ip1(i_i2c_U_dff_rx_mem[48]), .ip2(n9178), .op(n9105) );
  nand3_1 U11068 ( .ip1(n9107), .ip2(n9106), .ip3(n9105), .op(
        i_i2c_rx_pop_data[0]) );
  nand2_1 U11069 ( .ip1(i_i2c_U_dff_rx_mem[23]), .ip2(n9170), .op(n9116) );
  and2_1 U11070 ( .ip1(i_i2c_U_dff_rx_mem[7]), .ip2(n11190), .op(n9113) );
  nand2_1 U11071 ( .ip1(i_i2c_U_dff_rx_mem[47]), .ip2(n9167), .op(n9111) );
  nand2_1 U11072 ( .ip1(i_i2c_U_dff_rx_mem[55]), .ip2(n9178), .op(n9110) );
  nand2_1 U11073 ( .ip1(i_i2c_U_dff_rx_mem[15]), .ip2(n9177), .op(n9109) );
  nand2_1 U11074 ( .ip1(i_i2c_U_dff_rx_mem[39]), .ip2(n9169), .op(n9108) );
  nand4_1 U11075 ( .ip1(n9111), .ip2(n9110), .ip3(n9109), .ip4(n9108), .op(
        n9112) );
  not_ab_or_c_or_d U11076 ( .ip1(n9168), .ip2(i_i2c_U_dff_rx_mem[63]), .ip3(
        n9113), .ip4(n9112), .op(n9115) );
  nand2_1 U11077 ( .ip1(i_i2c_U_dff_rx_mem[31]), .ip2(n9166), .op(n9114) );
  nand3_1 U11078 ( .ip1(n9116), .ip2(n9115), .ip3(n9114), .op(
        i_i2c_rx_pop_data[7]) );
  nand2_1 U11079 ( .ip1(i_i2c_U_dff_rx_mem[20]), .ip2(n9170), .op(n9125) );
  and2_1 U11080 ( .ip1(i_i2c_U_dff_rx_mem[4]), .ip2(n11190), .op(n9122) );
  nand2_1 U11081 ( .ip1(i_i2c_U_dff_rx_mem[28]), .ip2(n9166), .op(n9120) );
  nand2_1 U11082 ( .ip1(i_i2c_U_dff_rx_mem[60]), .ip2(n9168), .op(n9119) );
  nand2_1 U11083 ( .ip1(i_i2c_U_dff_rx_mem[52]), .ip2(n9178), .op(n9118) );
  nand2_1 U11084 ( .ip1(i_i2c_U_dff_rx_mem[12]), .ip2(n9177), .op(n9117) );
  nand4_1 U11085 ( .ip1(n9120), .ip2(n9119), .ip3(n9118), .ip4(n9117), .op(
        n9121) );
  not_ab_or_c_or_d U11086 ( .ip1(n9169), .ip2(i_i2c_U_dff_rx_mem[36]), .ip3(
        n9122), .ip4(n9121), .op(n9124) );
  nand2_1 U11087 ( .ip1(i_i2c_U_dff_rx_mem[44]), .ip2(n9167), .op(n9123) );
  nand3_1 U11088 ( .ip1(n9125), .ip2(n9124), .ip3(n9123), .op(
        i_i2c_rx_pop_data[4]) );
  nand2_1 U11089 ( .ip1(i_i2c_U_dff_rx_mem[21]), .ip2(n9170), .op(n9134) );
  and2_1 U11090 ( .ip1(i_i2c_U_dff_rx_mem[5]), .ip2(n11190), .op(n9131) );
  nand2_1 U11091 ( .ip1(i_i2c_U_dff_rx_mem[29]), .ip2(n9166), .op(n9129) );
  nand2_1 U11092 ( .ip1(i_i2c_U_dff_rx_mem[61]), .ip2(n9168), .op(n9128) );
  nand2_1 U11093 ( .ip1(i_i2c_U_dff_rx_mem[13]), .ip2(n9177), .op(n9127) );
  nand2_1 U11094 ( .ip1(i_i2c_U_dff_rx_mem[37]), .ip2(n9169), .op(n9126) );
  nand4_1 U11095 ( .ip1(n9129), .ip2(n9128), .ip3(n9127), .ip4(n9126), .op(
        n9130) );
  not_ab_or_c_or_d U11096 ( .ip1(n9167), .ip2(i_i2c_U_dff_rx_mem[45]), .ip3(
        n9131), .ip4(n9130), .op(n9133) );
  nand2_1 U11097 ( .ip1(i_i2c_U_dff_rx_mem[53]), .ip2(n9178), .op(n9132) );
  nand3_1 U11098 ( .ip1(n9134), .ip2(n9133), .ip3(n9132), .op(
        i_i2c_rx_pop_data[5]) );
  nand2_1 U11099 ( .ip1(i_i2c_U_dff_rx_mem[22]), .ip2(n9170), .op(n9143) );
  and2_1 U11100 ( .ip1(i_i2c_U_dff_rx_mem[6]), .ip2(n11190), .op(n9140) );
  nand2_1 U11101 ( .ip1(i_i2c_U_dff_rx_mem[54]), .ip2(n9178), .op(n9138) );
  nand2_1 U11102 ( .ip1(i_i2c_U_dff_rx_mem[46]), .ip2(n9167), .op(n9137) );
  nand2_1 U11103 ( .ip1(i_i2c_U_dff_rx_mem[14]), .ip2(n9177), .op(n9136) );
  nand2_1 U11104 ( .ip1(i_i2c_U_dff_rx_mem[30]), .ip2(n9166), .op(n9135) );
  nand4_1 U11105 ( .ip1(n9138), .ip2(n9137), .ip3(n9136), .ip4(n9135), .op(
        n9139) );
  not_ab_or_c_or_d U11106 ( .ip1(n9169), .ip2(i_i2c_U_dff_rx_mem[38]), .ip3(
        n9140), .ip4(n9139), .op(n9142) );
  nand2_1 U11107 ( .ip1(i_i2c_U_dff_rx_mem[62]), .ip2(n9168), .op(n9141) );
  nand3_1 U11108 ( .ip1(n9143), .ip2(n9142), .ip3(n9141), .op(
        i_i2c_rx_pop_data[6]) );
  nand2_1 U11109 ( .ip1(i_i2c_U_dff_rx_mem[27]), .ip2(n9166), .op(n9152) );
  and2_1 U11110 ( .ip1(i_i2c_U_dff_rx_mem[3]), .ip2(n11190), .op(n9149) );
  nand2_1 U11111 ( .ip1(i_i2c_U_dff_rx_mem[59]), .ip2(n9168), .op(n9147) );
  nand2_1 U11112 ( .ip1(i_i2c_U_dff_rx_mem[35]), .ip2(n9169), .op(n9146) );
  nand2_1 U11113 ( .ip1(i_i2c_U_dff_rx_mem[11]), .ip2(n9177), .op(n9145) );
  nand2_1 U11114 ( .ip1(i_i2c_U_dff_rx_mem[51]), .ip2(n9178), .op(n9144) );
  nand4_1 U11115 ( .ip1(n9147), .ip2(n9146), .ip3(n9145), .ip4(n9144), .op(
        n9148) );
  not_ab_or_c_or_d U11116 ( .ip1(n9170), .ip2(i_i2c_U_dff_rx_mem[19]), .ip3(
        n9149), .ip4(n9148), .op(n9151) );
  nand2_1 U11117 ( .ip1(i_i2c_U_dff_rx_mem[43]), .ip2(n9167), .op(n9150) );
  nand3_1 U11118 ( .ip1(n9152), .ip2(n9151), .ip3(n9150), .op(
        i_i2c_rx_pop_data[3]) );
  xor2_1 U11119 ( .ip1(n9153), .ip2(i_i2c_tx_abrt_source[6]), .op(n5189) );
  nor2_1 U11120 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_scl_edg_hl_q), .ip2(n9154), 
        .op(n9156) );
  nand2_1 U11121 ( .ip1(i_i2c_slv_tx_ack_vld), .ip2(i_i2c_sda_vld), .op(n9155)
         );
  mux2_1 U11122 ( .ip1(n10579), .ip2(n9156), .s(n9155), .op(n5072) );
  nand2_1 U11123 ( .ip1(i_i2c_U_dff_rx_mem[34]), .ip2(n9169), .op(n9165) );
  and2_1 U11124 ( .ip1(i_i2c_U_dff_rx_mem[2]), .ip2(n11190), .op(n9162) );
  nand2_1 U11125 ( .ip1(i_i2c_U_dff_rx_mem[10]), .ip2(n9177), .op(n9160) );
  nand2_1 U11126 ( .ip1(i_i2c_U_dff_rx_mem[58]), .ip2(n9168), .op(n9159) );
  nand2_1 U11127 ( .ip1(i_i2c_U_dff_rx_mem[18]), .ip2(n9170), .op(n9158) );
  nand2_1 U11128 ( .ip1(i_i2c_U_dff_rx_mem[26]), .ip2(n9166), .op(n9157) );
  nand4_1 U11129 ( .ip1(n9160), .ip2(n9159), .ip3(n9158), .ip4(n9157), .op(
        n9161) );
  not_ab_or_c_or_d U11130 ( .ip1(n9167), .ip2(i_i2c_U_dff_rx_mem[42]), .ip3(
        n9162), .ip4(n9161), .op(n9164) );
  nand2_1 U11131 ( .ip1(i_i2c_U_dff_rx_mem[50]), .ip2(n9178), .op(n9163) );
  nand3_1 U11132 ( .ip1(n9165), .ip2(n9164), .ip3(n9163), .op(
        i_i2c_rx_pop_data[2]) );
  nand2_1 U11133 ( .ip1(i_i2c_U_dff_rx_mem[25]), .ip2(n9166), .op(n9181) );
  and2_1 U11134 ( .ip1(i_i2c_U_dff_rx_mem[1]), .ip2(n11190), .op(n9176) );
  nand2_1 U11135 ( .ip1(i_i2c_U_dff_rx_mem[41]), .ip2(n9167), .op(n9174) );
  nand2_1 U11136 ( .ip1(i_i2c_U_dff_rx_mem[57]), .ip2(n9168), .op(n9173) );
  nand2_1 U11137 ( .ip1(i_i2c_U_dff_rx_mem[33]), .ip2(n9169), .op(n9172) );
  nand2_1 U11138 ( .ip1(i_i2c_U_dff_rx_mem[17]), .ip2(n9170), .op(n9171) );
  nand4_1 U11139 ( .ip1(n9174), .ip2(n9173), .ip3(n9172), .ip4(n9171), .op(
        n9175) );
  not_ab_or_c_or_d U11140 ( .ip1(n9177), .ip2(i_i2c_U_dff_rx_mem[9]), .ip3(
        n9176), .ip4(n9175), .op(n9180) );
  nand2_1 U11141 ( .ip1(i_i2c_U_dff_rx_mem[49]), .ip2(n9178), .op(n9179) );
  nand3_1 U11142 ( .ip1(n9181), .ip2(n9180), .ip3(n9179), .op(
        i_i2c_rx_pop_data[1]) );
  and2_1 U11143 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_chk_win), .ip2(n9182), .op(n9184) );
  mux2_1 U11144 ( .ip1(i_i2c_ic_abort_sync), .ip2(n9184), .s(n9183), .op(n4181) );
  nor2_1 U11145 ( .ip1(n6470), .ip2(n9667), .op(n9185) );
  xor2_1 U11146 ( .ip1(i_i2c_tx_abrt_source[3]), .ip2(n9185), .op(n5193) );
  inv_1 U11147 ( .ip(i_i2c_rx_gen_call), .op(n9186) );
  nor2_1 U11148 ( .ip1(i_i2c_U_DW_apb_i2c_toggle_rx_gen_call_r), .ip2(n9186), 
        .op(n9187) );
  xor2_1 U11149 ( .ip1(i_i2c_rx_gen_call_flg), .ip2(n9187), .op(n4172) );
  nor2_1 U11150 ( .ip1(n9188), .ip2(n9414), .op(n9189) );
  xor2_1 U11151 ( .ip1(i_i2c_tx_abrt_source[9]), .ip2(n9189), .op(n4861) );
  mux2_1 U11152 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[5]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[5]), .s(n11359), .op(n4849) );
  mux2_1 U11153 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[12]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[12]), .s(n11359), .op(n4846) );
  mux2_1 U11154 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[3]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[3]), .s(n11359), .op(n4851) );
  mux2_1 U11155 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[7]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[7]), .s(n11359), .op(n4847) );
  mux2_1 U11156 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_hwrite_c), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite), .s(n11359), .op(n4853) );
  mux2_1 U11157 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[4]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[4]), .s(n11359), .op(n4850) );
  mux2_1 U11158 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[6]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[6]), .s(n11359), .op(n4848) );
  mux2_1 U11159 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[2]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[2]), .s(n11359), .op(n4852) );
  inv_1 U11160 ( .ip(i_ssi_U_mstfsm_bit_cnt[0]), .op(n9190) );
  xor2_1 U11161 ( .ip1(n9190), .ip2(n10473), .op(n9191) );
  nand2_1 U11162 ( .ip1(ex_i_ahb_AHB_Slave_PID_hresp[1]), .ip2(
        i_ahb_U_mux_hsel_prev[4]), .op(n9194) );
  nand2_1 U11163 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hresp[1]), .op(
        n9193) );
  nand2_1 U11164 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hresp[1]), .op(
        n9192) );
  nand2_1 U11165 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hresp[0]), .op(
        n9200) );
  nand2_1 U11166 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hresp[0]), .op(n9199) );
  nand3_1 U11167 ( .ip1(n9196), .ip2(i_ahb_hresp_none_0_), .ip3(n9195), .op(
        n9198) );
  nand2_1 U11168 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hresp[0]), .op(
        n9197) );
  nand2_1 U11169 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[27]), .op(
        n9204) );
  nand2_1 U11170 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[27]), .op(n9203) );
  nand2_1 U11171 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[27]), .op(
        n9202) );
  and2_1 U11172 ( .ip1(n9335), .ip2(n9358), .op(n9205) );
  nand2_1 U11173 ( .ip1(n9205), .ip2(i_ssi_prdata[27]), .op(n9201) );
  nand2_1 U11174 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[31]), .op(n9209) );
  nand2_1 U11175 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[31]), .op(
        n9208) );
  nand2_1 U11176 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[31]), .op(
        n9207) );
  nand2_1 U11177 ( .ip1(n9205), .ip2(i_ssi_prdata[31]), .op(n9206) );
  nand2_1 U11178 ( .ip1(n9358), .ip2(n9210), .op(n9214) );
  nand2_1 U11179 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[20]), .op(
        n9213) );
  nand2_1 U11180 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[20]), .op(
        n9212) );
  nand2_1 U11181 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[20]), .op(n9211) );
  nand2_1 U11182 ( .ip1(n9358), .ip2(n9215), .op(n9219) );
  nand2_1 U11183 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[13]), .op(
        n9218) );
  nand2_1 U11184 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[13]), .op(n9217) );
  nand2_1 U11185 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[13]), .op(
        n9216) );
  nand2_1 U11186 ( .ip1(n9358), .ip2(n9220), .op(n9224) );
  nand2_1 U11187 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[16]), .op(
        n9223) );
  nand2_1 U11188 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[16]), .op(n9222) );
  nand2_1 U11189 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[16]), .op(
        n9221) );
  nand2_1 U11190 ( .ip1(n9358), .ip2(n9225), .op(n9229) );
  nand2_1 U11191 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[2]), .op(
        n9228) );
  nand2_1 U11192 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[2]), .op(
        n9227) );
  nand2_1 U11193 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[2]), .op(n9226) );
  nand2_1 U11194 ( .ip1(n9358), .ip2(n9230), .op(n9234) );
  nand2_1 U11195 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[5]), .op(
        n9233) );
  nand2_1 U11196 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[5]), .op(n9232) );
  nand2_1 U11197 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[5]), .op(
        n9231) );
  nand2_1 U11198 ( .ip1(n9358), .ip2(n9235), .op(n9239) );
  nand2_1 U11199 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[12]), .op(
        n9238) );
  nand2_1 U11200 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[12]), .op(n9237) );
  nand2_1 U11201 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[12]), .op(
        n9236) );
  nand2_1 U11202 ( .ip1(n9358), .ip2(n9240), .op(n9244) );
  nand2_1 U11203 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[9]), .op(
        n9243) );
  nand2_1 U11204 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[9]), .op(n9242) );
  nand2_1 U11205 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[9]), .op(
        n9241) );
  nand2_1 U11206 ( .ip1(n9358), .ip2(n9245), .op(n9249) );
  nand2_1 U11207 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[10]), .op(
        n9248) );
  nand2_1 U11208 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[10]), .op(n9247) );
  nand2_1 U11209 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[10]), .op(
        n9246) );
  nand2_1 U11210 ( .ip1(n9358), .ip2(n9250), .op(n9254) );
  nand2_1 U11211 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[21]), .op(
        n9253) );
  nand2_1 U11212 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[21]), .op(
        n9252) );
  nand2_1 U11213 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[21]), .op(n9251) );
  nand2_1 U11214 ( .ip1(n9358), .ip2(n9255), .op(n9259) );
  nand2_1 U11215 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[11]), .op(
        n9258) );
  nand2_1 U11216 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[11]), .op(n9257) );
  nand2_1 U11217 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[11]), .op(
        n9256) );
  nand2_1 U11218 ( .ip1(n9358), .ip2(n9260), .op(n9264) );
  nand2_1 U11219 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[3]), .op(
        n9263) );
  nand2_1 U11220 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[3]), .op(n9262) );
  nand2_1 U11221 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[3]), .op(
        n9261) );
  nand2_1 U11222 ( .ip1(n9358), .ip2(n9265), .op(n9269) );
  nand2_1 U11223 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[17]), .op(
        n9268) );
  nand2_1 U11224 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[17]), .op(n9267) );
  nand2_1 U11225 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[17]), .op(
        n9266) );
  nand2_1 U11226 ( .ip1(n9358), .ip2(n9270), .op(n9274) );
  nand2_1 U11227 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[1]), .op(
        n9273) );
  nand2_1 U11228 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[1]), .op(n9272) );
  nand2_1 U11229 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[1]), .op(
        n9271) );
  nand2_1 U11230 ( .ip1(n9358), .ip2(n9275), .op(n9279) );
  nand2_1 U11231 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[4]), .op(
        n9278) );
  nand2_1 U11232 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[4]), .op(n9277) );
  nand2_1 U11233 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[4]), .op(
        n9276) );
  nand2_1 U11234 ( .ip1(n9358), .ip2(n9280), .op(n9284) );
  nand2_1 U11235 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[0]), .op(
        n9283) );
  nand2_1 U11236 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[0]), .op(
        n9282) );
  nand2_1 U11237 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[0]), .op(n9281) );
  nand2_1 U11238 ( .ip1(n9358), .ip2(n9285), .op(n9289) );
  nand2_1 U11239 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[14]), .op(
        n9288) );
  nand2_1 U11240 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[14]), .op(
        n9287) );
  nand2_1 U11241 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[14]), .op(n9286) );
  nand2_1 U11242 ( .ip1(n9358), .ip2(n9290), .op(n9294) );
  nand2_1 U11243 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[8]), .op(
        n9293) );
  nand2_1 U11244 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[8]), .op(n9292) );
  nand2_1 U11245 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[8]), .op(
        n9291) );
  nand2_1 U11246 ( .ip1(n9358), .ip2(n9295), .op(n9299) );
  nand2_1 U11247 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[7]), .op(
        n9298) );
  nand2_1 U11248 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[7]), .op(
        n9297) );
  nand2_1 U11249 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[7]), .op(n9296) );
  nand2_1 U11250 ( .ip1(n9358), .ip2(n9300), .op(n9304) );
  nand2_1 U11251 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[18]), .op(
        n9303) );
  nand2_1 U11252 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[18]), .op(
        n9302) );
  nand2_1 U11253 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[18]), .op(n9301) );
  nand2_1 U11254 ( .ip1(n9358), .ip2(n9305), .op(n9309) );
  nand2_1 U11255 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[6]), .op(
        n9308) );
  nand2_1 U11256 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[6]), .op(n9307) );
  nand2_1 U11257 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[6]), .op(
        n9306) );
  nand2_1 U11258 ( .ip1(n9358), .ip2(n9310), .op(n9314) );
  nand2_1 U11259 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[19]), .op(
        n9313) );
  nand2_1 U11260 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[19]), .op(
        n9312) );
  nand2_1 U11261 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[19]), .op(n9311) );
  nand2_1 U11262 ( .ip1(n9358), .ip2(n9315), .op(n9319) );
  nand2_1 U11263 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[15]), .op(
        n9318) );
  nand2_1 U11264 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[15]), .op(
        n9317) );
  nand2_1 U11265 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[15]), .op(n9316) );
  nand2_1 U11266 ( .ip1(n9358), .ip2(n9320), .op(n9324) );
  nand2_1 U11267 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[25]), .op(
        n9323) );
  nand2_1 U11268 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[25]), .op(
        n9322) );
  nand2_1 U11269 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[25]), .op(n9321) );
  nand2_1 U11270 ( .ip1(n9358), .ip2(n9325), .op(n9329) );
  nand2_1 U11271 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[23]), .op(
        n9328) );
  nand2_1 U11272 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[23]), .op(
        n9327) );
  nand2_1 U11273 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[23]), .op(n9326) );
  nand2_1 U11274 ( .ip1(n9358), .ip2(n9330), .op(n9334) );
  nand2_1 U11275 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[26]), .op(
        n9333) );
  nand2_1 U11276 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[26]), .op(
        n9332) );
  nand2_1 U11277 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[26]), .op(n9331) );
  nand2_1 U11278 ( .ip1(n9358), .ip2(n9336), .op(n9340) );
  nand2_1 U11279 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[22]), .op(
        n9339) );
  nand2_1 U11280 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[22]), .op(n9338) );
  nand2_1 U11281 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[22]), .op(
        n9337) );
  nand2_1 U11282 ( .ip1(n9358), .ip2(n9341), .op(n9345) );
  nand2_1 U11283 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[29]), .op(
        n9344) );
  nand2_1 U11284 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[29]), .op(
        n9343) );
  nand2_1 U11285 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[29]), .op(n9342) );
  nand2_1 U11286 ( .ip1(n9358), .ip2(n9346), .op(n9350) );
  nand2_1 U11287 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[24]), .op(
        n9349) );
  nand2_1 U11288 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[24]), .op(n9348) );
  nand2_1 U11289 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[24]), .op(
        n9347) );
  nand2_1 U11290 ( .ip1(n9358), .ip2(n9351), .op(n9355) );
  nand2_1 U11291 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[28]), .op(
        n9354) );
  nand2_1 U11292 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[28]), .op(
        n9353) );
  nand2_1 U11293 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[28]), .op(n9352) );
  nand2_1 U11294 ( .ip1(n9358), .ip2(n9357), .op(n9364) );
  nand2_1 U11295 ( .ip1(n9359), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[30]), .op(
        n9363) );
  nand2_1 U11296 ( .ip1(n9360), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[30]), .op(
        n9362) );
  nand2_1 U11297 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[30]), .op(n9361) );
  and2_1 U11298 ( .ip1(i_ssi_U_mstfsm_bit_cnt[0]), .ip2(
        i_ssi_U_mstfsm_bit_cnt[1]), .op(n9365) );
  and2_1 U11299 ( .ip1(n10473), .ip2(n9365), .op(n10476) );
  nand2_1 U11300 ( .ip1(n10476), .ip2(i_ssi_U_mstfsm_bit_cnt[2]), .op(n10481)
         );
  nor2_1 U11301 ( .ip1(n10482), .ip2(n10481), .op(n10479) );
  xor2_1 U11302 ( .ip1(n9366), .ip2(n10479), .op(n9367) );
  buf_2 U11303 ( .ip(n9372), .op(n9395) );
  nand3_1 U11304 ( .ip1(i_apb_U_DW_apb_ahbsif_state[1]), .ip2(n10106), .ip3(
        n10108), .op(n9373) );
  nand3_1 U11305 ( .ip1(n9897), .ip2(n9377), .ip3(n9373), .op(n9393) );
  or2_1 U11306 ( .ip1(i_apb_pclk_en), .ip2(n10024), .op(n9376) );
  or2_1 U11307 ( .ip1(n9374), .ip2(n10024), .op(n9375) );
  nor2_1 U11308 ( .ip1(n10108), .ip2(n9377), .op(n9390) );
  nor2_1 U11309 ( .ip1(n9380), .ip2(n9379), .op(n10025) );
  nor4_1 U11310 ( .ip1(n10025), .ip2(n9383), .ip3(n9382), .ip4(n10106), .op(
        n9389) );
  nand2_1 U11311 ( .ip1(i_apb_U_DW_apb_ahbsif_state[0]), .ip2(n9384), .op(
        n9387) );
  nand2_1 U11312 ( .ip1(i_apb_U_DW_apb_ahbsif_state[1]), .ip2(n10106), .op(
        n9386) );
  nor2_1 U11313 ( .ip1(n10108), .ip2(n9387), .op(n9385) );
  not_ab_or_c_or_d U11314 ( .ip1(n10108), .ip2(n9387), .ip3(n9386), .ip4(n9385), .op(n9388) );
  and3_1 U11315 ( .ip1(n9999), .ip2(i_i2c_U_DW_apb_i2c_tx_shift_slv_data_sda), 
        .ip3(i_i2c_U_DW_apb_i2c_tx_shift_data_sda), .op(n9394) );
  xor2_1 U11316 ( .ip1(n5739), .ip2(i_ssi_tx_pop), .op(n4585) );
  mux2_1 U11317 ( .ip1(n11110), .ip2(n11283), .s(i_i2c_tx_abrt_source[12]), 
        .op(n4182) );
  mux2_1 U11318 ( .ip1(n9401), .ip2(n9400), .s(i_i2c_tx_abrt_source[16]), .op(
        n5205) );
  inv_1 U11319 ( .ip(n9404), .op(n9406) );
  nor2_1 U11320 ( .ip1(n9406), .ip2(n9405), .op(n9407) );
  mux2_1 U11321 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_sda_data_int), .ip2(n9408), 
        .s(n9407), .op(n5136) );
  mux2_1 U11322 ( .ip1(i_i2c_prdata[29]), .ip2(i_i2c_iprdata[29]), .s(n11762), 
        .op(n4690) );
  mux2_1 U11323 ( .ip1(i_i2c_prdata[19]), .ip2(i_i2c_iprdata[19]), .s(n11762), 
        .op(n4680) );
  mux2_1 U11324 ( .ip1(i_i2c_prdata[16]), .ip2(i_i2c_iprdata[16]), .s(n11762), 
        .op(n4677) );
  mux2_1 U11325 ( .ip1(i_i2c_prdata[20]), .ip2(i_i2c_iprdata[20]), .s(n11762), 
        .op(n4681) );
  mux2_1 U11326 ( .ip1(i_i2c_prdata[17]), .ip2(i_i2c_iprdata[17]), .s(n11762), 
        .op(n4678) );
  inv_1 U11327 ( .ip(i_i2c_tx_abrt_source[4]), .op(n9412) );
  nand2_1 U11328 ( .ip1(n9410), .ip2(n9409), .op(n9411) );
  mux2_1 U11329 ( .ip1(n9412), .ip2(i_i2c_tx_abrt_source[4]), .s(n9411), .op(
        n5186) );
  mux2_1 U11330 ( .ip1(i_i2c_prdata[15]), .ip2(i_i2c_iprdata[15]), .s(n11762), 
        .op(n4676) );
  mux2_1 U11331 ( .ip1(i_i2c_prdata[14]), .ip2(i_i2c_iprdata[14]), .s(n11762), 
        .op(n4675) );
  mux2_1 U11332 ( .ip1(i_i2c_prdata[13]), .ip2(i_i2c_iprdata[13]), .s(n11762), 
        .op(n4674) );
  mux2_1 U11333 ( .ip1(i_i2c_prdata[9]), .ip2(i_i2c_iprdata[9]), .s(n11762), 
        .op(n4670) );
  nand3_1 U11334 ( .ip1(i_i2c_rx_push_sync), .ip2(i_i2c_rx_wr_addr[0]), .ip3(
        n11191), .op(n11194) );
  inv_1 U11335 ( .ip(i_i2c_rx_wr_addr[2]), .op(n9767) );
  or3_1 U11336 ( .ip1(n11194), .ip2(n9767), .ip3(i_i2c_rx_wr_addr[1]), .op(
        n9413) );
  mux2_1 U11337 ( .ip1(i_i2c_rx_push_data[1]), .ip2(i_i2c_U_dff_rx_mem[17]), 
        .s(n9413), .op(n4918) );
  mux2_1 U11338 ( .ip1(i_i2c_rx_push_data[7]), .ip2(i_i2c_U_dff_rx_mem[23]), 
        .s(n9413), .op(n4870) );
  mux2_1 U11339 ( .ip1(i_i2c_rx_push_data[5]), .ip2(i_i2c_U_dff_rx_mem[21]), 
        .s(n9413), .op(n4886) );
  mux2_1 U11340 ( .ip1(i_i2c_rx_push_data[0]), .ip2(i_i2c_U_dff_rx_mem[16]), 
        .s(n9413), .op(n4926) );
  mux2_1 U11341 ( .ip1(i_i2c_rx_push_data[4]), .ip2(i_i2c_U_dff_rx_mem[20]), 
        .s(n9413), .op(n4894) );
  mux2_1 U11342 ( .ip1(i_i2c_rx_push_data[2]), .ip2(i_i2c_U_dff_rx_mem[18]), 
        .s(n9413), .op(n4910) );
  mux2_1 U11343 ( .ip1(i_i2c_rx_push_data[3]), .ip2(i_i2c_U_dff_rx_mem[19]), 
        .s(n9413), .op(n4902) );
  mux2_1 U11344 ( .ip1(i_i2c_rx_push_data[6]), .ip2(i_i2c_U_dff_rx_mem[22]), 
        .s(n9413), .op(n4878) );
  nor2_1 U11345 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv), .ip2(n9414), 
        .op(n9415) );
  xor2_1 U11346 ( .ip1(i_i2c_tx_abrt_source[8]), .ip2(n9415), .op(n4863) );
  nand2_1 U11347 ( .ip1(n9735), .ip2(i_i2c_ic_tar[2]), .op(n9419) );
  nand2_1 U11348 ( .ip1(n9429), .ip2(i_i2c_ic_tar[9]), .op(n9418) );
  nand2_1 U11349 ( .ip1(n9448), .ip2(i_i2c_ic_tar[1]), .op(n9417) );
  nand3_1 U11350 ( .ip1(n9419), .ip2(n9418), .ip3(n9417), .op(n9420) );
  ab_or_c_or_d U11351 ( .ip1(n9740), .ip2(i_i2c_ic_hs_maddr[2]), .ip3(n9421), 
        .ip4(n9420), .op(n9422) );
  nor2_1 U11352 ( .ip1(i_i2c_debug_wr), .ip2(n11160), .op(n9743) );
  mux2_1 U11353 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[2]), .ip2(
        n9422), .s(n9743), .op(n5045) );
  nand2_1 U11354 ( .ip1(n9735), .ip2(i_i2c_ic_tar[3]), .op(n9426) );
  inv_1 U11355 ( .ip(n10413), .op(n9423) );
  nand2_1 U11356 ( .ip1(n9423), .ip2(i_i2c_tx_fifo_data_buf[3]), .op(n9425) );
  nand2_1 U11357 ( .ip1(n9448), .ip2(i_i2c_ic_tar[2]), .op(n9424) );
  nand4_1 U11358 ( .ip1(n9725), .ip2(n9426), .ip3(n9425), .ip4(n9424), .op(
        n9427) );
  mux2_1 U11359 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[3]), .ip2(
        n9427), .s(n9743), .op(n5044) );
  nand2_1 U11360 ( .ip1(n9735), .ip2(i_i2c_ic_tar[1]), .op(n9432) );
  nand2_1 U11361 ( .ip1(n9429), .ip2(i_i2c_ic_tar[8]), .op(n9431) );
  nand2_1 U11362 ( .ip1(n9448), .ip2(i_i2c_ic_tar[0]), .op(n9430) );
  nand3_1 U11363 ( .ip1(n9432), .ip2(n9431), .ip3(n9430), .op(n9433) );
  ab_or_c_or_d U11364 ( .ip1(n9740), .ip2(i_i2c_ic_hs_maddr[1]), .ip3(n9434), 
        .ip4(n9433), .op(n9435) );
  mux2_1 U11365 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[1]), .ip2(
        n9435), .s(n9743), .op(n5046) );
  nand2_1 U11366 ( .ip1(n9448), .ip2(i_i2c_ic_tar[3]), .op(n9438) );
  nand2_1 U11367 ( .ip1(n9449), .ip2(i_i2c_tx_fifo_data_buf[4]), .op(n9437) );
  nand2_1 U11368 ( .ip1(n9735), .ip2(i_i2c_ic_tar[4]), .op(n9436) );
  mux2_1 U11369 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[4]), .ip2(
        n9439), .s(n9743), .op(n5043) );
  nand2_1 U11370 ( .ip1(n9448), .ip2(i_i2c_ic_tar[4]), .op(n9442) );
  nand2_1 U11371 ( .ip1(n9449), .ip2(i_i2c_tx_fifo_data_buf[5]), .op(n9441) );
  nand2_1 U11372 ( .ip1(n9735), .ip2(i_i2c_ic_tar[5]), .op(n9440) );
  mux2_1 U11373 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[5]), .ip2(
        n9443), .s(n9743), .op(n5042) );
  nand2_1 U11374 ( .ip1(n9448), .ip2(i_i2c_ic_tar[6]), .op(n9446) );
  nand2_1 U11375 ( .ip1(n9449), .ip2(i_i2c_tx_fifo_data_buf[7]), .op(n9445) );
  nand2_1 U11376 ( .ip1(n9735), .ip2(i_i2c_ic_tar[7]), .op(n9444) );
  mux2_1 U11377 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[7]), .ip2(
        n9447), .s(n9743), .op(n5040) );
  nand2_1 U11378 ( .ip1(n9448), .ip2(i_i2c_ic_tar[5]), .op(n9452) );
  nand2_1 U11379 ( .ip1(n9449), .ip2(i_i2c_tx_fifo_data_buf[6]), .op(n9451) );
  nand2_1 U11380 ( .ip1(n9735), .ip2(i_i2c_ic_tar[6]), .op(n9450) );
  mux2_1 U11381 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[6]), .ip2(
        n9453), .s(n9743), .op(n5041) );
  nor3_1 U11382 ( .ip1(i_i2c_tx_rd_addr[2]), .ip2(i_i2c_tx_rd_addr[1]), .ip3(
        n9456), .op(n9559) );
  nand2_1 U11383 ( .ip1(n9559), .ip2(i_i2c_U_dff_tx_mem[55]), .op(n9467) );
  inv_1 U11384 ( .ip(i_i2c_tx_rd_addr[1]), .op(n9455) );
  nor3_1 U11385 ( .ip1(i_i2c_tx_rd_addr[2]), .ip2(i_i2c_tx_rd_addr[0]), .ip3(
        n9455), .op(n9551) );
  nand3_1 U11386 ( .ip1(i_i2c_tx_rd_addr[2]), .ip2(i_i2c_tx_rd_addr[1]), .ip3(
        i_i2c_tx_rd_addr[0]), .op(n9548) );
  inv_1 U11387 ( .ip(i_i2c_U_dff_tx_mem[1]), .op(n9454) );
  nor2_1 U11388 ( .ip1(n9548), .ip2(n9454), .op(n9463) );
  nor3_1 U11389 ( .ip1(i_i2c_tx_rd_addr[2]), .ip2(i_i2c_tx_rd_addr[1]), .ip3(
        i_i2c_tx_rd_addr[0]), .op(n9552) );
  nand2_1 U11390 ( .ip1(n9552), .ip2(i_i2c_U_dff_tx_mem[64]), .op(n9461) );
  nor3_1 U11391 ( .ip1(i_i2c_tx_rd_addr[0]), .ip2(n9455), .ip3(n9457), .op(
        n9549) );
  nand2_1 U11392 ( .ip1(n9549), .ip2(i_i2c_U_dff_tx_mem[10]), .op(n9460) );
  nor3_1 U11393 ( .ip1(i_i2c_tx_rd_addr[1]), .ip2(n9457), .ip3(n9456), .op(
        n9550) );
  nand2_1 U11394 ( .ip1(n9550), .ip2(i_i2c_U_dff_tx_mem[19]), .op(n9459) );
  nor3_1 U11395 ( .ip1(i_i2c_tx_rd_addr[1]), .ip2(i_i2c_tx_rd_addr[0]), .ip3(
        n9457), .op(n9546) );
  nand2_1 U11396 ( .ip1(n9546), .ip2(i_i2c_U_dff_tx_mem[28]), .op(n9458) );
  nand4_1 U11397 ( .ip1(n9461), .ip2(n9460), .ip3(n9459), .ip4(n9458), .op(
        n9462) );
  not_ab_or_c_or_d U11398 ( .ip1(n9551), .ip2(i_i2c_U_dff_tx_mem[46]), .ip3(
        n9463), .ip4(n9462), .op(n9466) );
  nor2_1 U11399 ( .ip1(i_i2c_tx_rd_addr[2]), .ip2(n9464), .op(n9560) );
  nand2_1 U11400 ( .ip1(n9560), .ip2(i_i2c_U_dff_tx_mem[37]), .op(n9465) );
  nand3_1 U11401 ( .ip1(n9467), .ip2(n9466), .ip3(n9465), .op(n9468) );
  mux2_1 U11402 ( .ip1(i_i2c_tx_fifo_data_buf[1]), .ip2(n9468), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .op(n5228) );
  nand2_1 U11403 ( .ip1(i_i2c_U_dff_tx_mem[16]), .ip2(n9549), .op(n9478) );
  inv_1 U11404 ( .ip(i_i2c_U_dff_tx_mem[7]), .op(n9469) );
  nor2_1 U11405 ( .ip1(n9548), .ip2(n9469), .op(n9475) );
  nand2_1 U11406 ( .ip1(n9546), .ip2(i_i2c_U_dff_tx_mem[34]), .op(n9473) );
  nand2_1 U11407 ( .ip1(n9559), .ip2(i_i2c_U_dff_tx_mem[61]), .op(n9472) );
  nand2_1 U11408 ( .ip1(n9560), .ip2(i_i2c_U_dff_tx_mem[43]), .op(n9471) );
  nand2_1 U11409 ( .ip1(n9552), .ip2(i_i2c_U_dff_tx_mem[70]), .op(n9470) );
  nand4_1 U11410 ( .ip1(n9473), .ip2(n9472), .ip3(n9471), .ip4(n9470), .op(
        n9474) );
  not_ab_or_c_or_d U11411 ( .ip1(n9550), .ip2(i_i2c_U_dff_tx_mem[25]), .ip3(
        n9475), .ip4(n9474), .op(n9477) );
  nand2_1 U11412 ( .ip1(n9551), .ip2(i_i2c_U_dff_tx_mem[52]), .op(n9476) );
  nand3_1 U11413 ( .ip1(n9478), .ip2(n9477), .ip3(n9476), .op(n9479) );
  mux2_1 U11414 ( .ip1(i_i2c_tx_fifo_data_buf[7]), .ip2(n9479), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .op(n5222) );
  nand2_1 U11415 ( .ip1(i_i2c_U_dff_tx_mem[29]), .ip2(n9546), .op(n9489) );
  inv_1 U11416 ( .ip(i_i2c_U_dff_tx_mem[2]), .op(n9480) );
  nor2_1 U11417 ( .ip1(n9548), .ip2(n9480), .op(n9486) );
  nand2_1 U11418 ( .ip1(n9551), .ip2(i_i2c_U_dff_tx_mem[47]), .op(n9484) );
  nand2_1 U11419 ( .ip1(n9552), .ip2(i_i2c_U_dff_tx_mem[65]), .op(n9483) );
  nand2_1 U11420 ( .ip1(n9550), .ip2(i_i2c_U_dff_tx_mem[20]), .op(n9482) );
  nand2_1 U11421 ( .ip1(n9559), .ip2(i_i2c_U_dff_tx_mem[56]), .op(n9481) );
  nand4_1 U11422 ( .ip1(n9484), .ip2(n9483), .ip3(n9482), .ip4(n9481), .op(
        n9485) );
  not_ab_or_c_or_d U11423 ( .ip1(i_i2c_U_dff_tx_mem[11]), .ip2(n9549), .ip3(
        n9486), .ip4(n9485), .op(n9488) );
  nand2_1 U11424 ( .ip1(n9560), .ip2(i_i2c_U_dff_tx_mem[38]), .op(n9487) );
  nand3_1 U11425 ( .ip1(n9489), .ip2(n9488), .ip3(n9487), .op(n9490) );
  mux2_1 U11426 ( .ip1(i_i2c_tx_fifo_data_buf[2]), .ip2(n9490), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .op(n5227) );
  nand2_1 U11427 ( .ip1(i_i2c_U_dff_tx_mem[54]), .ip2(n9559), .op(n9500) );
  inv_1 U11428 ( .ip(i_i2c_U_dff_tx_mem[0]), .op(n9491) );
  nor2_1 U11429 ( .ip1(n9491), .ip2(n9548), .op(n9497) );
  nand2_1 U11430 ( .ip1(i_i2c_U_dff_tx_mem[9]), .ip2(n9549), .op(n9495) );
  nand2_1 U11431 ( .ip1(i_i2c_U_dff_tx_mem[45]), .ip2(n9551), .op(n9494) );
  nand2_1 U11432 ( .ip1(i_i2c_U_dff_tx_mem[63]), .ip2(n9552), .op(n9493) );
  nand2_1 U11433 ( .ip1(i_i2c_U_dff_tx_mem[36]), .ip2(n9560), .op(n9492) );
  nand4_1 U11434 ( .ip1(n9495), .ip2(n9494), .ip3(n9493), .ip4(n9492), .op(
        n9496) );
  not_ab_or_c_or_d U11435 ( .ip1(n9550), .ip2(i_i2c_U_dff_tx_mem[18]), .ip3(
        n9497), .ip4(n9496), .op(n9499) );
  nand2_1 U11436 ( .ip1(i_i2c_U_dff_tx_mem[27]), .ip2(n9546), .op(n9498) );
  nand3_1 U11437 ( .ip1(n9500), .ip2(n9499), .ip3(n9498), .op(n9501) );
  mux2_1 U11438 ( .ip1(i_i2c_tx_fifo_data_buf[0]), .ip2(n9501), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .op(n5229) );
  nand2_1 U11439 ( .ip1(n9546), .ip2(i_i2c_U_dff_tx_mem[35]), .op(n9511) );
  inv_1 U11440 ( .ip(i_i2c_U_dff_tx_mem[8]), .op(n9502) );
  nor2_1 U11441 ( .ip1(n9548), .ip2(n9502), .op(n9508) );
  nand2_1 U11442 ( .ip1(n9559), .ip2(i_i2c_U_dff_tx_mem[62]), .op(n9506) );
  nand2_1 U11443 ( .ip1(n9552), .ip2(i_i2c_U_dff_tx_mem[71]), .op(n9505) );
  nand2_1 U11444 ( .ip1(n9549), .ip2(i_i2c_U_dff_tx_mem[17]), .op(n9504) );
  nand2_1 U11445 ( .ip1(n9550), .ip2(i_i2c_U_dff_tx_mem[26]), .op(n9503) );
  nand4_1 U11446 ( .ip1(n9506), .ip2(n9505), .ip3(n9504), .ip4(n9503), .op(
        n9507) );
  not_ab_or_c_or_d U11447 ( .ip1(n9560), .ip2(i_i2c_U_dff_tx_mem[44]), .ip3(
        n9508), .ip4(n9507), .op(n9510) );
  nand2_1 U11448 ( .ip1(n9551), .ip2(i_i2c_U_dff_tx_mem[53]), .op(n9509) );
  nand3_1 U11449 ( .ip1(n9511), .ip2(n9510), .ip3(n9509), .op(n9512) );
  mux2_1 U11450 ( .ip1(i_i2c_tx_fifo_data_buf[8]), .ip2(n9512), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .op(n5221) );
  nand2_1 U11451 ( .ip1(i_i2c_U_dff_tx_mem[33]), .ip2(n9546), .op(n9522) );
  inv_1 U11452 ( .ip(i_i2c_U_dff_tx_mem[6]), .op(n9513) );
  nor2_1 U11453 ( .ip1(n9548), .ip2(n9513), .op(n9519) );
  nand2_1 U11454 ( .ip1(n9550), .ip2(i_i2c_U_dff_tx_mem[24]), .op(n9517) );
  nand2_1 U11455 ( .ip1(n9559), .ip2(i_i2c_U_dff_tx_mem[60]), .op(n9516) );
  nand2_1 U11456 ( .ip1(n9552), .ip2(i_i2c_U_dff_tx_mem[69]), .op(n9515) );
  nand2_1 U11457 ( .ip1(n9549), .ip2(i_i2c_U_dff_tx_mem[15]), .op(n9514) );
  nand4_1 U11458 ( .ip1(n9517), .ip2(n9516), .ip3(n9515), .ip4(n9514), .op(
        n9518) );
  not_ab_or_c_or_d U11459 ( .ip1(n9560), .ip2(i_i2c_U_dff_tx_mem[42]), .ip3(
        n9519), .ip4(n9518), .op(n9521) );
  nand2_1 U11460 ( .ip1(n9551), .ip2(i_i2c_U_dff_tx_mem[51]), .op(n9520) );
  nand3_1 U11461 ( .ip1(n9522), .ip2(n9521), .ip3(n9520), .op(n9523) );
  mux2_1 U11462 ( .ip1(i_i2c_tx_fifo_data_buf[6]), .ip2(n9523), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .op(n5223) );
  nand2_1 U11463 ( .ip1(n9552), .ip2(i_i2c_U_dff_tx_mem[68]), .op(n9533) );
  inv_1 U11464 ( .ip(i_i2c_U_dff_tx_mem[5]), .op(n9524) );
  nor2_1 U11465 ( .ip1(n9548), .ip2(n9524), .op(n9530) );
  nand2_1 U11466 ( .ip1(n9550), .ip2(i_i2c_U_dff_tx_mem[23]), .op(n9528) );
  nand2_1 U11467 ( .ip1(n9546), .ip2(i_i2c_U_dff_tx_mem[32]), .op(n9527) );
  nand2_1 U11468 ( .ip1(n9551), .ip2(i_i2c_U_dff_tx_mem[50]), .op(n9526) );
  nand2_1 U11469 ( .ip1(n9559), .ip2(i_i2c_U_dff_tx_mem[59]), .op(n9525) );
  nand4_1 U11470 ( .ip1(n9528), .ip2(n9527), .ip3(n9526), .ip4(n9525), .op(
        n9529) );
  not_ab_or_c_or_d U11471 ( .ip1(i_i2c_U_dff_tx_mem[14]), .ip2(n9549), .ip3(
        n9530), .ip4(n9529), .op(n9532) );
  nand2_1 U11472 ( .ip1(n9560), .ip2(i_i2c_U_dff_tx_mem[41]), .op(n9531) );
  nand3_1 U11473 ( .ip1(n9533), .ip2(n9532), .ip3(n9531), .op(n9534) );
  mux2_1 U11474 ( .ip1(i_i2c_tx_fifo_data_buf[5]), .ip2(n9534), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .op(n5224) );
  nand2_1 U11475 ( .ip1(i_i2c_U_dff_tx_mem[22]), .ip2(n9550), .op(n9544) );
  inv_1 U11476 ( .ip(i_i2c_U_dff_tx_mem[4]), .op(n9535) );
  nor2_1 U11477 ( .ip1(n9548), .ip2(n9535), .op(n9541) );
  nand2_1 U11478 ( .ip1(n9549), .ip2(i_i2c_U_dff_tx_mem[13]), .op(n9539) );
  nand2_1 U11479 ( .ip1(n9551), .ip2(i_i2c_U_dff_tx_mem[49]), .op(n9538) );
  nand2_1 U11480 ( .ip1(n9546), .ip2(i_i2c_U_dff_tx_mem[31]), .op(n9537) );
  nand2_1 U11481 ( .ip1(n9552), .ip2(i_i2c_U_dff_tx_mem[67]), .op(n9536) );
  nand4_1 U11482 ( .ip1(n9539), .ip2(n9538), .ip3(n9537), .ip4(n9536), .op(
        n9540) );
  not_ab_or_c_or_d U11483 ( .ip1(i_i2c_U_dff_tx_mem[58]), .ip2(n9559), .ip3(
        n9541), .ip4(n9540), .op(n9543) );
  nand2_1 U11484 ( .ip1(n9560), .ip2(i_i2c_U_dff_tx_mem[40]), .op(n9542) );
  nand3_1 U11485 ( .ip1(n9544), .ip2(n9543), .ip3(n9542), .op(n9545) );
  mux2_1 U11486 ( .ip1(i_i2c_tx_fifo_data_buf[4]), .ip2(n9545), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .op(n5225) );
  nand2_1 U11487 ( .ip1(n9546), .ip2(i_i2c_U_dff_tx_mem[30]), .op(n9563) );
  inv_1 U11488 ( .ip(i_i2c_U_dff_tx_mem[3]), .op(n9547) );
  nor2_1 U11489 ( .ip1(n9548), .ip2(n9547), .op(n9558) );
  nand2_1 U11490 ( .ip1(n9549), .ip2(i_i2c_U_dff_tx_mem[12]), .op(n9556) );
  nand2_1 U11491 ( .ip1(n9550), .ip2(i_i2c_U_dff_tx_mem[21]), .op(n9555) );
  nand2_1 U11492 ( .ip1(n9551), .ip2(i_i2c_U_dff_tx_mem[48]), .op(n9554) );
  nand2_1 U11493 ( .ip1(n9552), .ip2(i_i2c_U_dff_tx_mem[66]), .op(n9553) );
  nand4_1 U11494 ( .ip1(n9556), .ip2(n9555), .ip3(n9554), .ip4(n9553), .op(
        n9557) );
  not_ab_or_c_or_d U11495 ( .ip1(n9559), .ip2(i_i2c_U_dff_tx_mem[57]), .ip3(
        n9558), .ip4(n9557), .op(n9562) );
  nand2_1 U11496 ( .ip1(n9560), .ip2(i_i2c_U_dff_tx_mem[39]), .op(n9561) );
  nand3_1 U11497 ( .ip1(n9563), .ip2(n9562), .ip3(n9561), .op(n9564) );
  mux2_1 U11498 ( .ip1(i_i2c_tx_fifo_data_buf[3]), .ip2(n9564), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .op(n5226) );
  inv_1 U11499 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[6]), .op(
        n11346) );
  inv_1 U11500 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[4]), .op(
        n11339) );
  inv_1 U11501 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[5]), .op(
        n11342) );
  inv_1 U11502 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[7]), .op(
        n11352) );
  nor4_1 U11503 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[1]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[2]), .ip3(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[3]), .ip4(n9571), .op(
        n9602) );
  inv_1 U11504 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[0]), .op(
        n11326) );
  and3_1 U11505 ( .ip1(n9638), .ip2(n9602), .ip3(n11326), .op(n9565) );
  and2_1 U11506 ( .ip1(n9565), .ip2(n11113), .op(n9567) );
  nand3_1 U11507 ( .ip1(n11115), .ip2(i_i2c_sda_vld), .ip3(n11113), .op(n11328) );
  mux2_1 U11508 ( .ip1(n9638), .ip2(i_i2c_rx_gen_call), .s(n9568), .op(n5091)
         );
  inv_1 U11509 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[3]), .op(
        n11336) );
  nor2_1 U11510 ( .ip1(n11336), .ip2(n9571), .op(n9634) );
  nand4_1 U11511 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[6]), 
        .ip2(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[4]), .ip3(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[5]), .ip4(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[7]), .op(n9572) );
  nor2_1 U11512 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[3]), .ip2(
        n9572), .op(n9620) );
  inv_1 U11513 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[1]), .op(
        n11330) );
  nor2_1 U11514 ( .ip1(n11330), .ip2(i_i2c_ic_sar[8]), .op(n9573) );
  not_ab_or_c_or_d U11515 ( .ip1(n11330), .ip2(i_i2c_ic_sar[8]), .ip3(n9573), 
        .ip4(i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_slv_1_sync_N2), .op(n9575) );
  inv_1 U11516 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[2]), .op(
        n11333) );
  mux2_1 U11517 ( .ip1(n11333), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[2]), .s(i_i2c_ic_sar[9]), 
        .op(n9574) );
  or2_1 U11518 ( .ip1(n9576), .ip2(n9647), .op(n9648) );
  or2_1 U11519 ( .ip1(n9577), .ip2(n9647), .op(n9578) );
  nand2_1 U11520 ( .ip1(n9648), .ip2(n9578), .op(n9599) );
  mux2_1 U11521 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[4]), .ip2(
        n11339), .s(i_i2c_ic_sar[4]), .op(n9582) );
  mux2_1 U11522 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[5]), .ip2(
        n11342), .s(i_i2c_ic_sar[5]), .op(n9581) );
  mux2_1 U11523 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[3]), .ip2(
        n11336), .s(i_i2c_ic_sar[3]), .op(n9580) );
  mux2_1 U11524 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[7]), .ip2(
        n11352), .s(i_i2c_ic_sar[7]), .op(n9579) );
  mux2_1 U11525 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[1]), .ip2(
        n11330), .s(i_i2c_ic_sar[1]), .op(n9584) );
  mux2_1 U11526 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[2]), .ip2(
        n11333), .s(i_i2c_ic_sar[2]), .op(n9583) );
  nand2_1 U11527 ( .ip1(n11301), .ip2(n9600), .op(n9607) );
  mux2_1 U11528 ( .ip1(n11326), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[0]), .s(i_i2c_ic_sar[0]), 
        .op(n9586) );
  mux2_1 U11529 ( .ip1(n11346), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[6]), .s(i_i2c_ic_sar[6]), 
        .op(n9585) );
  nand2_1 U11530 ( .ip1(n9589), .ip2(
        i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_slv_1_sync_N2), .op(n9617) );
  mux2_1 U11531 ( .ip1(n11346), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[6]), .s(i_i2c_ic_sar[5]), 
        .op(n9593) );
  mux2_1 U11532 ( .ip1(n11339), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[4]), .s(i_i2c_ic_sar[3]), 
        .op(n9592) );
  mux2_1 U11533 ( .ip1(n11333), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[2]), .s(i_i2c_ic_sar[1]), 
        .op(n9591) );
  mux2_1 U11534 ( .ip1(n11342), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[5]), .s(i_i2c_ic_sar[4]), 
        .op(n9590) );
  nand4_1 U11535 ( .ip1(n9593), .ip2(n9592), .ip3(n9591), .ip4(n9590), .op(
        n9594) );
  mux2_1 U11536 ( .ip1(n11330), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[1]), .s(i_i2c_ic_sar[0]), 
        .op(n9597) );
  mux2_1 U11537 ( .ip1(n11352), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[7]), .s(i_i2c_ic_sar[6]), 
        .op(n9596) );
  mux2_1 U11538 ( .ip1(n11336), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[3]), .s(i_i2c_ic_sar[2]), 
        .op(n9595) );
  nand2_1 U11539 ( .ip1(n9606), .ip2(n9623), .op(n9650) );
  not_ab_or_c_or_d U11540 ( .ip1(n9600), .ip2(n9570), .ip3(n9599), .ip4(n9650), 
        .op(n9601) );
  or2_1 U11541 ( .ip1(n9601), .ip2(n11721), .op(n9604) );
  nand4_1 U11542 ( .ip1(n9638), .ip2(n9602), .ip3(
        i_i2c_ic_ack_general_call_sync), .ip4(n11326), .op(n9603) );
  nand2_1 U11543 ( .ip1(n9604), .ip2(n9603), .op(n9611) );
  or2_1 U11544 ( .ip1(n11769), .ip2(n9606), .op(n9653) );
  nand3_1 U11545 ( .ip1(n11714), .ip2(n9608), .ip3(n9607), .op(n9609) );
  mux2_1 U11546 ( .ip1(i_i2c_slv_rx_ack_vld), .ip2(n9611), .s(n9610), .op(
        n5089) );
  nand3_1 U11547 ( .ip1(n11773), .ip2(i_i2c_mst_rx_bit_count[0]), .ip3(n9612), 
        .op(n9613) );
  nor3_1 U11548 ( .ip1(i_i2c_mst_rx_bit_count[2]), .ip2(n9642), .ip3(n9613), 
        .op(n11309) );
  mux2_1 U11549 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[4]), .ip2(
        i_i2c_sda_int), .s(n11309), .op(n4932) );
  nor2_1 U11550 ( .ip1(i_i2c_mst_rx_bit_count[2]), .ip2(n9632), .op(n9614) );
  mux2_1 U11551 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[6]), .ip2(
        i_i2c_sda_int), .s(n9614), .op(n4930) );
  inv_1 U11552 ( .ip(i_i2c_tx_wr_addr[1]), .op(n11253) );
  mux2_1 U11553 ( .ip1(i_i2c_U_dff_tx_mem[53]), .ip2(i_apb_pwdata_int[8]), .s(
        n9615), .op(n4966) );
  mux2_1 U11554 ( .ip1(i_i2c_U_dff_tx_mem[71]), .ip2(i_apb_pwdata_int[8]), .s(
        n9616), .op(n4964) );
  mux2_1 U11555 ( .ip1(i_i2c_U_dff_tx_mem[51]), .ip2(i_apb_pwdata_int[6]), .s(
        n9615), .op(n4982) );
  mux2_1 U11556 ( .ip1(i_i2c_U_dff_tx_mem[52]), .ip2(i_apb_pwdata_int[7]), .s(
        n9615), .op(n4974) );
  mux2_1 U11557 ( .ip1(i_i2c_U_dff_tx_mem[69]), .ip2(i_apb_pwdata_int[6]), .s(
        n9616), .op(n4980) );
  mux2_1 U11558 ( .ip1(i_i2c_U_dff_tx_mem[49]), .ip2(i_apb_pwdata_int[4]), .s(
        n9615), .op(n4998) );
  mux2_1 U11559 ( .ip1(i_i2c_U_dff_tx_mem[70]), .ip2(i_apb_pwdata_int[7]), .s(
        n9616), .op(n4972) );
  mux2_1 U11560 ( .ip1(i_i2c_U_dff_tx_mem[67]), .ip2(i_apb_pwdata_int[4]), .s(
        n9616), .op(n4996) );
  mux2_1 U11561 ( .ip1(i_i2c_U_dff_tx_mem[50]), .ip2(i_apb_pwdata_int[5]), .s(
        n9615), .op(n4990) );
  mux2_1 U11562 ( .ip1(i_i2c_U_dff_tx_mem[66]), .ip2(i_apb_pwdata_int[3]), .s(
        n9616), .op(n5004) );
  mux2_1 U11563 ( .ip1(i_i2c_U_dff_tx_mem[48]), .ip2(i_apb_pwdata_int[3]), .s(
        n9615), .op(n5006) );
  mux2_1 U11564 ( .ip1(i_i2c_U_dff_tx_mem[46]), .ip2(i_apb_pwdata_int[1]), .s(
        n9615), .op(n5022) );
  mux2_1 U11565 ( .ip1(i_i2c_U_dff_tx_mem[64]), .ip2(i_apb_pwdata_int[1]), .s(
        n9616), .op(n5020) );
  mux2_1 U11566 ( .ip1(i_i2c_U_dff_tx_mem[68]), .ip2(i_apb_pwdata_int[5]), .s(
        n9616), .op(n4988) );
  mux2_1 U11567 ( .ip1(i_i2c_U_dff_tx_mem[45]), .ip2(i_apb_pwdata_int[0]), .s(
        n9615), .op(n5030) );
  mux2_1 U11568 ( .ip1(i_i2c_U_dff_tx_mem[47]), .ip2(i_apb_pwdata_int[2]), .s(
        n9615), .op(n5014) );
  mux2_1 U11569 ( .ip1(i_i2c_U_dff_tx_mem[65]), .ip2(i_apb_pwdata_int[2]), .s(
        n9616), .op(n5012) );
  mux2_1 U11570 ( .ip1(i_i2c_U_dff_tx_mem[63]), .ip2(i_apb_pwdata_int[0]), .s(
        n9616), .op(n5028) );
  inv_1 U11571 ( .ip(n9617), .op(n9619) );
  inv_1 U11572 ( .ip(n9647), .op(n9618) );
  or2_1 U11573 ( .ip1(n9619), .ip2(n9618), .op(n9621) );
  nand2_1 U11574 ( .ip1(n9621), .ip2(n9620), .op(n9622) );
  inv_1 U11575 ( .ip(n9622), .op(n9626) );
  and2_1 U11576 ( .ip1(n9623), .ip2(n9622), .op(n9624) );
  mux2_1 U11577 ( .ip1(n9626), .ip2(i_i2c_rx_addr_10bit), .s(n9654), .op(n5093) );
  nor2_1 U11578 ( .ip1(n9628), .ip2(n9627), .op(n9630) );
  mux2_1 U11579 ( .ip1(n9631), .ip2(n9630), .s(n9629), .op(n4145) );
  mux2_1 U11580 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[2]), .ip2(
        i_i2c_sda_int), .s(n11310), .op(n4934) );
  mux2_1 U11581 ( .ip1(i_i2c_rx_hs_mcode), .ip2(n9638), .s(n9637), .op(n5090)
         );
  mux2_1 U11582 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[0]), .ip2(
        i_i2c_sda_int), .s(n9639), .op(n4936) );
  nor3_1 U11583 ( .ip1(i_i2c_mst_rx_bit_count[1]), .ip2(n9643), .ip3(n9645), 
        .op(n9640) );
  mux2_1 U11584 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[3]), .ip2(
        i_i2c_sda_int), .s(n9640), .op(n4933) );
  nor3_1 U11585 ( .ip1(i_i2c_mst_rx_bit_count[2]), .ip2(n9642), .ip3(n9645), 
        .op(n9641) );
  mux2_1 U11586 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[5]), .ip2(
        i_i2c_sda_int), .s(n9641), .op(n4931) );
  mux2_1 U11587 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[1]), .ip2(
        i_i2c_sda_int), .s(n9644), .op(n4935) );
  nor3_1 U11588 ( .ip1(i_i2c_mst_rx_bit_count[2]), .ip2(
        i_i2c_mst_rx_bit_count[1]), .ip3(n9645), .op(n9646) );
  mux2_1 U11589 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[7]), .ip2(
        i_i2c_sda_int), .s(n9646), .op(n4929) );
  or2_1 U11590 ( .ip1(i_i2c_rx_slv_read), .ip2(n9647), .op(n9649) );
  nand2_1 U11591 ( .ip1(n9649), .ip2(n9648), .op(n9651) );
  nor2_1 U11592 ( .ip1(n9651), .ip2(n9650), .op(n9652) );
  nor2_1 U11593 ( .ip1(n11721), .ip2(n9652), .op(n9656) );
  mux2_1 U11594 ( .ip1(i_i2c_rx_addr_match), .ip2(n9656), .s(n9655), .op(n5092) );
  xor2_1 U11595 ( .ip1(n9657), .ip2(i_i2c_rx_done_flg), .op(n5071) );
  nor3_1 U11596 ( .ip1(i_i2c_slv_ack_det), .ip2(n9658), .ip3(n5245), .op(n9659) );
  xor2_1 U11597 ( .ip1(n9659), .ip2(i_i2c_slv_clr_leftover_flg), .op(n5038) );
  xor2_1 U11598 ( .ip1(i_i2c_tx_pop_flg), .ip2(i_i2c_tx_pop), .op(n4180) );
  xor2_1 U11599 ( .ip1(i_i2c_p_det_flg), .ip2(i_i2c_p_det_intr), .op(n4169) );
  xor2_1 U11600 ( .ip1(i_i2c_rx_push_flg), .ip2(i_i2c_rx_push), .op(n4170) );
  xor2_1 U11601 ( .ip1(i_i2c_set_tx_empty_en_flg), .ip2(i_i2c_set_tx_empty_en), 
        .op(n4143) );
  mux2_1 U11602 ( .ip1(n11606), .ip2(i_ssi_prdata[25]), .s(n9660), .op(n4219)
         );
  mux2_1 U11603 ( .ip1(n11606), .ip2(i_ssi_prdata[29]), .s(n9660), .op(n4215)
         );
  mux2_1 U11604 ( .ip1(n11606), .ip2(i_ssi_prdata[28]), .s(n9660), .op(n4216)
         );
  mux2_1 U11605 ( .ip1(i_ssi_imr[3]), .ip2(i_apb_pwdata_int[3]), .s(n9917), 
        .op(n4647) );
  mux2_1 U11606 ( .ip1(i_ssi_imr[4]), .ip2(i_apb_pwdata_int[4]), .s(n9917), 
        .op(n4646) );
  mux2_1 U11607 ( .ip1(i_ssi_imr[1]), .ip2(i_apb_pwdata_int[1]), .s(n9917), 
        .op(n4649) );
  mux2_1 U11608 ( .ip1(i_ssi_imr[2]), .ip2(i_apb_pwdata_int[2]), .s(n9917), 
        .op(n4648) );
  mux2_1 U11609 ( .ip1(i_ssi_imr[0]), .ip2(i_apb_pwdata_int[0]), .s(n9917), 
        .op(n4650) );
  xor2_1 U11610 ( .ip1(n9661), .ip2(i_i2c_tx_abrt_source[5]), .op(n4940) );
  xor2_1 U11611 ( .ip1(i_i2c_tx_abrt_source[2]), .ip2(n9663), .op(n5188) );
  nor2_1 U11612 ( .ip1(n9667), .ip2(n9664), .op(n9665) );
  xor2_1 U11613 ( .ip1(i_i2c_tx_abrt_source[0]), .ip2(n9665), .op(n5194) );
  nor2_1 U11614 ( .ip1(n9667), .ip2(n9666), .op(n9668) );
  xor2_1 U11615 ( .ip1(i_i2c_tx_abrt_source[1]), .ip2(n9668), .op(n5192) );
  nor2_1 U11616 ( .ip1(n11760), .ip2(n11148), .op(n9670) );
  or4_1 U11617 ( .ip1(i_ssi_U_regfile_rxflr[0]), .ip2(i_ssi_U_regfile_rxflr[1]), .ip3(i_ssi_U_regfile_rxflr[2]), .ip4(i_ssi_U_regfile_rxflr[3]), .op(n9669)
         );
  nor2_1 U11618 ( .ip1(n9671), .ip2(n11165), .op(n11522) );
  inv_1 U11619 ( .ip(n11522), .op(n9674) );
  nor2_1 U11620 ( .ip1(i_ssi_U_regfile_rxflr[3]), .ip2(n11148), .op(n9672) );
  and2_1 U11621 ( .ip1(n11165), .ip2(n5453), .op(n9680) );
  inv_1 U11622 ( .ip(n9680), .op(n9673) );
  nor3_1 U11623 ( .ip1(n9680), .ip2(n11148), .ip3(n11522), .op(n9679) );
  inv_1 U11624 ( .ip(i_ssi_U_regfile_rxflr[1]), .op(n11531) );
  inv_1 U11625 ( .ip(i_ssi_U_regfile_rxflr[0]), .op(n11529) );
  nand2_1 U11626 ( .ip1(n9680), .ip2(n9676), .op(n11524) );
  nor2_1 U11627 ( .ip1(i_ssi_U_regfile_rxflr[1]), .ip2(
        i_ssi_U_regfile_rxflr[0]), .op(n9677) );
  nand2_1 U11628 ( .ip1(n11522), .ip2(n9677), .op(n11535) );
  nand2_1 U11629 ( .ip1(n11524), .ip2(n11535), .op(n9682) );
  nand2_1 U11630 ( .ip1(n11522), .ip2(i_ssi_U_regfile_rxflr[1]), .op(n9681) );
  nor2_1 U11631 ( .ip1(n9679), .ip2(n9678), .op(n11532) );
  nand2_1 U11632 ( .ip1(n9680), .ip2(n11531), .op(n11530) );
  nand3_1 U11633 ( .ip1(n9681), .ip2(n11532), .ip3(n11530), .op(n11526) );
  nand2_1 U11634 ( .ip1(n9687), .ip2(n9686), .op(n9688) );
  nand2_1 U11635 ( .ip1(n9689), .ip2(n9688), .op(n9690) );
  mux2_1 U11636 ( .ip1(n9691), .ip2(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[0]), .s(n10051), .op(n4394) );
  inv_1 U11637 ( .ip(i_ssi_tx_wr_addr[2]), .op(n10165) );
  inv_1 U11638 ( .ip(i_ssi_tx_wr_addr[1]), .op(n11212) );
  nand2_1 U11639 ( .ip1(n9692), .ip2(i_ssi_tx_full), .op(n9693) );
  inv_1 U11640 ( .ip(n9695), .op(n9694) );
  nor3_2 U11641 ( .ip1(n10165), .ip2(n11212), .ip3(n11211), .op(n10034) );
  nor2_1 U11642 ( .ip1(n11212), .ip2(n9695), .op(n11214) );
  inv_1 U11643 ( .ip(i_ssi_tx_wr_addr[0]), .op(n9698) );
  xor2_1 U11644 ( .ip1(i_i2c_tx_abrt_source[7]), .ip2(n9700), .op(n5187) );
  or2_1 U11645 ( .ip1(n10246), .ip2(n5279), .op(n9703) );
  nand2_1 U11646 ( .ip1(n10346), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[2]), 
        .op(n9702) );
  nand2_1 U11647 ( .ip1(n9714), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[1]), .op(n9701) );
  nand4_1 U11648 ( .ip1(n9703), .ip2(n9717), .ip3(n9702), .ip4(n9701), .op(
        n9706) );
  nor2_1 U11649 ( .ip1(n5334), .ip2(n9704), .op(n9705) );
  or2_1 U11650 ( .ip1(n9707), .ip2(n5279), .op(n9711) );
  nand2_1 U11651 ( .ip1(n9708), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[8]), 
        .op(n9710) );
  nand2_1 U11652 ( .ip1(n9714), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[7]), .op(n9709) );
  nand4_1 U11653 ( .ip1(n9711), .ip2(n9717), .ip3(n9710), .ip4(n9709), .op(
        n9713) );
  or2_1 U11654 ( .ip1(n10251), .ip2(n5279), .op(n9718) );
  nand2_1 U11655 ( .ip1(n10346), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[4]), 
        .op(n9716) );
  nand2_1 U11656 ( .ip1(n9714), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[3]), .op(n9715) );
  nand4_1 U11657 ( .ip1(n9718), .ip2(n9717), .ip3(n9716), .ip4(n9715), .op(
        n9719) );
  inv_1 U11658 ( .ip(i_i2c_ic_master), .op(
        i_i2c_U_DW_apb_i2c_sync_U_ic_master_1_sync_N2) );
  nor2_1 U11659 ( .ip1(i_ssi_U_regfile_ctrlr0_ir_int[5]), .ip2(
        i_ssi_U_regfile_ctrlr0_ir_int[4]), .op(n9720) );
  nand2_1 U11660 ( .ip1(n9720), .ip2(i_ssi_U_regfile_ctrlr0_ir_int_7), .op(
        n5242) );
  nor2_1 U11661 ( .ip1(i_ssi_U_fifo_U_tx_fifo_almost_empty_n), .ip2(n11148), 
        .op(i_ssi_U_intctl_N2) );
  mux2_1 U11662 ( .ip1(i_i2c_s_det), .ip2(n10801), .s(i_i2c_s_det_flg), .op(
        n4178) );
  inv_1 U11663 ( .ip(n9721), .op(n9722) );
  nand2_1 U11664 ( .ip1(n9726), .ip2(n9725), .op(i_i2c_U_DW_apb_i2c_toggle_N32) );
  nand2_1 U11665 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv), .ip2(
        n9727), .op(n9728) );
  xnor2_1 U11666 ( .ip1(i_i2c_tx_abrt_source[11]), .ip2(n9728), .op(n4862) );
  nor2_1 U11667 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[0]), 
        .ip2(n10561), .op(i_i2c_U_DW_apb_i2c_rx_filter_N82) );
  inv_1 U11668 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt[0]), .op(n9729) );
  nor2_1 U11669 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt[1]), .ip2(n9729), 
        .op(n9730) );
  nor2_1 U11670 ( .ip1(n9730), .ip2(n10584), .op(n5094) );
  nor2_1 U11671 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt[1]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt[0]), .op(n9731) );
  nor2_1 U11672 ( .ip1(n9731), .ip2(n10584), .op(n5095) );
  mux2_1 U11673 ( .ip1(i_i2c_prdata[24]), .ip2(i_i2c_iprdata[24]), .s(n11762), 
        .op(n4685) );
  inv_1 U11674 ( .ip(n9732), .op(n9733) );
  mux2_1 U11675 ( .ip1(n9733), .ip2(n9732), .s(i_i2c_ic_rd_req_flg), .op(n5037) );
  mux2_1 U11676 ( .ip1(i_i2c_prdata[18]), .ip2(i_i2c_iprdata[18]), .s(n11762), 
        .op(n4679) );
  mux2_1 U11677 ( .ip1(i_i2c_prdata[22]), .ip2(i_i2c_iprdata[22]), .s(n11762), 
        .op(n4683) );
  mux2_1 U11678 ( .ip1(i_i2c_prdata[21]), .ip2(i_i2c_iprdata[21]), .s(n11762), 
        .op(n4682) );
  mux2_1 U11679 ( .ip1(i_i2c_prdata[23]), .ip2(i_i2c_iprdata[23]), .s(n11762), 
        .op(n4684) );
  inv_1 U11680 ( .ip(i_i2c_ic_clk_in_a), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_U_SYNC_N2) );
  nand2_1 U11681 ( .ip1(n9735), .ip2(i_i2c_ic_tar[0]), .op(n9736) );
  not_ab_or_c_or_d U11682 ( .ip1(n9740), .ip2(i_i2c_ic_hs_maddr[0]), .ip3(
        n9739), .ip4(n9738), .op(n9741) );
  nand2_1 U11683 ( .ip1(n9742), .ip2(n9741), .op(n9744) );
  mux2_1 U11684 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[0]), .ip2(
        n9744), .s(n9743), .op(n5047) );
  nand2_1 U11685 ( .ip1(i_i2c_rx_wr_addr[1]), .ip2(i_i2c_rx_wr_addr[2]), .op(
        n9746) );
  or2_1 U11686 ( .ip1(i_i2c_rx_wr_addr[0]), .ip2(n11197), .op(n9769) );
  mux2_1 U11687 ( .ip1(i_i2c_U_dff_rx_mem[11]), .ip2(i_i2c_rx_push_data[3]), 
        .s(n9745), .op(n4903) );
  mux2_1 U11688 ( .ip1(i_i2c_U_dff_rx_mem[15]), .ip2(i_i2c_rx_push_data[7]), 
        .s(n9745), .op(n4871) );
  mux2_1 U11689 ( .ip1(i_i2c_U_dff_rx_mem[9]), .ip2(i_i2c_rx_push_data[1]), 
        .s(n9745), .op(n4919) );
  mux2_1 U11690 ( .ip1(i_i2c_U_dff_rx_mem[14]), .ip2(i_i2c_rx_push_data[6]), 
        .s(n9745), .op(n4879) );
  mux2_1 U11691 ( .ip1(i_i2c_U_dff_rx_mem[10]), .ip2(i_i2c_rx_push_data[2]), 
        .s(n9745), .op(n4911) );
  mux2_1 U11692 ( .ip1(i_i2c_U_dff_rx_mem[12]), .ip2(i_i2c_rx_push_data[4]), 
        .s(n9745), .op(n4895) );
  mux2_1 U11693 ( .ip1(i_i2c_U_dff_rx_mem[13]), .ip2(i_i2c_rx_push_data[5]), 
        .s(n9745), .op(n4887) );
  mux2_1 U11694 ( .ip1(i_i2c_U_dff_rx_mem[8]), .ip2(i_i2c_rx_push_data[0]), 
        .s(n9745), .op(n4927) );
  mux2_1 U11695 ( .ip1(i_i2c_U_dff_rx_mem[6]), .ip2(i_i2c_rx_push_data[6]), 
        .s(n9747), .op(n4880) );
  mux2_1 U11696 ( .ip1(i_i2c_U_dff_rx_mem[0]), .ip2(i_i2c_rx_push_data[0]), 
        .s(n9747), .op(n4928) );
  mux2_1 U11697 ( .ip1(i_i2c_U_dff_rx_mem[4]), .ip2(i_i2c_rx_push_data[4]), 
        .s(n9747), .op(n4896) );
  mux2_1 U11698 ( .ip1(i_i2c_U_dff_rx_mem[3]), .ip2(i_i2c_rx_push_data[3]), 
        .s(n9747), .op(n4904) );
  mux2_1 U11699 ( .ip1(i_i2c_U_dff_rx_mem[1]), .ip2(i_i2c_rx_push_data[1]), 
        .s(n9747), .op(n4920) );
  mux2_1 U11700 ( .ip1(i_i2c_U_dff_rx_mem[7]), .ip2(i_i2c_rx_push_data[7]), 
        .s(n9747), .op(n4872) );
  mux2_1 U11701 ( .ip1(i_i2c_U_dff_rx_mem[5]), .ip2(i_i2c_rx_push_data[5]), 
        .s(n9747), .op(n4888) );
  mux2_1 U11702 ( .ip1(i_i2c_U_dff_rx_mem[2]), .ip2(i_i2c_rx_push_data[2]), 
        .s(n9747), .op(n4912) );
  nor2_1 U11703 ( .ip1(i_i2c_tx_wr_addr[0]), .ip2(n9783), .op(n9748) );
  nand3_1 U11704 ( .ip1(i_i2c_tx_wr_addr[2]), .ip2(n9748), .ip3(n11253), .op(
        n9749) );
  mux2_1 U11705 ( .ip1(i_apb_pwdata_int[8]), .ip2(i_i2c_U_dff_tx_mem[35]), .s(
        n9749), .op(n4968) );
  mux2_1 U11706 ( .ip1(i_apb_pwdata_int[7]), .ip2(i_i2c_U_dff_tx_mem[34]), .s(
        n9749), .op(n4976) );
  mux2_1 U11707 ( .ip1(i_apb_pwdata_int[3]), .ip2(i_i2c_U_dff_tx_mem[30]), .s(
        n9749), .op(n5008) );
  mux2_1 U11708 ( .ip1(i_apb_pwdata_int[6]), .ip2(i_i2c_U_dff_tx_mem[33]), .s(
        n9749), .op(n4984) );
  mux2_1 U11709 ( .ip1(i_apb_pwdata_int[4]), .ip2(i_i2c_U_dff_tx_mem[31]), .s(
        n9749), .op(n5000) );
  mux2_1 U11710 ( .ip1(i_apb_pwdata_int[1]), .ip2(i_i2c_U_dff_tx_mem[28]), .s(
        n9749), .op(n5024) );
  mux2_1 U11711 ( .ip1(i_apb_pwdata_int[5]), .ip2(i_i2c_U_dff_tx_mem[32]), .s(
        n9749), .op(n4992) );
  mux2_1 U11712 ( .ip1(i_apb_pwdata_int[0]), .ip2(i_i2c_U_dff_tx_mem[27]), .s(
        n9749), .op(n5032) );
  mux2_1 U11713 ( .ip1(i_apb_pwdata_int[2]), .ip2(i_i2c_U_dff_tx_mem[29]), .s(
        n9749), .op(n5016) );
  inv_1 U11714 ( .ip(n9754), .op(n9756) );
  or4_1 U11715 ( .ip1(n9758), .ip2(n9757), .ip3(n9756), .ip4(n9755), .op(n9759) );
  not_ab_or_c_or_d U11716 ( .ip1(i_i2c_ic_sda_rx_hold_sync[0]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[0]), .ip3(n9760), 
        .ip4(n9759), .op(n9761) );
  nand2_1 U11717 ( .ip1(n9762), .ip2(n9761), .op(n9763) );
  nand2_1 U11718 ( .ip1(n11776), .ip2(n9763), .op(n9764) );
  mux2_1 U11719 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_sda_post_hold_done), .ip2(
        n9765), .s(n9764), .op(n5104) );
  nand2_1 U11720 ( .ip1(i_i2c_tx_wr_addr[0]), .ip2(n9766), .op(n11252) );
  mux2_1 U11721 ( .ip1(i_i2c_U_dff_tx_mem[8]), .ip2(i_apb_pwdata_int[8]), .s(
        n11255), .op(n4971) );
  mux2_1 U11722 ( .ip1(i_i2c_U_dff_tx_mem[6]), .ip2(i_apb_pwdata_int[6]), .s(
        n11255), .op(n4987) );
  mux2_1 U11723 ( .ip1(i_i2c_U_dff_tx_mem[3]), .ip2(i_apb_pwdata_int[3]), .s(
        n11255), .op(n5011) );
  mux2_1 U11724 ( .ip1(i_i2c_U_dff_tx_mem[7]), .ip2(i_apb_pwdata_int[7]), .s(
        n11255), .op(n4979) );
  mux2_1 U11725 ( .ip1(i_i2c_U_dff_tx_mem[1]), .ip2(i_apb_pwdata_int[1]), .s(
        n11255), .op(n5027) );
  mux2_1 U11726 ( .ip1(i_i2c_U_dff_tx_mem[5]), .ip2(i_apb_pwdata_int[5]), .s(
        n11255), .op(n4995) );
  mux2_1 U11727 ( .ip1(i_i2c_U_dff_tx_mem[4]), .ip2(i_apb_pwdata_int[4]), .s(
        n11255), .op(n5003) );
  mux2_1 U11728 ( .ip1(i_i2c_U_dff_tx_mem[0]), .ip2(i_apb_pwdata_int[0]), .s(
        n11255), .op(n5035) );
  mux2_1 U11729 ( .ip1(i_i2c_U_dff_tx_mem[2]), .ip2(i_apb_pwdata_int[2]), .s(
        n11255), .op(n5019) );
  nor3_1 U11730 ( .ip1(i_i2c_rx_wr_addr[1]), .ip2(n9767), .ip3(n9769), .op(
        n9768) );
  mux2_1 U11731 ( .ip1(i_i2c_U_dff_rx_mem[26]), .ip2(i_i2c_rx_push_data[2]), 
        .s(n9768), .op(n4909) );
  mux2_1 U11732 ( .ip1(i_i2c_U_dff_rx_mem[24]), .ip2(i_i2c_rx_push_data[0]), 
        .s(n9768), .op(n4925) );
  mux2_1 U11733 ( .ip1(i_i2c_U_dff_rx_mem[30]), .ip2(i_i2c_rx_push_data[6]), 
        .s(n9768), .op(n4877) );
  mux2_1 U11734 ( .ip1(i_i2c_U_dff_rx_mem[28]), .ip2(i_i2c_rx_push_data[4]), 
        .s(n9768), .op(n4893) );
  mux2_1 U11735 ( .ip1(i_i2c_U_dff_rx_mem[25]), .ip2(i_i2c_rx_push_data[1]), 
        .s(n9768), .op(n4917) );
  mux2_1 U11736 ( .ip1(i_i2c_U_dff_rx_mem[27]), .ip2(i_i2c_rx_push_data[3]), 
        .s(n9768), .op(n4901) );
  mux2_1 U11737 ( .ip1(i_i2c_U_dff_rx_mem[29]), .ip2(i_i2c_rx_push_data[5]), 
        .s(n9768), .op(n4885) );
  mux2_1 U11738 ( .ip1(i_i2c_U_dff_rx_mem[31]), .ip2(i_i2c_rx_push_data[7]), 
        .s(n9768), .op(n4869) );
  nor3_1 U11739 ( .ip1(i_i2c_rx_wr_addr[1]), .ip2(i_i2c_rx_wr_addr[2]), .ip3(
        n9769), .op(n9771) );
  mux2_1 U11740 ( .ip1(i_i2c_U_dff_rx_mem[57]), .ip2(i_i2c_rx_push_data[1]), 
        .s(n9771), .op(n4913) );
  mux2_1 U11741 ( .ip1(i_i2c_U_dff_rx_mem[58]), .ip2(i_i2c_rx_push_data[2]), 
        .s(n9771), .op(n4905) );
  mux2_1 U11742 ( .ip1(i_i2c_U_dff_rx_mem[60]), .ip2(i_i2c_rx_push_data[4]), 
        .s(n9771), .op(n4889) );
  inv_1 U11743 ( .ip(i_i2c_rx_wr_addr[1]), .op(n11193) );
  nor3_1 U11744 ( .ip1(i_i2c_rx_wr_addr[2]), .ip2(n11193), .ip3(n9769), .op(
        n9770) );
  mux2_1 U11745 ( .ip1(i_i2c_U_dff_rx_mem[44]), .ip2(i_i2c_rx_push_data[4]), 
        .s(n9770), .op(n4891) );
  mux2_1 U11746 ( .ip1(i_i2c_U_dff_rx_mem[46]), .ip2(i_i2c_rx_push_data[6]), 
        .s(n9770), .op(n4875) );
  mux2_1 U11747 ( .ip1(i_i2c_U_dff_rx_mem[56]), .ip2(i_i2c_rx_push_data[0]), 
        .s(n9771), .op(n4921) );
  mux2_1 U11748 ( .ip1(i_i2c_U_dff_rx_mem[41]), .ip2(i_i2c_rx_push_data[1]), 
        .s(n9770), .op(n4915) );
  mux2_1 U11749 ( .ip1(i_i2c_U_dff_rx_mem[45]), .ip2(i_i2c_rx_push_data[5]), 
        .s(n9770), .op(n4883) );
  mux2_1 U11750 ( .ip1(i_i2c_U_dff_rx_mem[40]), .ip2(i_i2c_rx_push_data[0]), 
        .s(n9770), .op(n4923) );
  mux2_1 U11751 ( .ip1(i_i2c_U_dff_rx_mem[59]), .ip2(i_i2c_rx_push_data[3]), 
        .s(n9771), .op(n4897) );
  mux2_1 U11752 ( .ip1(i_i2c_U_dff_rx_mem[42]), .ip2(i_i2c_rx_push_data[2]), 
        .s(n9770), .op(n4907) );
  mux2_1 U11753 ( .ip1(i_i2c_U_dff_rx_mem[47]), .ip2(i_i2c_rx_push_data[7]), 
        .s(n9770), .op(n4867) );
  mux2_1 U11754 ( .ip1(i_i2c_U_dff_rx_mem[61]), .ip2(i_i2c_rx_push_data[5]), 
        .s(n9771), .op(n4881) );
  mux2_1 U11755 ( .ip1(i_i2c_U_dff_rx_mem[63]), .ip2(i_i2c_rx_push_data[7]), 
        .s(n9771), .op(n4865) );
  mux2_1 U11756 ( .ip1(i_i2c_U_dff_rx_mem[43]), .ip2(i_i2c_rx_push_data[3]), 
        .s(n9770), .op(n4899) );
  mux2_1 U11757 ( .ip1(i_i2c_U_dff_rx_mem[62]), .ip2(i_i2c_rx_push_data[6]), 
        .s(n9771), .op(n4873) );
  inv_1 U11758 ( .ip(i_i2c_rx_hs_mcode), .op(n9772) );
  nand3_1 U11759 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_rx_hs_mcode_r), .ip3(n9772), .op(n9776)
         );
  inv_1 U11760 ( .ip(i_i2c_hs_mcode_en), .op(n9774) );
  nand3_1 U11761 ( .ip1(n9774), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_hs_mcode_en_r), .ip3(n9773), .op(n9775)
         );
  nand2_1 U11762 ( .ip1(n9776), .ip2(n9775), .op(n9778) );
  mux2_1 U11763 ( .ip1(n9778), .ip2(n9777), .s(
        i_i2c_U_DW_apb_i2c_rx_filter_hs_mcode_fed_dtctd_r), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_N50) );
  nor3_1 U11764 ( .ip1(i_i2c_rx_wr_addr[2]), .ip2(n11193), .ip3(n11194), .op(
        n9780) );
  mux2_1 U11765 ( .ip1(i_i2c_U_dff_rx_mem[36]), .ip2(i_i2c_rx_push_data[4]), 
        .s(n9780), .op(n4892) );
  mux2_1 U11766 ( .ip1(i_i2c_U_dff_rx_mem[39]), .ip2(i_i2c_rx_push_data[7]), 
        .s(n9780), .op(n4868) );
  mux2_1 U11767 ( .ip1(i_i2c_U_dff_rx_mem[37]), .ip2(i_i2c_rx_push_data[5]), 
        .s(n9780), .op(n4884) );
  nor3_1 U11768 ( .ip1(i_i2c_rx_wr_addr[1]), .ip2(i_i2c_rx_wr_addr[2]), .ip3(
        n11194), .op(n9779) );
  mux2_1 U11769 ( .ip1(i_i2c_U_dff_rx_mem[49]), .ip2(i_i2c_rx_push_data[1]), 
        .s(n9779), .op(n4914) );
  mux2_1 U11770 ( .ip1(i_i2c_U_dff_rx_mem[32]), .ip2(i_i2c_rx_push_data[0]), 
        .s(n9780), .op(n4924) );
  mux2_1 U11771 ( .ip1(i_i2c_U_dff_rx_mem[52]), .ip2(i_i2c_rx_push_data[4]), 
        .s(n9779), .op(n4890) );
  mux2_1 U11772 ( .ip1(i_i2c_U_dff_rx_mem[51]), .ip2(i_i2c_rx_push_data[3]), 
        .s(n9779), .op(n4898) );
  mux2_1 U11773 ( .ip1(i_i2c_U_dff_rx_mem[50]), .ip2(i_i2c_rx_push_data[2]), 
        .s(n9779), .op(n4906) );
  mux2_1 U11774 ( .ip1(i_i2c_U_dff_rx_mem[38]), .ip2(i_i2c_rx_push_data[6]), 
        .s(n9780), .op(n4876) );
  mux2_1 U11775 ( .ip1(i_i2c_U_dff_rx_mem[48]), .ip2(i_i2c_rx_push_data[0]), 
        .s(n9779), .op(n4922) );
  mux2_1 U11776 ( .ip1(i_i2c_U_dff_rx_mem[55]), .ip2(i_i2c_rx_push_data[7]), 
        .s(n9779), .op(n4866) );
  mux2_1 U11777 ( .ip1(i_i2c_U_dff_rx_mem[53]), .ip2(i_i2c_rx_push_data[5]), 
        .s(n9779), .op(n4882) );
  mux2_1 U11778 ( .ip1(i_i2c_U_dff_rx_mem[33]), .ip2(i_i2c_rx_push_data[1]), 
        .s(n9780), .op(n4916) );
  mux2_1 U11779 ( .ip1(i_i2c_U_dff_rx_mem[34]), .ip2(i_i2c_rx_push_data[2]), 
        .s(n9780), .op(n4908) );
  mux2_1 U11780 ( .ip1(i_i2c_U_dff_rx_mem[54]), .ip2(i_i2c_rx_push_data[6]), 
        .s(n9779), .op(n4874) );
  mux2_1 U11781 ( .ip1(i_i2c_U_dff_rx_mem[35]), .ip2(i_i2c_rx_push_data[3]), 
        .s(n9780), .op(n4900) );
  nor2_1 U11782 ( .ip1(i_i2c_tx_wr_addr[2]), .ip2(n11256), .op(n9781) );
  mux2_1 U11783 ( .ip1(i_i2c_U_dff_tx_mem[44]), .ip2(i_apb_pwdata_int[8]), .s(
        n9781), .op(n4967) );
  mux2_1 U11784 ( .ip1(i_i2c_U_dff_tx_mem[42]), .ip2(i_apb_pwdata_int[6]), .s(
        n9781), .op(n4983) );
  mux2_1 U11785 ( .ip1(i_i2c_U_dff_tx_mem[43]), .ip2(i_apb_pwdata_int[7]), .s(
        n9781), .op(n4975) );
  mux2_1 U11786 ( .ip1(i_i2c_U_dff_tx_mem[41]), .ip2(i_apb_pwdata_int[5]), .s(
        n9781), .op(n4991) );
  mux2_1 U11787 ( .ip1(i_i2c_U_dff_tx_mem[40]), .ip2(i_apb_pwdata_int[4]), .s(
        n9781), .op(n4999) );
  mux2_1 U11788 ( .ip1(i_i2c_U_dff_tx_mem[39]), .ip2(i_apb_pwdata_int[3]), .s(
        n9781), .op(n5007) );
  mux2_1 U11789 ( .ip1(i_i2c_U_dff_tx_mem[37]), .ip2(i_apb_pwdata_int[1]), .s(
        n9781), .op(n5023) );
  mux2_1 U11790 ( .ip1(i_i2c_U_dff_tx_mem[36]), .ip2(i_apb_pwdata_int[0]), .s(
        n9781), .op(n5031) );
  mux2_1 U11791 ( .ip1(i_i2c_U_dff_tx_mem[38]), .ip2(i_apb_pwdata_int[2]), .s(
        n9781), .op(n5015) );
  nor3_1 U11792 ( .ip1(i_i2c_tx_wr_addr[0]), .ip2(n9783), .ip3(n9782), .op(
        n9784) );
  mux2_1 U11793 ( .ip1(i_i2c_U_dff_tx_mem[12]), .ip2(i_apb_pwdata_int[3]), .s(
        n9784), .op(n5010) );
  mux2_1 U11794 ( .ip1(i_i2c_U_dff_tx_mem[10]), .ip2(i_apb_pwdata_int[1]), .s(
        n9784), .op(n5026) );
  mux2_1 U11795 ( .ip1(i_i2c_U_dff_tx_mem[15]), .ip2(i_apb_pwdata_int[6]), .s(
        n9784), .op(n4986) );
  mux2_1 U11796 ( .ip1(i_i2c_U_dff_tx_mem[11]), .ip2(i_apb_pwdata_int[2]), .s(
        n9784), .op(n5018) );
  mux2_1 U11797 ( .ip1(i_i2c_U_dff_tx_mem[14]), .ip2(i_apb_pwdata_int[5]), .s(
        n9784), .op(n4994) );
  mux2_1 U11798 ( .ip1(i_i2c_U_dff_tx_mem[13]), .ip2(i_apb_pwdata_int[4]), .s(
        n9784), .op(n5002) );
  mux2_1 U11799 ( .ip1(i_i2c_U_dff_tx_mem[17]), .ip2(i_apb_pwdata_int[8]), .s(
        n9784), .op(n4970) );
  mux2_1 U11800 ( .ip1(i_i2c_U_dff_tx_mem[16]), .ip2(i_apb_pwdata_int[7]), .s(
        n9784), .op(n4978) );
  mux2_1 U11801 ( .ip1(i_i2c_U_dff_tx_mem[9]), .ip2(i_apb_pwdata_int[0]), .s(
        n9784), .op(n5034) );
  nor2_1 U11802 ( .ip1(n9786), .ip2(n9785), .op(n11563) );
  nand2_1 U11803 ( .ip1(n9838), .ip2(n11563), .op(n9787) );
  mux2_1 U11804 ( .ip1(i_apb_pwdata_int[0]), .ip2(i_ssi_ser_0_), .s(n9787), 
        .op(n4634) );
  inv_1 U11805 ( .ip(n11599), .op(n9790) );
  nor2_1 U11806 ( .ip1(i_ssi_U_regfile_rxflr[3]), .ip2(n9790), .op(n9789) );
  or2_1 U11807 ( .ip1(n9790), .ip2(n9789), .op(n9798) );
  nand2_1 U11808 ( .ip1(n10310), .ip2(n11691), .op(n9793) );
  nand2_1 U11809 ( .ip1(i_ssi_U_regfile_ctrlr1_int[3]), .ip2(n11693), .op(
        n9792) );
  nand2_1 U11810 ( .ip1(n5358), .ip2(n11692), .op(n9791) );
  nand4_1 U11811 ( .ip1(n9793), .ip2(n9855), .ip3(n9792), .ip4(n9791), .op(
        n9795) );
  inv_1 U11812 ( .ip(i_ssi_U_fifo_U_rx_fifo_empty_n), .op(n9904) );
  nand2_1 U11813 ( .ip1(n9904), .ip2(n11576), .op(n9794) );
  nand2_1 U11814 ( .ip1(n9795), .ip2(n9794), .op(n9796) );
  mux2_1 U11815 ( .ip1(n11518), .ip2(n9796), .s(n9846), .op(n9797) );
  nand2_1 U11816 ( .ip1(n9798), .ip2(n9797), .op(n9813) );
  nand2_1 U11817 ( .ip1(n11677), .ip2(i_ssi_U_dff_rx_mem[51]), .op(n9802) );
  nand2_1 U11818 ( .ip1(n11674), .ip2(i_ssi_U_dff_rx_mem[115]), .op(n9801) );
  nand2_1 U11819 ( .ip1(n11686), .ip2(i_ssi_U_dff_rx_mem[67]), .op(n9800) );
  nand2_1 U11820 ( .ip1(n11679), .ip2(i_ssi_U_dff_rx_mem[35]), .op(n9799) );
  nand4_1 U11821 ( .ip1(n9802), .ip2(n9801), .ip3(n9800), .ip4(n9799), .op(
        n9808) );
  nand2_1 U11822 ( .ip1(n11676), .ip2(i_ssi_U_dff_rx_mem[19]), .op(n9806) );
  nand2_1 U11823 ( .ip1(n11687), .ip2(i_ssi_U_dff_rx_mem[99]), .op(n9805) );
  nand2_1 U11824 ( .ip1(n11678), .ip2(i_ssi_U_dff_rx_mem[83]), .op(n9804) );
  nand2_1 U11825 ( .ip1(n11675), .ip2(i_ssi_U_dff_rx_mem[3]), .op(n9803) );
  nand4_1 U11826 ( .ip1(n9806), .ip2(n9805), .ip3(n9804), .ip4(n9803), .op(
        n9807) );
  nor2_1 U11827 ( .ip1(n9808), .ip2(n9807), .op(n9809) );
  inv_1 U11828 ( .ip(n11598), .op(n9887) );
  nor2_1 U11829 ( .ip1(n9809), .ip2(n9887), .op(n9811) );
  nor2_1 U11830 ( .ip1(n11584), .ip2(i_ssi_ssi_rxo_intr_n), .op(n9810) );
  ab_or_c_or_d U11831 ( .ip1(i_ssi_risr[3]), .ip2(n11587), .ip3(n9811), .ip4(
        n9810), .op(n9812) );
  not_ab_or_c_or_d U11832 ( .ip1(i_ssi_imr[3]), .ip2(n11600), .ip3(n9813), 
        .ip4(n9812), .op(n9815) );
  nand2_1 U11833 ( .ip1(n9815), .ip2(n9814), .op(n9816) );
  mux2_1 U11834 ( .ip1(i_ssi_prdata[3]), .ip2(n9816), .s(n9832), .op(n4241) );
  mux2_1 U11835 ( .ip1(i_apb_pwdata_int[2]), .ip2(i_ssi_mwcr[2]), .s(n9817), 
        .op(n4635) );
  mux2_1 U11836 ( .ip1(i_apb_pwdata_int[12]), .ip2(i_ssi_cfs[0]), .s(n9837), 
        .op(n4599) );
  mux2_1 U11837 ( .ip1(i_apb_pwdata_int[13]), .ip2(i_ssi_cfs[1]), .s(n9837), 
        .op(n4600) );
  mux2_1 U11838 ( .ip1(i_apb_pwdata_int[10]), .ip2(i_ssi_ctrlr0[10]), .s(n9837), .op(n4597) );
  mux2_1 U11839 ( .ip1(i_apb_pwdata_int[15]), .ip2(i_ssi_cfs[3]), .s(n9837), 
        .op(n4602) );
  inv_1 U11840 ( .ip(i_i2c_tx_wr_addr[2]), .op(n11257) );
  nor3_1 U11841 ( .ip1(i_i2c_tx_wr_addr[1]), .ip2(n11257), .ip3(n11252), .op(
        n9818) );
  mux2_1 U11842 ( .ip1(i_i2c_U_dff_tx_mem[24]), .ip2(i_apb_pwdata_int[6]), .s(
        n9818), .op(n4985) );
  mux2_1 U11843 ( .ip1(i_i2c_U_dff_tx_mem[26]), .ip2(i_apb_pwdata_int[8]), .s(
        n9818), .op(n4969) );
  mux2_1 U11844 ( .ip1(i_i2c_U_dff_tx_mem[22]), .ip2(i_apb_pwdata_int[4]), .s(
        n9818), .op(n5001) );
  mux2_1 U11845 ( .ip1(i_i2c_U_dff_tx_mem[18]), .ip2(i_apb_pwdata_int[0]), .s(
        n9818), .op(n5033) );
  mux2_1 U11846 ( .ip1(i_i2c_U_dff_tx_mem[25]), .ip2(i_apb_pwdata_int[7]), .s(
        n9818), .op(n4977) );
  mux2_1 U11847 ( .ip1(i_i2c_U_dff_tx_mem[20]), .ip2(i_apb_pwdata_int[2]), .s(
        n9818), .op(n5017) );
  mux2_1 U11848 ( .ip1(i_i2c_U_dff_tx_mem[19]), .ip2(i_apb_pwdata_int[1]), .s(
        n9818), .op(n5025) );
  mux2_1 U11849 ( .ip1(i_i2c_U_dff_tx_mem[21]), .ip2(i_apb_pwdata_int[3]), .s(
        n9818), .op(n5009) );
  mux2_1 U11850 ( .ip1(i_i2c_U_dff_tx_mem[23]), .ip2(i_apb_pwdata_int[5]), .s(
        n9818), .op(n4993) );
  nor3_1 U11851 ( .ip1(i_i2c_tx_wr_addr[2]), .ip2(i_i2c_tx_wr_addr[1]), .ip3(
        n11252), .op(n9819) );
  mux2_1 U11852 ( .ip1(i_i2c_U_dff_tx_mem[57]), .ip2(i_apb_pwdata_int[3]), .s(
        n9819), .op(n5005) );
  mux2_1 U11853 ( .ip1(i_i2c_U_dff_tx_mem[61]), .ip2(i_apb_pwdata_int[7]), .s(
        n9819), .op(n4973) );
  mux2_1 U11854 ( .ip1(i_i2c_U_dff_tx_mem[58]), .ip2(i_apb_pwdata_int[4]), .s(
        n9819), .op(n4997) );
  mux2_1 U11855 ( .ip1(i_i2c_U_dff_tx_mem[55]), .ip2(i_apb_pwdata_int[1]), .s(
        n9819), .op(n5021) );
  mux2_1 U11856 ( .ip1(i_i2c_U_dff_tx_mem[62]), .ip2(i_apb_pwdata_int[8]), .s(
        n9819), .op(n4965) );
  mux2_1 U11857 ( .ip1(i_i2c_U_dff_tx_mem[59]), .ip2(i_apb_pwdata_int[5]), .s(
        n9819), .op(n4989) );
  mux2_1 U11858 ( .ip1(i_i2c_U_dff_tx_mem[56]), .ip2(i_apb_pwdata_int[2]), .s(
        n9819), .op(n5013) );
  mux2_1 U11859 ( .ip1(i_i2c_U_dff_tx_mem[60]), .ip2(i_apb_pwdata_int[6]), .s(
        n9819), .op(n4981) );
  mux2_1 U11860 ( .ip1(i_i2c_U_dff_tx_mem[54]), .ip2(i_apb_pwdata_int[0]), .s(
        n9819), .op(n5029) );
  or2_1 U11861 ( .ip1(n11616), .ip2(n11615), .op(n9821) );
  or3_1 U11862 ( .ip1(n9909), .ip2(i_ssi_reg_addr[0]), .ip3(i_ssi_reg_addr[2]), 
        .op(n9902) );
  nor2_1 U11863 ( .ip1(n9820), .ip2(n9902), .op(n11620) );
  inv_1 U11864 ( .ip(n11620), .op(n9830) );
  nand2_1 U11865 ( .ip1(n9821), .ip2(n9830), .op(n9822) );
  nand2_1 U11866 ( .ip1(n9822), .ip2(n9832), .op(n9823) );
  nand2_1 U11867 ( .ip1(n9823), .ip2(i_ssi_risr[3]), .op(n9826) );
  inv_1 U11868 ( .ip(i_ssi_U_fifo_rx_pop_dly), .op(n9824) );
  nand3_1 U11869 ( .ip1(i_ssi_U_fifo_rx_error_ir), .ip2(
        i_ssi_U_fifo_rx_push_sync_dly), .ip3(n9824), .op(n9825) );
  nand2_1 U11870 ( .ip1(n9826), .ip2(n9825), .op(n9827) );
  and2_1 U11871 ( .ip1(n9827), .ip2(n11569), .op(n4450) );
  nand2_1 U11872 ( .ip1(i_ssi_U_fifo_tx_error_ir), .ip2(
        i_ssi_U_fifo_tx_push_dly), .op(n9828) );
  nor2_1 U11873 ( .ip1(i_ssi_U_fifo_tx_pop_sync_dly), .ip2(n9828), .op(n9835)
         );
  or2_1 U11874 ( .ip1(n11616), .ip2(n9829), .op(n11562) );
  nand2_1 U11875 ( .ip1(n9830), .ip2(n11562), .op(n9831) );
  nand2_1 U11876 ( .ip1(n9832), .ip2(n9831), .op(n9833) );
  and2_1 U11877 ( .ip1(n9833), .ip2(i_ssi_risr[1]), .op(n9834) );
  nor2_1 U11878 ( .ip1(n9835), .ip2(n9834), .op(n9836) );
  nor2_1 U11879 ( .ip1(n9836), .ip2(n11148), .op(n4584) );
  mux2_1 U11880 ( .ip1(i_apb_pwdata_int[7]), .ip2(
        i_ssi_U_regfile_ctrlr0_ir_int_7), .s(n9837), .op(n4594) );
  inv_1 U11881 ( .ip(n9838), .op(n9840) );
  or3_1 U11882 ( .ip1(i_apb_pwdata_int[3]), .ip2(i_apb_pwdata_int[5]), .ip3(
        i_apb_pwdata_int[7]), .op(n9839) );
  nor4_1 U11883 ( .ip1(i_apb_pwdata_int[6]), .ip2(i_apb_pwdata_int[4]), .ip3(
        n9840), .ip4(n9839), .op(n9841) );
  mux2_1 U11884 ( .ip1(i_apb_pwdata_int[1]), .ip2(i_ssi_rxftlr[1]), .s(n9842), 
        .op(n4643) );
  mux2_1 U11885 ( .ip1(i_apb_pwdata_int[1]), .ip2(i_ssi_txftlr[1]), .s(n9843), 
        .op(n4640) );
  mux2_1 U11886 ( .ip1(i_apb_pwdata_int[2]), .ip2(i_ssi_rxftlr[2]), .s(n9842), 
        .op(n4642) );
  mux2_1 U11887 ( .ip1(i_apb_pwdata_int[2]), .ip2(i_ssi_txftlr[2]), .s(n9843), 
        .op(n4639) );
  mux2_1 U11888 ( .ip1(i_apb_pwdata_int[0]), .ip2(i_ssi_rxftlr[0]), .s(n9842), 
        .op(n4644) );
  mux2_1 U11889 ( .ip1(i_apb_pwdata_int[0]), .ip2(i_ssi_txftlr[0]), .s(n9843), 
        .op(n4641) );
  mux2_1 U11890 ( .ip1(ex_i_ahb_AHB_Slave_PID_hmastlock), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hlock), .s(ex_i_ahb_AHB_Slave_PID_hready), 
        .op(n4855) );
  mux2_1 U11891 ( .ip1(n11606), .ip2(i_ssi_prdata[24]), .s(n11697), .op(n4220)
         );
  mux2_1 U11892 ( .ip1(n11606), .ip2(i_ssi_prdata[20]), .s(n11697), .op(n4224)
         );
  mux2_1 U11893 ( .ip1(n11606), .ip2(i_ssi_prdata[21]), .s(n11697), .op(n4223)
         );
  mux2_1 U11894 ( .ip1(n11606), .ip2(i_ssi_prdata[17]), .s(n11697), .op(n4227)
         );
  nor2_1 U11895 ( .ip1(n11584), .ip2(i_ssi_ssi_txo_intr_n), .op(n9860) );
  nor2_1 U11896 ( .ip1(i_ssi_U_regfile_txflr[1]), .ip2(n9846), .op(n9845) );
  or2_1 U11897 ( .ip1(n9846), .ip2(n9845), .op(n9858) );
  inv_1 U11898 ( .ip(i_ssi_txftlr[1]), .op(n10185) );
  nor2_1 U11899 ( .ip1(n9900), .ip2(n10293), .op(n9849) );
  nor2_1 U11900 ( .ip1(n9847), .ip2(n11543), .op(n9848) );
  not_ab_or_c_or_d U11901 ( .ip1(n5395), .ip2(n11693), .ip3(n9849), .ip4(n9848), .op(n9851) );
  inv_1 U11902 ( .ip(n9852), .op(n11571) );
  mux2_1 U11903 ( .ip1(n10185), .ip2(n9853), .s(n11571), .op(n9854) );
  inv_1 U11904 ( .ip(i_ssi_rxftlr[1]), .op(n11228) );
  mux2_1 U11905 ( .ip1(n9854), .ip2(n11228), .s(n11573), .op(n9856) );
  mux2_1 U11906 ( .ip1(i_ssi_tx_full), .ip2(n9856), .s(n9855), .op(n9857) );
  nand2_1 U11907 ( .ip1(n9858), .ip2(n9857), .op(n9859) );
  not_ab_or_c_or_d U11908 ( .ip1(n11599), .ip2(i_ssi_U_regfile_rxflr[1]), 
        .ip3(n9860), .ip4(n9859), .op(n9874) );
  nand2_1 U11909 ( .ip1(i_ssi_U_dff_rx_mem[97]), .ip2(n11687), .op(n9869) );
  and2_1 U11910 ( .ip1(n11675), .ip2(i_ssi_U_dff_rx_mem[1]), .op(n9866) );
  nand2_1 U11911 ( .ip1(n11686), .ip2(i_ssi_U_dff_rx_mem[65]), .op(n9864) );
  nand2_1 U11912 ( .ip1(n11678), .ip2(i_ssi_U_dff_rx_mem[81]), .op(n9863) );
  nand2_1 U11913 ( .ip1(n11676), .ip2(i_ssi_U_dff_rx_mem[17]), .op(n9862) );
  nand2_1 U11914 ( .ip1(n11679), .ip2(i_ssi_U_dff_rx_mem[33]), .op(n9861) );
  nand4_1 U11915 ( .ip1(n9864), .ip2(n9863), .ip3(n9862), .ip4(n9861), .op(
        n9865) );
  not_ab_or_c_or_d U11916 ( .ip1(i_ssi_U_dff_rx_mem[113]), .ip2(n11674), .ip3(
        n9866), .ip4(n9865), .op(n9868) );
  nand2_1 U11917 ( .ip1(n11677), .ip2(i_ssi_U_dff_rx_mem[49]), .op(n9867) );
  nand3_1 U11918 ( .ip1(n9869), .ip2(n9868), .ip3(n9867), .op(n9870) );
  nand2_1 U11919 ( .ip1(n11598), .ip2(n9870), .op(n9873) );
  nand2_1 U11920 ( .ip1(n11600), .ip2(i_ssi_imr[1]), .op(n9872) );
  nand2_1 U11921 ( .ip1(n11587), .ip2(i_ssi_risr[1]), .op(n9871) );
  nand4_1 U11922 ( .ip1(n9874), .ip2(n9873), .ip3(n9872), .ip4(n9871), .op(
        n9875) );
  or2_1 U11923 ( .ip1(n9875), .ip2(n11606), .op(n9876) );
  mux2_1 U11924 ( .ip1(n9876), .ip2(i_ssi_prdata[1]), .s(n11697), .op(n4243)
         );
  nand2_1 U11925 ( .ip1(n11679), .ip2(i_ssi_U_dff_rx_mem[37]), .op(n9880) );
  nand2_1 U11926 ( .ip1(n11678), .ip2(i_ssi_U_dff_rx_mem[85]), .op(n9879) );
  nand2_1 U11927 ( .ip1(n11677), .ip2(i_ssi_U_dff_rx_mem[53]), .op(n9878) );
  nand2_1 U11928 ( .ip1(n11675), .ip2(i_ssi_U_dff_rx_mem[5]), .op(n9877) );
  nand4_1 U11929 ( .ip1(n9880), .ip2(n9879), .ip3(n9878), .ip4(n9877), .op(
        n9886) );
  nand2_1 U11930 ( .ip1(n11676), .ip2(i_ssi_U_dff_rx_mem[21]), .op(n9884) );
  nand2_1 U11931 ( .ip1(n11687), .ip2(i_ssi_U_dff_rx_mem[101]), .op(n9883) );
  nand2_1 U11932 ( .ip1(n11674), .ip2(i_ssi_U_dff_rx_mem[117]), .op(n9882) );
  nand2_1 U11933 ( .ip1(n11686), .ip2(i_ssi_U_dff_rx_mem[69]), .op(n9881) );
  nand4_1 U11934 ( .ip1(n9884), .ip2(n9883), .ip3(n9882), .ip4(n9881), .op(
        n9885) );
  nor2_1 U11935 ( .ip1(n9886), .ip2(n9885), .op(n9888) );
  nor2_1 U11936 ( .ip1(n9888), .ip2(n9887), .op(n9890) );
  nor2_1 U11937 ( .ip1(i_ssi_ssi_mst_intr_n), .ip2(n11584), .op(n9889) );
  not_ab_or_c_or_d U11938 ( .ip1(n11600), .ip2(i_ssi_imr[5]), .ip3(n9890), 
        .ip4(n9889), .op(n9894) );
  and2_1 U11939 ( .ip1(n11693), .ip2(i_ssi_U_regfile_ctrlr1_int[5]), .op(n9891) );
  not_ab_or_c_or_d U11940 ( .ip1(i_ssi_baudr[5]), .ip2(n11691), .ip3(n11606), 
        .ip4(n9891), .op(n9893) );
  nand2_1 U11941 ( .ip1(n11587), .ip2(i_ssi_risr[5]), .op(n9892) );
  nand3_1 U11942 ( .ip1(n9894), .ip2(n9893), .ip3(n9892), .op(n9895) );
  mux2_1 U11943 ( .ip1(n9895), .ip2(i_ssi_prdata[5]), .s(n11697), .op(n4239)
         );
  nand2_1 U11944 ( .ip1(i_apb_U_DW_apb_ahbsif_state[2]), .ip2(n11367), .op(
        n10016) );
  nand2_1 U11945 ( .ip1(n10016), .ip2(n9897), .op(n9898) );
  mux2_1 U11946 ( .ip1(i_apb_penable), .ip2(n9898), .s(i_apb_pclk_en), .op(
        n4211) );
  and2_1 U11947 ( .ip1(i_ssi_fsm_sleep), .ip2(n11148), .op(
        i_ssi_U_regfile_N451) );
  or2_1 U11948 ( .ip1(n11697), .ip2(n9902), .op(n9903) );
  nand2_1 U11949 ( .ip1(n9903), .ip2(i_ssi_risr[2]), .op(n9906) );
  nand3_1 U11950 ( .ip1(i_ssi_U_fifo_rx_pop_dly), .ip2(
        i_ssi_U_fifo_rx_error_ir), .ip3(n9904), .op(n9905) );
  nand2_1 U11951 ( .ip1(n9906), .ip2(n9905), .op(n9907) );
  and2_1 U11952 ( .ip1(n9907), .ip2(n11569), .op(n4449) );
  or2_1 U11953 ( .ip1(i_ssi_reg_addr[0]), .ip2(n11620), .op(n9911) );
  nor2_1 U11954 ( .ip1(n9909), .ip2(n9908), .op(n11605) );
  or2_1 U11955 ( .ip1(n11605), .ip2(n11620), .op(n9910) );
  nand2_1 U11956 ( .ip1(n9911), .ip2(n9910), .op(n11614) );
  nor2_1 U11957 ( .ip1(n11697), .ip2(n11614), .op(n9915) );
  inv_1 U11958 ( .ip(n9915), .op(n9912) );
  nand2_1 U11959 ( .ip1(n9912), .ip2(i_ssi_risr[5]), .op(n9913) );
  and2_1 U11960 ( .ip1(n9914), .ip2(n11569), .op(n4247) );
  nand2_1 U11961 ( .ip1(i_ssi_mst_contention), .ip2(i_ssi_risr[5]), .op(n9916)
         );
  nor2_1 U11962 ( .ip1(n9916), .ip2(n9915), .op(n9919) );
  inv_1 U11963 ( .ip(n9917), .op(n9918) );
  inv_1 U11964 ( .ip(i_ssi_risr[5]), .op(n9921) );
  and2_1 U11965 ( .ip1(n9925), .ip2(n11569), .op(n4246) );
  fulladder U11966 ( .a(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[6]), .b(n9927), .ci(n9926), .co(n9929), .s(n6962) );
  xor2_1 U11967 ( .ip1(n9927), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[7]), .op(n9928) );
  xor2_1 U11968 ( .ip1(n9929), .ip2(n9928), .op(n9931) );
  nand2_1 U11969 ( .ip1(n9931), .ip2(n9930), .op(n9934) );
  nand2_1 U11970 ( .ip1(n9932), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[7]), .op(n9933) );
  nand2_1 U11971 ( .ip1(n9934), .ip2(n9933), .op(n4135) );
  inv_1 U11972 ( .ip(n9935), .op(n9936) );
  nor2_1 U11973 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_hcnt_cmplt_int), .ip2(
        n9936), .op(n9937) );
  nor2_1 U11974 ( .ip1(n10275), .ip2(n9937), .op(n4166) );
  inv_1 U11975 ( .ip(n10958), .op(n10960) );
  nor2_1 U11976 ( .ip1(n10960), .ip2(i_i2c_scl_s_setup_cmplt), .op(n9938) );
  nor2_1 U11977 ( .ip1(n9938), .ip2(n10994), .op(n5197) );
  inv_1 U11978 ( .ip(n10634), .op(n10636) );
  nor2_1 U11979 ( .ip1(n10636), .ip2(i_i2c_scl_p_setup_cmplt), .op(n9939) );
  nor2_1 U11980 ( .ip1(n9939), .ip2(n10677), .op(n5051) );
  inv_1 U11981 ( .ip(n10918), .op(n10920) );
  nor2_1 U11982 ( .ip1(n10920), .ip2(i_i2c_U_DW_apb_i2c_mstfsm_N382), .op(
        n9940) );
  nor2_1 U11983 ( .ip1(n9940), .ip2(n10955), .op(n5119) );
  inv_1 U11984 ( .ip(n10997), .op(n10999) );
  nor2_1 U11985 ( .ip1(n10999), .ip2(i_i2c_scl_s_hld_cmplt), .op(n9941) );
  nor2_1 U11986 ( .ip1(n11041), .ip2(n9941), .op(n5195) );
  nand2_1 U11987 ( .ip1(n9942), .ip2(n6404), .op(n9943) );
  nand2_1 U11988 ( .ip1(n9944), .ip2(n9943), .op(n9945) );
  nor2_1 U11989 ( .ip1(n10275), .ip2(n9945), .op(n4163) );
  nand2_1 U11990 ( .ip1(n9973), .ip2(n9969), .op(n9948) );
  inv_1 U11991 ( .ip(n9946), .op(n9947) );
  nand2_1 U11992 ( .ip1(n10965), .ip2(n9950), .op(n9951) );
  nand2_1 U11993 ( .ip1(i_i2c_scl_s_setup_en), .ip2(n9951), .op(n9952) );
  nor2_1 U11994 ( .ip1(n10969), .ip2(n9952), .op(n5150) );
  and2_1 U11995 ( .ip1(n11767), .ip2(n9954), .op(i_ssi_U_fifo_U_tx_fifo_N39)
         );
  nand2_1 U11996 ( .ip1(n10061), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_start_sda_gate_r), .op(n11103) );
  and3_1 U11997 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda_r), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_start_sda), .op(n11104) );
  or3_1 U11998 ( .ip1(i_i2c_ic_clk_oe), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_start_sda_gate_r), .ip3(n11104), .op(n9955) );
  nand2_1 U11999 ( .ip1(n11103), .ip2(n9955), .op(
        i_i2c_U_DW_apb_i2c_tx_shift_N272) );
  nand2_1 U12000 ( .ip1(n9956), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[3]), .op(n9957) );
  nand2_1 U12001 ( .ip1(n9957), .ip2(n6409), .op(n9958) );
  nand2_1 U12002 ( .ip1(n9980), .ip2(n9958), .op(n9959) );
  nor2_1 U12003 ( .ip1(n10275), .ip2(n9959), .op(n4161) );
  inv_1 U12004 ( .ip(i_ssi_U_mstfsm_ctrl_cnt[1]), .op(n11704) );
  inv_1 U12005 ( .ip(i_ssi_U_mstfsm_ctrl_cnt[2]), .op(n11706) );
  xor2_1 U12006 ( .ip1(i_ssi_cfs[3]), .ip2(i_ssi_U_mstfsm_ctrl_cnt[3]), .op(
        n9962) );
  xor2_1 U12007 ( .ip1(i_ssi_cfs[0]), .ip2(i_ssi_U_mstfsm_ctrl_cnt[0]), .op(
        n9961) );
  nor2_1 U12008 ( .ip1(n9968), .ip2(n9967), .op(n4587) );
  inv_1 U12009 ( .ip(i_ssi_U_regfile_txflr[1]), .op(n10545) );
  inv_1 U12010 ( .ip(n11519), .op(n9978) );
  inv_1 U12011 ( .ip(i_ssi_U_regfile_txflr[2]), .op(n11514) );
  inv_1 U12012 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[5]), .op(n9979)
         );
  nand2_1 U12013 ( .ip1(n9980), .ip2(n9979), .op(n9981) );
  nand2_1 U12014 ( .ip1(n9982), .ip2(n9981), .op(n9983) );
  nor2_1 U12015 ( .ip1(n10275), .ip2(n9983), .op(n4160) );
  mux2_1 U12016 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[0]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[1]), .s(n10051), .op(n4393) );
  mux2_1 U12017 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[1]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[2]), .s(n10051), .op(n4392) );
  mux2_1 U12018 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[6]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[7]), .s(n10051), .op(n4387) );
  mux2_1 U12019 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[2]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[3]), .s(n10051), .op(n4391) );
  mux2_1 U12020 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[4]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[5]), .s(n10051), .op(n4389) );
  mux2_1 U12021 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[3]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[4]), .s(n10051), .op(n4390) );
  nand2_1 U12022 ( .ip1(i_ssi_U_mstfsm_ss_in_n_sync), .ip2(n9986), .op(n9987)
         );
  nand2_1 U12023 ( .ip1(n11569), .ip2(n9987), .op(i_ssi_U_mstfsm_N221) );
  inv_1 U12024 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[7]), .op(n9990)
         );
  nand2_1 U12025 ( .ip1(n9988), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[6]), .op(n9989) );
  nand2_1 U12026 ( .ip1(n9990), .ip2(n9989), .op(n9991) );
  nand2_1 U12027 ( .ip1(n10058), .ip2(n9991), .op(n9992) );
  nor2_1 U12028 ( .ip1(n10275), .ip2(n9992), .op(n4158) );
  nor3_1 U12029 ( .ip1(i_i2c_scl_s_setup_en), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_scl_hld_low_en_r), .ip3(n9993), .op(n9995)
         );
  inv_1 U12030 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_re_scl_s_hld_en), .op(n9994)
         );
  nand4_1 U12031 ( .ip1(n9995), .ip2(n11771), .ip3(n10677), .ip4(n9994), .op(
        n9996) );
  nor4_1 U12032 ( .ip1(n5109), .ip2(i_i2c_rx_scl_lcnt_en), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_data_scl_lcnt_en), .ip4(n9996), .op(n9998)
         );
  nand4_1 U12033 ( .ip1(i_i2c_mst_rx_data_scl), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_stop_scl), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl), .ip4(
        i_i2c_U_DW_apb_i2c_tx_shift_data_scl), .op(n10000) );
  nor3_1 U12034 ( .ip1(n11105), .ip2(i_i2c_scl_hld_low_en), .ip3(n10000), .op(
        n10001) );
  not_ab_or_c_or_d U12035 ( .ip1(n11105), .ip2(n10005), .ip3(n10001), .ip4(
        n11110), .op(n10007) );
  not_ab_or_c_or_d U12036 ( .ip1(n10061), .ip2(n10003), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_mst_slv_ack_ext_r), .ip4(n10002), .op(
        n11106) );
  nor3_1 U12037 ( .ip1(n11106), .ip2(n10005), .ip3(n10004), .op(n10006) );
  or2_1 U12038 ( .ip1(n10007), .ip2(n10006), .op(n4958) );
  inv_1 U12039 ( .ip(n10008), .op(n10010) );
  or2_1 U12040 ( .ip1(n10009), .ip2(n10010), .op(n10013) );
  nand2_1 U12041 ( .ip1(n10013), .ip2(n10012), .op(n10014) );
  or2_1 U12042 ( .ip1(n10014), .ip2(i_apb_U_DW_apb_ahbsif_nextstate[2]), .op(
        n10015) );
  nand2_1 U12043 ( .ip1(n10016), .ip2(n10015), .op(n10030) );
  nor3_2 U12044 ( .ip1(n10017), .ip2(i_apb_U_DW_apb_ahbsif_nextstate[2]), 
        .ip3(n5311), .op(n11361) );
  not_ab_or_c_or_d U12045 ( .ip1(n10026), .ip2(n10110), .ip3(n10018), .ip4(
        n11361), .op(n10023) );
  nor3_1 U12046 ( .ip1(n10021), .ip2(n10020), .ip3(n10019), .op(n10022) );
  not_ab_or_c_or_d U12047 ( .ip1(n10025), .ip2(n10024), .ip3(n10023), .ip4(
        n10022), .op(n10028) );
  nand3_1 U12048 ( .ip1(i_apb_U_DW_apb_ahbsif_nextstate[1]), .ip2(n10026), 
        .ip3(i_apb_U_DW_apb_ahbsif_pipeline_c), .op(n10027) );
  nand2_1 U12049 ( .ip1(n10028), .ip2(n10027), .op(n10029) );
  nor3_2 U12050 ( .ip1(i_ssi_tx_wr_addr[1]), .ip2(n10165), .ip3(n11211), .op(
        n10033) );
  nand2_1 U12051 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[15]), .ip2(n11461), 
        .op(n10044) );
  nand2_1 U12052 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[15]), .ip2(n5270), 
        .op(n10043) );
  nand2_1 U12053 ( .ip1(n10044), .ip2(n10043), .op(n4750) );
  nand2_1 U12054 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[13]), .ip2(n11461), 
        .op(n10046) );
  nand2_1 U12055 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[13]), .ip2(n5270), 
        .op(n10045) );
  nand2_1 U12056 ( .ip1(n10046), .ip2(n10045), .op(n4752) );
  inv_1 U12057 ( .ip(n11221), .op(n10048) );
  mux2_1 U12058 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[14]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[15]), .s(n10051), .op(n4379)
         );
  mux2_1 U12059 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[10]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[11]), .s(n10051), .op(n4383)
         );
  mux2_1 U12060 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[9]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[10]), .s(n10051), .op(n4384)
         );
  mux2_1 U12061 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[12]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[13]), .s(n10051), .op(n4381)
         );
  mux2_1 U12062 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[8]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[9]), .s(n10051), .op(n4385) );
  mux2_1 U12063 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[11]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[12]), .s(n10051), .op(n4382)
         );
  mux2_1 U12064 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[7]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[8]), .s(n10051), .op(n4386) );
  mux2_1 U12065 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[13]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[14]), .s(n10051), .op(n4380)
         );
  mux2_1 U12066 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[5]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[6]), .s(n10051), .op(n4388) );
  inv_1 U12067 ( .ip(n10052), .op(n10053) );
  nand2_1 U12068 ( .ip1(n10053), .ip2(i_ssi_U_fifo_unconnected_tx_wrd_count[0]), .op(n10054) );
  nand2_1 U12069 ( .ip1(n10055), .ip2(n10054), .op(n10188) );
  and2_1 U12070 ( .ip1(n10188), .ip2(n11219), .op(i_ssi_U_fifo_U_tx_fifo_N47)
         );
  nor3_1 U12071 ( .ip1(i_ssi_U_fifo_U_tx_fifo_N37), .ip2(
        i_ssi_U_fifo_U_tx_fifo_N47), .ip3(n11779), .op(n10057) );
  inv_1 U12072 ( .ip(i_ssi_U_fifo_U_tx_fifo_N48), .op(n10056) );
  nand2_1 U12073 ( .ip1(n10057), .ip2(n10056), .op(i_ssi_U_fifo_U_tx_fifo_N33)
         );
  nand2_1 U12074 ( .ip1(n10058), .ip2(n6429), .op(n10059) );
  nand2_1 U12075 ( .ip1(n10216), .ip2(n10059), .op(n10060) );
  nor2_1 U12076 ( .ip1(n10275), .ip2(n10060), .op(n4157) );
  inv_1 U12077 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_stop_sda), .op(n10063) );
  nand2_1 U12078 ( .ip1(n10061), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_stop_sda_gate_r), .op(n10062) );
  nand2_1 U12079 ( .ip1(n10063), .ip2(n10062), .op(
        i_i2c_U_DW_apb_i2c_tx_shift_N281) );
  inv_1 U12080 ( .ip(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[3]), .op(n10068)
         );
  nor2_1 U12081 ( .ip1(n11543), .ip2(n10198), .op(n11558) );
  inv_1 U12082 ( .ip(n10205), .op(n10066) );
  mux2_1 U12083 ( .ip1(i_ssi_rx_push_data[3]), .ip2(n10069), .s(n5266), .op(
        n4442) );
  inv_1 U12084 ( .ip(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[4]), .op(n10070)
         );
  nor2_1 U12085 ( .ip1(n10070), .ip2(n10205), .op(n10071) );
  mux2_1 U12086 ( .ip1(i_ssi_rx_push_data[4]), .ip2(n10071), .s(n5266), .op(
        n4441) );
  mux2_1 U12087 ( .ip1(i_ssi_rx_push_data[0]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[0]), .s(n5266), .op(n4378) );
  nand2_1 U12088 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[29]), .ip2(n11465), 
        .op(n10073) );
  nand2_1 U12089 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[29]), .ip2(n5270), 
        .op(n10072) );
  nand2_1 U12090 ( .ip1(n10073), .ip2(n10072), .op(n4736) );
  nand2_1 U12091 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[16]), .ip2(n11461), 
        .op(n10075) );
  nand2_1 U12092 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[16]), .ip2(n5270), 
        .op(n10074) );
  nand2_1 U12093 ( .ip1(n10075), .ip2(n10074), .op(n4749) );
  nand2_1 U12094 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[22]), .ip2(n11461), 
        .op(n10077) );
  nand2_1 U12095 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[22]), .ip2(n5270), 
        .op(n10076) );
  nand2_1 U12096 ( .ip1(n10077), .ip2(n10076), .op(n4743) );
  nand2_1 U12097 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[21]), .ip2(n11465), 
        .op(n10079) );
  nand2_1 U12098 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[21]), .ip2(n5270), 
        .op(n10078) );
  nand2_1 U12099 ( .ip1(n10079), .ip2(n10078), .op(n4744) );
  nand2_1 U12100 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[28]), .ip2(n11461), 
        .op(n10081) );
  nand2_1 U12101 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[28]), .ip2(n5270), 
        .op(n10080) );
  nand2_1 U12102 ( .ip1(n10081), .ip2(n10080), .op(n4737) );
  nand2_1 U12103 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[19]), .ip2(n11461), 
        .op(n10083) );
  nand2_1 U12104 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[19]), .ip2(n5270), 
        .op(n10082) );
  nand2_1 U12105 ( .ip1(n10083), .ip2(n10082), .op(n4746) );
  nand2_1 U12106 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[20]), .ip2(n11461), 
        .op(n10085) );
  nand2_1 U12107 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[20]), .ip2(n5270), 
        .op(n10084) );
  nand2_1 U12108 ( .ip1(n10085), .ip2(n10084), .op(n4745) );
  nand2_1 U12109 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[18]), .ip2(n11461), 
        .op(n10087) );
  nand2_1 U12110 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[18]), .ip2(n5270), 
        .op(n10086) );
  nand2_1 U12111 ( .ip1(n10087), .ip2(n10086), .op(n4747) );
  nand2_1 U12112 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[30]), .ip2(n11461), 
        .op(n10089) );
  nand2_1 U12113 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[30]), .ip2(n5270), 
        .op(n10088) );
  nand2_1 U12114 ( .ip1(n10089), .ip2(n10088), .op(n4735) );
  nand2_1 U12115 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[26]), .ip2(n11461), 
        .op(n10091) );
  nand2_1 U12116 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[26]), .ip2(n5270), 
        .op(n10090) );
  nand2_1 U12117 ( .ip1(n10091), .ip2(n10090), .op(n4739) );
  nand2_1 U12118 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[24]), .ip2(n11461), 
        .op(n10093) );
  nand2_1 U12119 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[24]), .ip2(n5270), 
        .op(n10092) );
  nand2_1 U12120 ( .ip1(n10093), .ip2(n10092), .op(n4741) );
  nand2_1 U12121 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[25]), .ip2(n11461), 
        .op(n10095) );
  nand2_1 U12122 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[25]), .ip2(n5270), 
        .op(n10094) );
  nand2_1 U12123 ( .ip1(n10095), .ip2(n10094), .op(n4740) );
  nand2_1 U12124 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[23]), .ip2(n11465), 
        .op(n10097) );
  nand2_1 U12125 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[23]), .ip2(n5270), 
        .op(n10096) );
  nand2_1 U12126 ( .ip1(n10097), .ip2(n10096), .op(n4742) );
  nand2_1 U12127 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[27]), .ip2(n11461), 
        .op(n10099) );
  nand2_1 U12128 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[27]), .ip2(n5270), 
        .op(n10098) );
  nand2_1 U12129 ( .ip1(n10099), .ip2(n10098), .op(n4738) );
  nand2_1 U12130 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[14]), .ip2(n11465), 
        .op(n10101) );
  nand2_1 U12131 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[14]), .ip2(n5270), 
        .op(n10100) );
  nand2_1 U12132 ( .ip1(n10101), .ip2(n10100), .op(n4751) );
  nand2_1 U12133 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[31]), .ip2(n11461), 
        .op(n10103) );
  nand2_1 U12134 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[31]), .ip2(n5270), 
        .op(n10102) );
  nand2_1 U12135 ( .ip1(n10103), .ip2(n10102), .op(n4734) );
  nand2_1 U12136 ( .ip1(i_apb_pclk_en), .ip2(n11361), .op(n10104) );
  nor2_1 U12137 ( .ip1(n10106), .ip2(n10105), .op(n10109) );
  nand2_1 U12138 ( .ip1(i_apb_paddr[21]), .ip2(n11497), .op(n10115) );
  nor2_1 U12139 ( .ip1(n10108), .ip2(n10107), .op(n11470) );
  nand2_1 U12140 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[21]), .ip2(n11507), 
        .op(n10114) );
  nand3_1 U12141 ( .ip1(n10110), .ip2(n10109), .ip3(n11471), .op(n10112) );
  nand2_1 U12142 ( .ip1(i_apb_U_DW_apb_ahbsif_use_saved_c), .ip2(n11369), .op(
        n10111) );
  nand2_1 U12143 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[21]), .ip2(n5269), 
        .op(n10113) );
  nand3_1 U12144 ( .ip1(n10115), .ip2(n10114), .ip3(n10113), .op(n4718) );
  nand2_1 U12145 ( .ip1(i_apb_paddr[13]), .ip2(n11497), .op(n10119) );
  nand2_1 U12146 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[13]), .ip2(n11507), 
        .op(n10118) );
  nand2_1 U12147 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[13]), .ip2(n5269), 
        .op(n10117) );
  nand3_1 U12148 ( .ip1(n10119), .ip2(n10118), .ip3(n10117), .op(n4726) );
  nand2_1 U12149 ( .ip1(i_apb_paddr[18]), .ip2(n11497), .op(n10122) );
  nand2_1 U12150 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[18]), .ip2(n11507), 
        .op(n10121) );
  nand2_1 U12151 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[18]), .ip2(n5269), 
        .op(n10120) );
  nand3_1 U12152 ( .ip1(n10122), .ip2(n10121), .ip3(n10120), .op(n4721) );
  nand2_1 U12153 ( .ip1(i_apb_paddr[15]), .ip2(n11497), .op(n10125) );
  nand2_1 U12154 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[15]), .ip2(n11507), 
        .op(n10124) );
  nand2_1 U12155 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[15]), .ip2(n5269), 
        .op(n10123) );
  nand3_1 U12156 ( .ip1(n10125), .ip2(n10124), .ip3(n10123), .op(n4724) );
  nand2_1 U12157 ( .ip1(i_apb_paddr[14]), .ip2(n11497), .op(n10128) );
  nand2_1 U12158 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[14]), .ip2(n11507), 
        .op(n10127) );
  nand2_1 U12159 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[14]), .ip2(n5269), 
        .op(n10126) );
  nand3_1 U12160 ( .ip1(n10128), .ip2(n10127), .ip3(n10126), .op(n4725) );
  nand2_1 U12161 ( .ip1(i_apb_paddr[23]), .ip2(n11497), .op(n10131) );
  nand2_1 U12162 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[23]), .ip2(n11507), 
        .op(n10130) );
  nand2_1 U12163 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[23]), .ip2(n5269), 
        .op(n10129) );
  nand3_1 U12164 ( .ip1(n10131), .ip2(n10130), .ip3(n10129), .op(n4716) );
  nand2_1 U12165 ( .ip1(i_apb_paddr[25]), .ip2(n11497), .op(n10134) );
  nand2_1 U12166 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[25]), .ip2(n11507), 
        .op(n10133) );
  nand2_1 U12167 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[25]), .ip2(n5269), 
        .op(n10132) );
  nand3_1 U12168 ( .ip1(n10134), .ip2(n10133), .ip3(n10132), .op(n4714) );
  nand2_1 U12169 ( .ip1(i_apb_paddr[29]), .ip2(n11497), .op(n10137) );
  nand2_1 U12170 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[29]), .ip2(n11507), 
        .op(n10136) );
  nand2_1 U12171 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[29]), .ip2(n5269), 
        .op(n10135) );
  nand3_1 U12172 ( .ip1(n10137), .ip2(n10136), .ip3(n10135), .op(n4710) );
  nand2_1 U12173 ( .ip1(i_apb_paddr[26]), .ip2(n11497), .op(n10140) );
  nand2_1 U12174 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[26]), .ip2(n11507), 
        .op(n10139) );
  nand2_1 U12175 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[26]), .ip2(n5269), 
        .op(n10138) );
  nand3_1 U12176 ( .ip1(n10140), .ip2(n10139), .ip3(n10138), .op(n4713) );
  nand2_1 U12177 ( .ip1(i_apb_paddr[22]), .ip2(n11497), .op(n10143) );
  nand2_1 U12178 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[22]), .ip2(n11507), 
        .op(n10142) );
  nand2_1 U12179 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[22]), .ip2(n5269), 
        .op(n10141) );
  nand3_1 U12180 ( .ip1(n10143), .ip2(n10142), .ip3(n10141), .op(n4717) );
  nand2_1 U12181 ( .ip1(i_apb_paddr[31]), .ip2(n11497), .op(n10146) );
  nand2_1 U12182 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[31]), .ip2(n11507), 
        .op(n10145) );
  nand2_1 U12183 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[31]), .ip2(n5269), 
        .op(n10144) );
  nand3_1 U12184 ( .ip1(n10146), .ip2(n10145), .ip3(n10144), .op(n4708) );
  nand2_1 U12185 ( .ip1(i_apb_paddr[16]), .ip2(n11497), .op(n10149) );
  nand2_1 U12186 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[16]), .ip2(n11507), 
        .op(n10148) );
  nand2_1 U12187 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[16]), .ip2(n5269), 
        .op(n10147) );
  nand3_1 U12188 ( .ip1(n10149), .ip2(n10148), .ip3(n10147), .op(n4723) );
  nand2_1 U12189 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[30]), .ip2(n11507), 
        .op(n10152) );
  nand2_1 U12190 ( .ip1(i_apb_paddr[30]), .ip2(n11497), .op(n10151) );
  nand2_1 U12191 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[30]), .ip2(n5269), 
        .op(n10150) );
  nand3_1 U12192 ( .ip1(n10152), .ip2(n10151), .ip3(n10150), .op(n4709) );
  nand2_1 U12193 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[27]), .ip2(n11507), 
        .op(n10155) );
  nand2_1 U12194 ( .ip1(i_apb_paddr[27]), .ip2(n11497), .op(n10154) );
  nand2_1 U12195 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[27]), .ip2(n5269), 
        .op(n10153) );
  nand3_1 U12196 ( .ip1(n10155), .ip2(n10154), .ip3(n10153), .op(n4712) );
  nand2_1 U12197 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[24]), .ip2(n11507), 
        .op(n10158) );
  nand2_1 U12198 ( .ip1(i_apb_paddr[24]), .ip2(n11497), .op(n10157) );
  nand2_1 U12199 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[24]), .ip2(n5269), 
        .op(n10156) );
  nand3_1 U12200 ( .ip1(n10158), .ip2(n10157), .ip3(n10156), .op(n4715) );
  nand2_1 U12201 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[20]), .ip2(n11507), 
        .op(n10161) );
  nand2_1 U12202 ( .ip1(i_apb_paddr[20]), .ip2(n11497), .op(n10160) );
  nand2_1 U12203 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[20]), .ip2(n5269), 
        .op(n10159) );
  nand3_1 U12204 ( .ip1(n10161), .ip2(n10160), .ip3(n10159), .op(n4719) );
  nand2_1 U12205 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[19]), .ip2(n11507), 
        .op(n10164) );
  nand2_1 U12206 ( .ip1(i_apb_paddr[19]), .ip2(n11497), .op(n10163) );
  nand2_1 U12207 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[19]), .ip2(n5269), 
        .op(n10162) );
  nand3_1 U12208 ( .ip1(n10164), .ip2(n10163), .ip3(n10162), .op(n4720) );
  nor2_1 U12209 ( .ip1(i_ssi_txftlr[1]), .ip2(n11227), .op(n10179) );
  nor2_1 U12210 ( .ip1(n10179), .ip2(i_ssi_U_fifo_U_tx_fifo_N48), .op(n10180)
         );
  or2_1 U12211 ( .ip1(i_ssi_txftlr[2]), .ip2(n10180), .op(n10183) );
  nand2_4 U12212 ( .ip1(n10184), .ip2(i_ssi_txftlr[1]), .op(n10181) );
  nand2_1 U12213 ( .ip1(n11779), .ip2(n10181), .op(n10182) );
  nand2_1 U12214 ( .ip1(n10183), .ip2(n10182), .op(n10192) );
  inv_4 U12215 ( .ip(n10184), .op(n10186) );
  nand2_1 U12216 ( .ip1(n10186), .ip2(n10185), .op(n10190) );
  inv_1 U12217 ( .ip(i_ssi_txftlr[0]), .op(n10187) );
  nand2_1 U12218 ( .ip1(n10190), .ip2(n10189), .op(n10191) );
  nand2_1 U12219 ( .ip1(n10192), .ip2(n10191), .op(n10196) );
  inv_1 U12220 ( .ip(i_ssi_txftlr[2]), .op(n10193) );
  and2_1 U12221 ( .ip1(n11779), .ip2(n10193), .op(n10194) );
  nand2_1 U12222 ( .ip1(n10196), .ip2(n10195), .op(i_ssi_U_fifo_U_tx_fifo_N34)
         );
  inv_1 U12223 ( .ip(i_ssi_rx_push_data[5]), .op(n10197) );
  nor2_1 U12224 ( .ip1(n10197), .ip2(n5266), .op(n10202) );
  nand2_1 U12225 ( .ip1(n5266), .ip2(n11555), .op(n10200) );
  nand2_1 U12226 ( .ip1(n5266), .ip2(n5358), .op(n11536) );
  inv_1 U12227 ( .ip(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[5]), .op(n10199)
         );
  not_ab_or_c_or_d U12228 ( .ip1(n10200), .ip2(n11536), .ip3(n10205), .ip4(
        n10199), .op(n10201) );
  or2_1 U12229 ( .ip1(n10202), .ip2(n10201), .op(n4440) );
  inv_1 U12230 ( .ip(i_ssi_rx_push_data[7]), .op(n10203) );
  nor2_1 U12231 ( .ip1(n10203), .ip2(n5266), .op(n10208) );
  nand2_1 U12232 ( .ip1(n5266), .ip2(n11558), .op(n10206) );
  inv_1 U12233 ( .ip(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[7]), .op(n10204)
         );
  not_ab_or_c_or_d U12234 ( .ip1(n10206), .ip2(n11536), .ip3(n10205), .ip4(
        n10204), .op(n10207) );
  or2_1 U12235 ( .ip1(n10208), .ip2(n10207), .op(n4438) );
  nor2_1 U12236 ( .ip1(n11547), .ip2(n11536), .op(n11559) );
  nand3_1 U12237 ( .ip1(n11559), .ip2(n5398), .ip3(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[14]), .op(n10210) );
  nand2_1 U12238 ( .ip1(n6655), .ip2(i_ssi_rx_push_data[14]), .op(n10209) );
  nand2_1 U12239 ( .ip1(n10210), .ip2(n10209), .op(n4431) );
  nand3_1 U12240 ( .ip1(n5266), .ip2(n5398), .ip3(n5356), .op(n10211) );
  nand2_1 U12241 ( .ip1(n10211), .ip2(n11536), .op(n10212) );
  nand2_1 U12242 ( .ip1(n10212), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[6]), .op(n10214) );
  nand2_1 U12243 ( .ip1(n6655), .ip2(i_ssi_rx_push_data[6]), .op(n10213) );
  nand2_1 U12244 ( .ip1(n10214), .ip2(n10213), .op(n4439) );
  inv_1 U12245 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[9]), .op(n10215)
         );
  nand2_1 U12246 ( .ip1(n10216), .ip2(n10215), .op(n10217) );
  nand2_1 U12247 ( .ip1(n10228), .ip2(n10217), .op(n10218) );
  nor2_1 U12248 ( .ip1(n10275), .ip2(n10218), .op(n4156) );
  or2_1 U12249 ( .ip1(n10219), .ip2(n10220), .op(n10222) );
  or2_1 U12250 ( .ip1(i_ssi_U_fifo_unconnected_rx_wrd_count[0]), .ip2(n10220), 
        .op(n10221) );
  nor2_1 U12251 ( .ip1(n11235), .ip2(n11227), .op(i_ssi_U_fifo_U_rx_fifo_N47)
         );
  nor2_1 U12252 ( .ip1(i_ssi_U_fifo_unconnected_rx_wrd_count[0]), .ip2(n10223), 
        .op(n10224) );
  nor2_1 U12253 ( .ip1(n10225), .ip2(n10224), .op(n10226) );
  xor2_1 U12254 ( .ip1(i_ssi_U_fifo_unconnected_rx_wrd_count[1]), .ip2(n10226), 
        .op(n11232) );
  inv_1 U12255 ( .ip(n11232), .op(n10227) );
  nor2_1 U12256 ( .ip1(n10227), .ip2(n11227), .op(i_ssi_U_fifo_U_rx_fifo_N48)
         );
  nand2_1 U12257 ( .ip1(n10228), .ip2(n6385), .op(n10229) );
  nand2_1 U12258 ( .ip1(n10237), .ip2(n10229), .op(n10230) );
  nor2_1 U12259 ( .ip1(n10275), .ip2(n10230), .op(n4155) );
  nand2_1 U12260 ( .ip1(n10232), .ip2(n10231), .op(n10235) );
  inv_1 U12261 ( .ip(n10542), .op(n10233) );
  nand2_1 U12262 ( .ip1(n10233), .ip2(i_ssi_U_mstfsm_abort_ir), .op(n10234) );
  nand2_1 U12263 ( .ip1(n10235), .ip2(n10234), .op(n4428) );
  inv_1 U12264 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[11]), .op(n10236) );
  nand2_1 U12265 ( .ip1(n10237), .ip2(n10236), .op(n10238) );
  nand2_1 U12266 ( .ip1(n10242), .ip2(n10238), .op(n10239) );
  nor2_1 U12267 ( .ip1(n10275), .ip2(n10239), .op(n4154) );
  nor3_1 U12268 ( .ip1(n10240), .ip2(n11148), .ip3(n5362), .op(
        i_ssi_U_mstfsm_N222) );
  nand2_1 U12269 ( .ip1(n10241), .ip2(n5400), .op(n4183) );
  nand2_1 U12270 ( .ip1(n10242), .ip2(n6446), .op(n10243) );
  nand2_1 U12271 ( .ip1(n10244), .ip2(n10243), .op(n10245) );
  nor2_1 U12272 ( .ip1(n10275), .ip2(n10245), .op(n4153) );
  nand2_1 U12273 ( .ip1(n10263), .ip2(i_ssi_U_mstfsm_ss_in_n_sync), .op(n10264) );
  nand2_1 U12274 ( .ip1(n11569), .ip2(n10264), .op(i_ssi_U_mstfsm_N220) );
  nand2_1 U12275 ( .ip1(n10265), .ip2(i_ssi_U_mstfsm_ss_in_n_sync), .op(n10266) );
  nand2_1 U12276 ( .ip1(n10266), .ip2(n11569), .op(i_ssi_U_mstfsm_N223) );
  inv_1 U12277 ( .ip(n10267), .op(n10995) );
  nor2_1 U12278 ( .ip1(n10995), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[14]), .op(n10269) );
  nor3_1 U12279 ( .ip1(n10269), .ip2(n10994), .ip3(n10268), .op(n5139) );
  inv_1 U12280 ( .ip(n10270), .op(n10271) );
  nand2_1 U12281 ( .ip1(n10271), .ip2(n6442), .op(n10272) );
  nand2_1 U12282 ( .ip1(n10273), .ip2(n10272), .op(n10274) );
  nor2_1 U12283 ( .ip1(n10275), .ip2(n10274), .op(n4151) );
  inv_1 U12284 ( .ip(i_ssi_U_shift_U_tx_shifter_tx_buffer[1]), .op(n10279) );
  nor2_1 U12285 ( .ip1(n10279), .ip2(n10278), .op(n10283) );
  nor4_1 U12286 ( .ip1(n10284), .ip2(n10283), .ip3(n10282), .ip4(n10281), .op(
        n10286) );
  nor2_1 U12287 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[1]), .ip2(n6144), .op(n10285) );
  nor2_1 U12288 ( .ip1(n10286), .ip2(n10285), .op(n4409) );
  inv_1 U12289 ( .ip(i_ssi_sclk_active), .op(n10332) );
  nor2_1 U12290 ( .ip1(n10287), .ip2(n10303), .op(n10290) );
  or2_1 U12291 ( .ip1(n10290), .ip2(n10289), .op(n10291) );
  nor2_1 U12292 ( .ip1(n5362), .ip2(n10291), .op(n10292) );
  nor2_1 U12293 ( .ip1(n10304), .ip2(n10292), .op(n10309) );
  nand2_1 U12294 ( .ip1(n10294), .ip2(n10293), .op(n10300) );
  nor4_1 U12295 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[5]), .ip2(
        i_ssi_U_sclkgen_ssi_cnt[6]), .ip3(i_ssi_U_sclkgen_ssi_cnt[7]), .ip4(
        i_ssi_U_sclkgen_ssi_cnt[8]), .op(n10298) );
  nand4_1 U12296 ( .ip1(n10298), .ip2(n10297), .ip3(n10296), .ip4(n10295), 
        .op(n10299) );
  nor2_1 U12297 ( .ip1(n10335), .ip2(i_ssi_sclk_active), .op(n10308) );
  nand2_1 U12298 ( .ip1(n10304), .ip2(n10303), .op(n10305) );
  nor3_1 U12299 ( .ip1(n5362), .ip2(i_ssi_sclk_active), .ip3(n10305), .op(
        n10307) );
  not_ab_or_c_or_d U12300 ( .ip1(n10332), .ip2(n10309), .ip3(n10307), .ip4(
        n10308), .op(n10339) );
  inv_1 U12301 ( .ip(n10309), .op(n10337) );
  inv_1 U12302 ( .ip(i_ssi_sclk_out), .op(n10331) );
  xnor2_1 U12303 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[8]), .ip2(n11652), .op(n10314)
         );
  and4_1 U12304 ( .ip1(n10314), .ip2(n10313), .ip3(n10312), .ip4(n10311), .op(
        n10329) );
  xor2_1 U12305 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[1]), .ip2(n10384), .op(n10318)
         );
  xor2_1 U12306 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[13]), .ip2(i_ssi_baudr[14]), 
        .op(n10317) );
  xor2_1 U12307 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[11]), .ip2(i_ssi_baudr[12]), 
        .op(n10316) );
  xor2_1 U12308 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[9]), .ip2(n5257), .op(n10315)
         );
  xor2_1 U12309 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[7]), .ip2(i_ssi_baudr[8]), .op(
        n10319) );
  xor2_1 U12310 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[10]), .ip2(n6224), .op(n10325)
         );
  xor2_1 U12311 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[12]), .ip2(i_ssi_baudr[13]), 
        .op(n10324) );
  nand4_1 U12312 ( .ip1(n10329), .ip2(n10328), .ip3(n10327), .ip4(n10326), 
        .op(n10330) );
  mux2_1 U12313 ( .ip1(n10332), .ip2(n10331), .s(n10330), .op(n10333) );
  inv_1 U12314 ( .ip(n10333), .op(n10336) );
  nand2_1 U12315 ( .ip1(n10339), .ip2(n10338), .op(n4249) );
  not_ab_or_c_or_d U12316 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_buffer[15]), 
        .ip2(n10346), .ip3(n10345), .ip4(n10344), .op(n10347) );
  nand2_1 U12317 ( .ip1(n10348), .ip2(n10347), .op(n10354) );
  inv_1 U12318 ( .ip(n10350), .op(n10351) );
  nor2_1 U12319 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[15]), .ip2(
        n10357), .op(n10358) );
  nor2_1 U12320 ( .ip1(n10359), .ip2(n10358), .op(n4396) );
  xor2_1 U12321 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[11]), .ip2(n6224), .op(n10360)
         );
  xor2_1 U12322 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[8]), .ip2(i_ssi_baudr[8]), .op(
        n10363) );
  nor2_1 U12323 ( .ip1(n5256), .ip2(n10380), .op(n10362) );
  xor2_1 U12324 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[13]), .ip2(i_ssi_baudr[13]), 
        .op(n10364) );
  xor2_1 U12325 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[15]), .ip2(i_ssi_baudr[15]), 
        .op(n10368) );
  xor2_1 U12326 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[12]), .ip2(i_ssi_baudr[12]), 
        .op(n10377) );
  xnor2_1 U12327 ( .ip1(n10377), .ip2(n10376), .op(n10394) );
  xor2_1 U12328 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[10]), .ip2(n5257), .op(n10379)
         );
  xor2_1 U12329 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[7]), .ip2(n5256), .op(n10381)
         );
  inv_1 U12330 ( .ip(i_ssi_U_sclkgen_ssi_cnt[4]), .op(n10441) );
  xor2_2 U12331 ( .ip1(n10383), .ip2(n10382), .op(n10390) );
  fulladder U12332 ( .a(i_ssi_U_sclkgen_ssi_cnt[2]), .b(n10385), .ci(n10384), 
        .s(n10387) );
  xor2_1 U12333 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[1]), .ip2(n10385), .op(n10386)
         );
  xor2_1 U12334 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[9]), .ip2(n11652), .op(n10396)
         );
  xor2_1 U12335 ( .ip1(n10396), .ip2(n10395), .op(n10400) );
  xor2_1 U12336 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[5]), .ip2(i_ssi_baudr[5]), .op(
        n10398) );
  xor2_1 U12337 ( .ip1(n10398), .ip2(n10397), .op(n10399) );
  xor2_1 U12338 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[6]), .ip2(i_ssi_baudr[6]), .op(
        n10402) );
  xor2_1 U12339 ( .ip1(n10402), .ip2(n10401), .op(n10403) );
  nor2_1 U12340 ( .ip1(n11148), .ip2(n10409), .op(i_ssi_U_sclkgen_N75) );
  nand2_1 U12341 ( .ip1(i_apb_paddr[28]), .ip2(n11497), .op(n10412) );
  nand2_1 U12342 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[28]), .ip2(n11507), 
        .op(n10411) );
  nand2_1 U12343 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[28]), .ip2(n5269), 
        .op(n10410) );
  nand3_1 U12344 ( .ip1(n10412), .ip2(n10411), .ip3(n10410), .op(n4711) );
  nand2_1 U12345 ( .ip1(n10414), .ip2(n10413), .op(
        i_i2c_U_DW_apb_i2c_mstfsm_N421) );
  nor2_1 U12346 ( .ip1(i_i2c_mst_rx_bwen), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_mst_tx_bwen), .op(n10415) );
  nor4_1 U12347 ( .ip1(n11776), .ip2(n11774), .ip3(
        i_i2c_U_DW_apb_i2c_toggle_N30), .ip4(n10415), .op(
        i_i2c_U_DW_apb_i2c_tx_shift_byte_wait_en) );
  and4_1 U12348 ( .ip1(n11776), .ip2(i_i2c_U_DW_apb_i2c_rx_filter_sda_int_q), 
        .ip3(i_i2c_U_DW_apb_i2c_rx_filter_scl_int_q), .ip4(n10579), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_s_det_int) );
  nand2_1 U12349 ( .ip1(n5386), .ip2(n5307), .op(n10418) );
  nand3_1 U12350 ( .ip1(n5307), .ip2(i_ssi_U_sclkgen_ssi_cnt[0]), .ip3(n10416), 
        .op(n10417) );
  nand2_1 U12351 ( .ip1(n10418), .ip2(n10417), .op(i_ssi_U_sclkgen_N41) );
  inv_1 U12352 ( .ip(i_ssi_U_sclkgen_ssi_cnt[13]), .op(n10467) );
  inv_1 U12353 ( .ip(i_ssi_U_sclkgen_ssi_cnt[9]), .op(n10455) );
  inv_1 U12354 ( .ip(i_ssi_U_sclkgen_ssi_cnt[5]), .op(n10443) );
  nand2_1 U12355 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[1]), .ip2(
        i_ssi_U_sclkgen_ssi_cnt[0]), .op(n10432) );
  and2_1 U12356 ( .ip1(n10434), .ip2(i_ssi_U_sclkgen_ssi_cnt[3]), .op(n10438)
         );
  nand2_1 U12357 ( .ip1(n10438), .ip2(i_ssi_U_sclkgen_ssi_cnt[4]), .op(n10442)
         );
  nand2_1 U12358 ( .ip1(n10444), .ip2(i_ssi_U_sclkgen_ssi_cnt[6]), .op(n10448)
         );
  nand2_1 U12359 ( .ip1(n10450), .ip2(i_ssi_U_sclkgen_ssi_cnt[8]), .op(n10454)
         );
  nand2_1 U12360 ( .ip1(n10456), .ip2(i_ssi_U_sclkgen_ssi_cnt[10]), .op(n10460) );
  nand2_1 U12361 ( .ip1(n10462), .ip2(i_ssi_U_sclkgen_ssi_cnt[12]), .op(n10466) );
  nand2_1 U12362 ( .ip1(n10468), .ip2(i_ssi_U_sclkgen_ssi_cnt[14]), .op(n10469) );
  xor2_1 U12363 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[15]), .ip2(n10469), .op(n10419)
         );
  and2_1 U12364 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[14]), 
        .ip2(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[13]), .op(n10420) );
  nand2_1 U12365 ( .ip1(n10420), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[12]), .op(n10430) );
  and2_1 U12366 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[10]), 
        .ip2(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[11]), .op(n10429) );
  inv_1 U12367 ( .ip(n10423), .op(n10426) );
  not_ab_or_c_or_d U12368 ( .ip1(n10427), .ip2(n10426), .ip3(n10425), .ip4(
        n10424), .op(n11063) );
  nand4_1 U12369 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[6]), 
        .ip2(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[5]), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[4]), .ip4(n11063), .op(
        n10428) );
  nor2_2 U12370 ( .ip1(n11065), .ip2(n10428), .op(n11077) );
  nand2_2 U12371 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[7]), 
        .ip2(n11077), .op(n11081) );
  nand2_2 U12372 ( .ip1(n10429), .ip2(n11084), .op(n11093) );
  nor2_1 U12373 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[15]), 
        .ip2(n5446), .op(n10431) );
  nor2_1 U12374 ( .ip1(n10431), .ip2(n11099), .op(n4942) );
  not_ab_or_c_or_d U12375 ( .ip1(n10433), .ip2(n10432), .ip3(n10434), .ip4(
        n10435), .op(i_ssi_U_sclkgen_N42) );
  inv_1 U12376 ( .ip(i_ssi_U_sclkgen_ssi_cnt[3]), .op(n10437) );
  not_ab_or_c_or_d U12377 ( .ip1(n10437), .ip2(n10436), .ip3(n10438), .ip4(
        n5391), .op(i_ssi_U_sclkgen_N43) );
  inv_1 U12378 ( .ip(n10438), .op(n10440) );
  inv_1 U12379 ( .ip(n10442), .op(n10439) );
  not_ab_or_c_or_d U12380 ( .ip1(n10441), .ip2(n10440), .ip3(n10439), .ip4(
        n10435), .op(i_ssi_U_sclkgen_N44) );
  not_ab_or_c_or_d U12381 ( .ip1(n10443), .ip2(n10442), .ip3(n10444), .ip4(
        n5391), .op(i_ssi_U_sclkgen_N45) );
  inv_1 U12382 ( .ip(i_ssi_U_sclkgen_ssi_cnt[6]), .op(n10447) );
  inv_1 U12383 ( .ip(n10448), .op(n10445) );
  not_ab_or_c_or_d U12384 ( .ip1(n10447), .ip2(n10446), .ip3(n10445), .ip4(
        n5391), .op(i_ssi_U_sclkgen_N46) );
  not_ab_or_c_or_d U12385 ( .ip1(n10449), .ip2(n10448), .ip3(n10450), .ip4(
        n10435), .op(i_ssi_U_sclkgen_N47) );
  inv_1 U12386 ( .ip(n10454), .op(n10451) );
  not_ab_or_c_or_d U12387 ( .ip1(n10453), .ip2(n10452), .ip3(n10451), .ip4(
        n10435), .op(i_ssi_U_sclkgen_N48) );
  not_ab_or_c_or_d U12388 ( .ip1(n10455), .ip2(n10454), .ip3(n10456), .ip4(
        n10435), .op(i_ssi_U_sclkgen_N49) );
  not_ab_or_c_or_d U12389 ( .ip1(n10459), .ip2(n10458), .ip3(n5391), .ip4(
        n10457), .op(i_ssi_U_sclkgen_N50) );
  not_ab_or_c_or_d U12390 ( .ip1(n10461), .ip2(n10460), .ip3(n5391), .ip4(
        n10462), .op(i_ssi_U_sclkgen_N51) );
  not_ab_or_c_or_d U12391 ( .ip1(n10465), .ip2(n10464), .ip3(n5391), .ip4(
        n10463), .op(i_ssi_U_sclkgen_N52) );
  not_ab_or_c_or_d U12392 ( .ip1(n10467), .ip2(n10466), .ip3(n10435), .ip4(
        n10468), .op(i_ssi_U_sclkgen_N53) );
  inv_1 U12393 ( .ip(i_ssi_U_sclkgen_ssi_cnt[14]), .op(n10472) );
  inv_1 U12394 ( .ip(n10469), .op(n10470) );
  not_ab_or_c_or_d U12395 ( .ip1(n10472), .ip2(n10471), .ip3(n5391), .ip4(
        n10470), .op(i_ssi_U_sclkgen_N54) );
  nand2_1 U12396 ( .ip1(n10473), .ip2(i_ssi_U_mstfsm_bit_cnt[0]), .op(n10474)
         );
  not_ab_or_c_or_d U12397 ( .ip1(n10475), .ip2(n10474), .ip3(n10476), .ip4(
        n10480), .op(n4209) );
  inv_1 U12398 ( .ip(n10476), .op(n10478) );
  not_ab_or_c_or_d U12399 ( .ip1(n5565), .ip2(n10478), .ip3(n10477), .ip4(
        n10480), .op(n4208) );
  not_ab_or_c_or_d U12400 ( .ip1(n10482), .ip2(n10481), .ip3(n10480), .ip4(
        n10479), .op(n4207) );
  inv_1 U12401 ( .ip(i_ssi_U_mstfsm_frame_cnt[0]), .op(n10494) );
  nor2_1 U12402 ( .ip1(n10484), .ip2(n10483), .op(n10485) );
  nand2_1 U12403 ( .ip1(n10486), .ip2(n10485), .op(n10488) );
  inv_1 U12404 ( .ip(n10502), .op(n10491) );
  not_ab_or_c_or_d U12405 ( .ip1(n10494), .ip2(n10493), .ip3(n10542), .ip4(
        n10495), .op(n4184) );
  inv_1 U12406 ( .ip(n10495), .op(n10497) );
  nand2_1 U12407 ( .ip1(n10495), .ip2(i_ssi_U_mstfsm_frame_cnt[1]), .op(n10503) );
  inv_1 U12408 ( .ip(n10503), .op(n10496) );
  not_ab_or_c_or_d U12409 ( .ip1(n10498), .ip2(n10497), .ip3(n10542), .ip4(
        n10496), .op(n4185) );
  not_ab_or_c_or_d U12410 ( .ip1(n10504), .ip2(n10503), .ip3(n10516), .ip4(
        n10542), .op(n4186) );
  inv_1 U12411 ( .ip(n10516), .op(n10506) );
  nand2_1 U12412 ( .ip1(n10516), .ip2(i_ssi_U_mstfsm_frame_cnt[3]), .op(n10508) );
  inv_1 U12413 ( .ip(n10508), .op(n10505) );
  not_ab_or_c_or_d U12414 ( .ip1(n10507), .ip2(n10506), .ip3(n10542), .ip4(
        n10505), .op(n4187) );
  not_ab_or_c_or_d U12415 ( .ip1(n10509), .ip2(n10508), .ip3(n10542), .ip4(
        n10510), .op(n4188) );
  inv_1 U12416 ( .ip(n10510), .op(n10512) );
  nand2_1 U12417 ( .ip1(n10510), .ip2(i_ssi_U_mstfsm_frame_cnt[5]), .op(n10518) );
  inv_1 U12418 ( .ip(n10518), .op(n10511) );
  not_ab_or_c_or_d U12419 ( .ip1(n10513), .ip2(n10512), .ip3(n10542), .ip4(
        n10511), .op(n4189) );
  inv_1 U12420 ( .ip(n10514), .op(n10515) );
  nand2_1 U12421 ( .ip1(n10516), .ip2(n10515), .op(n10520) );
  inv_1 U12422 ( .ip(n10520), .op(n10517) );
  not_ab_or_c_or_d U12423 ( .ip1(n10519), .ip2(n10518), .ip3(n10517), .ip4(
        n10542), .op(n4190) );
  not_ab_or_c_or_d U12424 ( .ip1(n10521), .ip2(n10520), .ip3(n10542), .ip4(
        n10522), .op(n4191) );
  inv_1 U12425 ( .ip(n10522), .op(n10524) );
  nand2_1 U12426 ( .ip1(n10522), .ip2(i_ssi_U_mstfsm_frame_cnt[8]), .op(n10526) );
  inv_1 U12427 ( .ip(n10526), .op(n10523) );
  not_ab_or_c_or_d U12428 ( .ip1(n10525), .ip2(n10524), .ip3(n10542), .ip4(
        n10523), .op(n4192) );
  not_ab_or_c_or_d U12429 ( .ip1(n10527), .ip2(n10526), .ip3(n10528), .ip4(
        n10542), .op(n4193) );
  inv_1 U12430 ( .ip(n10528), .op(n10530) );
  inv_1 U12431 ( .ip(n10532), .op(n10529) );
  not_ab_or_c_or_d U12432 ( .ip1(n10531), .ip2(n10530), .ip3(n10542), .ip4(
        n10529), .op(n4194) );
  not_ab_or_c_or_d U12433 ( .ip1(n10533), .ip2(n10532), .ip3(n10542), .ip4(
        n10536), .op(n4195) );
  inv_1 U12434 ( .ip(n10538), .op(n10534) );
  not_ab_or_c_or_d U12435 ( .ip1(n10535), .ip2(n5278), .ip3(n10542), .ip4(
        n10534), .op(n4196) );
  not_ab_or_c_or_d U12436 ( .ip1(n10539), .ip2(n10538), .ip3(n10542), .ip4(
        n10540), .op(n4197) );
  nand2_1 U12437 ( .ip1(n10540), .ip2(i_ssi_U_mstfsm_frame_cnt[14]), .op(
        n10543) );
  not_ab_or_c_or_d U12438 ( .ip1(n10544), .ip2(n10543), .ip3(n10542), .ip4(
        n5425), .op(n4199) );
  nand2_1 U12439 ( .ip1(n10545), .ip2(i_ssi_U_regfile_txflr[0]), .op(n10546)
         );
  nor4_1 U12440 ( .ip1(i_ssi_U_regfile_txflr[3]), .ip2(
        i_ssi_U_regfile_txflr[2]), .ip3(n11780), .ip4(n10546), .op(n10549) );
  inv_1 U12441 ( .ip(i_ssi_U_fifo_U_tx_fifo_empty_n), .op(n10548) );
  not_ab_or_c_or_d U12442 ( .ip1(n10549), .ip2(i_ssi_tx_pop_sync), .ip3(n10548), .ip4(n10547), .op(i_ssi_U_regfile_N452) );
  not_ab_or_c_or_d U12443 ( .ip1(n10552), .ip2(n10551), .ip3(n10550), .ip4(
        n10561), .op(i_i2c_U_DW_apb_i2c_rx_filter_N84) );
  not_ab_or_c_or_d U12444 ( .ip1(n10554), .ip2(n10553), .ip3(n10555), .ip4(
        n10561), .op(i_i2c_U_DW_apb_i2c_rx_filter_N85) );
  inv_1 U12445 ( .ip(n10555), .op(n10557) );
  not_ab_or_c_or_d U12446 ( .ip1(n10558), .ip2(n10557), .ip3(n10556), .ip4(
        n10561), .op(i_i2c_U_DW_apb_i2c_rx_filter_N86) );
  not_ab_or_c_or_d U12447 ( .ip1(n5318), .ip2(n10559), .ip3(n10560), .ip4(
        n10561), .op(i_i2c_U_DW_apb_i2c_rx_filter_N87) );
  inv_1 U12448 ( .ip(n5316), .op(n10564) );
  inv_1 U12449 ( .ip(n10560), .op(n10563) );
  not_ab_or_c_or_d U12450 ( .ip1(n10564), .ip2(n10563), .ip3(n10562), .ip4(
        n10561), .op(i_i2c_U_DW_apb_i2c_rx_filter_N88) );
  nand2_1 U12451 ( .ip1(n11776), .ip2(n10565), .op(n10568) );
  not_ab_or_c_or_d U12452 ( .ip1(n10572), .ip2(n10568), .ip3(n10567), .ip4(
        n10566), .op(n5202) );
  nor2_1 U12453 ( .ip1(n10573), .ip2(i_i2c_mst_rx_bwen), .op(n10570) );
  not_ab_or_c_or_d U12454 ( .ip1(n10573), .ip2(n10572), .ip3(n10571), .ip4(
        n10570), .op(n4167) );
  nand2_1 U12455 ( .ip1(n10575), .ip2(n10574), .op(n10578) );
  inv_1 U12456 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_mst_tx_bwen), .op(n10577) );
  nor2_1 U12457 ( .ip1(i_i2c_scl_hcnt_en), .ip2(n10578), .op(n10576) );
  not_ab_or_c_or_d U12458 ( .ip1(n10578), .ip2(n10577), .ip3(n11173), .ip4(
        n10576), .op(n4134) );
  nor2_1 U12459 ( .ip1(n10579), .ip2(n11167), .op(n10581) );
  inv_1 U12460 ( .ip(i_i2c_mst_tx_ack_vld), .op(n10580) );
  not_ab_or_c_or_d U12461 ( .ip1(n10582), .ip2(n11167), .ip3(n10581), .ip4(
        n10580), .op(n4168) );
  inv_1 U12462 ( .ip(n10583), .op(n10587) );
  nor2_1 U12463 ( .ip1(n10584), .ip2(n10583), .op(n10585) );
  nor2_1 U12464 ( .ip1(i_i2c_scl_hcnt_en), .ip2(n10585), .op(n10586) );
  not_ab_or_c_or_d U12465 ( .ip1(n10587), .ip2(n11158), .ip3(n10586), .ip4(
        n11160), .op(n4149) );
  inv_1 U12466 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[0]), .op(n10588)
         );
  not_ab_or_c_or_d U12467 ( .ip1(n10589), .ip2(n10588), .ip3(n10590), .ip4(
        n10630), .op(n5185) );
  inv_1 U12468 ( .ip(n10590), .op(n10592) );
  inv_1 U12469 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[1]), .op(n10591)
         );
  not_ab_or_c_or_d U12470 ( .ip1(n10592), .ip2(n10591), .ip3(n10593), .ip4(
        n10630), .op(n5184) );
  inv_1 U12471 ( .ip(n10593), .op(n10595) );
  inv_1 U12472 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[2]), .op(n10594)
         );
  not_ab_or_c_or_d U12473 ( .ip1(n10595), .ip2(n10594), .ip3(n10596), .ip4(
        n10630), .op(n5183) );
  inv_1 U12474 ( .ip(n10596), .op(n10598) );
  inv_1 U12475 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[3]), .op(n10597)
         );
  not_ab_or_c_or_d U12476 ( .ip1(n10598), .ip2(n10597), .ip3(n10599), .ip4(
        n10630), .op(n5182) );
  inv_1 U12477 ( .ip(n10599), .op(n10601) );
  inv_1 U12478 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[4]), .op(n10600)
         );
  not_ab_or_c_or_d U12479 ( .ip1(n10601), .ip2(n10600), .ip3(n10602), .ip4(
        n10630), .op(n5181) );
  inv_1 U12480 ( .ip(n10602), .op(n10604) );
  inv_1 U12481 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[5]), .op(n10603)
         );
  not_ab_or_c_or_d U12482 ( .ip1(n10604), .ip2(n10603), .ip3(n10605), .ip4(
        n10630), .op(n5180) );
  inv_1 U12483 ( .ip(n10605), .op(n10607) );
  inv_1 U12484 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[6]), .op(n10606)
         );
  not_ab_or_c_or_d U12485 ( .ip1(n10607), .ip2(n10606), .ip3(n10608), .ip4(
        n10630), .op(n5179) );
  inv_1 U12486 ( .ip(n10608), .op(n10610) );
  inv_1 U12487 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[7]), .op(n10609)
         );
  not_ab_or_c_or_d U12488 ( .ip1(n10610), .ip2(n10609), .ip3(n10611), .ip4(
        n10630), .op(n5178) );
  inv_1 U12489 ( .ip(n10611), .op(n10613) );
  inv_1 U12490 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[8]), .op(n10612)
         );
  not_ab_or_c_or_d U12491 ( .ip1(n10613), .ip2(n10612), .ip3(n10614), .ip4(
        n10630), .op(n5177) );
  inv_1 U12492 ( .ip(n10614), .op(n10616) );
  inv_1 U12493 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[9]), .op(n10615)
         );
  not_ab_or_c_or_d U12494 ( .ip1(n10616), .ip2(n10615), .ip3(n10617), .ip4(
        n10630), .op(n5176) );
  inv_1 U12495 ( .ip(n10617), .op(n10619) );
  inv_1 U12496 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[10]), .op(n10618)
         );
  not_ab_or_c_or_d U12497 ( .ip1(n10619), .ip2(n10618), .ip3(n10620), .ip4(
        n10630), .op(n5175) );
  inv_1 U12498 ( .ip(n10620), .op(n10622) );
  inv_1 U12499 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[11]), .op(n10621)
         );
  not_ab_or_c_or_d U12500 ( .ip1(n10622), .ip2(n10621), .ip3(n10623), .ip4(
        n10630), .op(n5174) );
  inv_1 U12501 ( .ip(n10623), .op(n10625) );
  inv_1 U12502 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[12]), .op(n10624)
         );
  not_ab_or_c_or_d U12503 ( .ip1(n10625), .ip2(n10624), .ip3(n10626), .ip4(
        n10630), .op(n5173) );
  inv_1 U12504 ( .ip(n10626), .op(n10628) );
  inv_1 U12505 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[13]), .op(n10627)
         );
  not_ab_or_c_or_d U12506 ( .ip1(n10628), .ip2(n10627), .ip3(n10629), .ip4(
        n10630), .op(n5172) );
  inv_1 U12507 ( .ip(n10629), .op(n10633) );
  inv_1 U12508 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[14]), .op(n10632)
         );
  not_ab_or_c_or_d U12509 ( .ip1(n10633), .ip2(n10632), .ip3(n10631), .ip4(
        n10630), .op(n5171) );
  inv_1 U12510 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[0]), .op(
        n10635) );
  and2_1 U12511 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[0]), .ip2(
        n10634), .op(n10637) );
  not_ab_or_c_or_d U12512 ( .ip1(n10636), .ip2(n10635), .ip3(n10637), .ip4(
        n10677), .op(n5066) );
  inv_1 U12513 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[1]), .op(
        n10640) );
  inv_1 U12514 ( .ip(n10637), .op(n10639) );
  nand2_1 U12515 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[1]), .ip2(
        n10637), .op(n10641) );
  inv_1 U12516 ( .ip(n10641), .op(n10638) );
  not_ab_or_c_or_d U12517 ( .ip1(n10640), .ip2(n10639), .ip3(n10638), .ip4(
        n10677), .op(n5065) );
  inv_1 U12518 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[2]), .op(
        n10642) );
  not_ab_or_c_or_d U12519 ( .ip1(n10642), .ip2(n10641), .ip3(n10643), .ip4(
        n10677), .op(n5064) );
  inv_1 U12520 ( .ip(n10643), .op(n10646) );
  inv_1 U12521 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[3]), .op(
        n10645) );
  inv_1 U12522 ( .ip(n10648), .op(n10644) );
  not_ab_or_c_or_d U12523 ( .ip1(n10646), .ip2(n10645), .ip3(n10644), .ip4(
        n10677), .op(n5063) );
  not_ab_or_c_or_d U12524 ( .ip1(n10648), .ip2(n10647), .ip3(n10649), .ip4(
        n10677), .op(n5062) );
  inv_1 U12525 ( .ip(n10649), .op(n10652) );
  inv_1 U12526 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[5]), .op(
        n10651) );
  inv_1 U12527 ( .ip(n10654), .op(n10650) );
  not_ab_or_c_or_d U12528 ( .ip1(n10652), .ip2(n10651), .ip3(n10650), .ip4(
        n10677), .op(n5061) );
  not_ab_or_c_or_d U12529 ( .ip1(n10654), .ip2(n10653), .ip3(n10655), .ip4(
        n10677), .op(n5060) );
  inv_1 U12530 ( .ip(n10655), .op(n10658) );
  inv_1 U12531 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[7]), .op(
        n10657) );
  inv_1 U12532 ( .ip(n10660), .op(n10656) );
  not_ab_or_c_or_d U12533 ( .ip1(n10658), .ip2(n10657), .ip3(n10656), .ip4(
        n10677), .op(n5059) );
  not_ab_or_c_or_d U12534 ( .ip1(n10660), .ip2(n10659), .ip3(n10661), .ip4(
        n10677), .op(n5058) );
  inv_1 U12535 ( .ip(n10661), .op(n10664) );
  inv_1 U12536 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[9]), .op(
        n10663) );
  inv_1 U12537 ( .ip(n10666), .op(n10662) );
  not_ab_or_c_or_d U12538 ( .ip1(n10664), .ip2(n10663), .ip3(n10662), .ip4(
        n10677), .op(n5057) );
  not_ab_or_c_or_d U12539 ( .ip1(n10666), .ip2(n10665), .ip3(n10667), .ip4(
        n10677), .op(n5056) );
  inv_1 U12540 ( .ip(n10667), .op(n10670) );
  inv_1 U12541 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[11]), .op(
        n10669) );
  inv_1 U12542 ( .ip(n10672), .op(n10668) );
  not_ab_or_c_or_d U12543 ( .ip1(n10670), .ip2(n10669), .ip3(n10668), .ip4(
        n10677), .op(n5055) );
  not_ab_or_c_or_d U12544 ( .ip1(n10672), .ip2(n10671), .ip3(n10673), .ip4(
        n10677), .op(n5054) );
  inv_1 U12545 ( .ip(n10673), .op(n10676) );
  inv_1 U12546 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[13]), .op(
        n10675) );
  inv_1 U12547 ( .ip(n10680), .op(n10674) );
  not_ab_or_c_or_d U12548 ( .ip1(n10676), .ip2(n10675), .ip3(n10674), .ip4(
        n10677), .op(n5053) );
  not_ab_or_c_or_d U12549 ( .ip1(n10680), .ip2(n10679), .ip3(n10678), .ip4(
        n10677), .op(n5052) );
  nand2_1 U12550 ( .ip1(i_i2c_ic_fs_lcnt[13]), .ip2(n10719), .op(n10682) );
  inv_4 U12551 ( .ip(n10719), .op(n10720) );
  nand2_1 U12552 ( .ip1(i_i2c_ic_lcnt[13]), .ip2(n10720), .op(n10681) );
  nand2_1 U12553 ( .ip1(i_i2c_ic_fs_lcnt[2]), .ip2(n10719), .op(n10688) );
  nand2_1 U12554 ( .ip1(i_i2c_ic_lcnt[2]), .ip2(n10720), .op(n10687) );
  nand2_1 U12555 ( .ip1(i_i2c_ic_fs_lcnt[3]), .ip2(n10719), .op(n10690) );
  nand2_1 U12556 ( .ip1(i_i2c_ic_lcnt[3]), .ip2(n10720), .op(n10689) );
  nand2_1 U12557 ( .ip1(i_i2c_ic_fs_lcnt[4]), .ip2(n10719), .op(n10692) );
  nand2_1 U12558 ( .ip1(i_i2c_ic_lcnt[4]), .ip2(n10720), .op(n10691) );
  nand2_1 U12559 ( .ip1(i_i2c_ic_fs_lcnt[5]), .ip2(n10719), .op(n10694) );
  nand2_1 U12560 ( .ip1(i_i2c_ic_lcnt[5]), .ip2(n10720), .op(n10693) );
  nand2_1 U12561 ( .ip1(i_i2c_ic_fs_lcnt[6]), .ip2(n10719), .op(n10696) );
  nand2_1 U12562 ( .ip1(i_i2c_ic_lcnt[6]), .ip2(n10720), .op(n10695) );
  nand2_1 U12563 ( .ip1(i_i2c_ic_fs_lcnt[7]), .ip2(n10719), .op(n10698) );
  nand2_1 U12564 ( .ip1(i_i2c_ic_lcnt[7]), .ip2(n10720), .op(n10697) );
  nand2_1 U12565 ( .ip1(i_i2c_ic_fs_lcnt[8]), .ip2(n10719), .op(n10700) );
  nand2_1 U12566 ( .ip1(i_i2c_ic_lcnt[8]), .ip2(n10720), .op(n10699) );
  nand2_1 U12567 ( .ip1(i_i2c_ic_fs_lcnt[9]), .ip2(n10719), .op(n10702) );
  nand2_1 U12568 ( .ip1(i_i2c_ic_lcnt[9]), .ip2(n10720), .op(n10701) );
  nand2_1 U12569 ( .ip1(i_i2c_ic_fs_lcnt[10]), .ip2(n10719), .op(n10704) );
  nand2_1 U12570 ( .ip1(i_i2c_ic_lcnt[10]), .ip2(n10720), .op(n10703) );
  nand2_1 U12571 ( .ip1(i_i2c_ic_fs_lcnt[11]), .ip2(n10719), .op(n10706) );
  nand2_1 U12572 ( .ip1(i_i2c_ic_lcnt[11]), .ip2(n10720), .op(n10705) );
  nand2_1 U12573 ( .ip1(i_i2c_ic_fs_lcnt[12]), .ip2(n10719), .op(n10708) );
  nand2_1 U12574 ( .ip1(i_i2c_ic_lcnt[12]), .ip2(n10720), .op(n10707) );
  xor2_1 U12575 ( .ip1(n10717), .ip2(n10718), .op(n10907) );
  inv_1 U12576 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[12]), .op(n10779) );
  xor2_1 U12577 ( .ip1(n10710), .ip2(n10709), .op(n10837) );
  nor2_1 U12578 ( .ip1(n10711), .ip2(n10712), .op(n10714) );
  nor2_1 U12579 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[13]), .ip2(
        n10712), .op(n10713) );
  or2_1 U12580 ( .ip1(n10714), .ip2(n10713), .op(n10729) );
  nand2_1 U12581 ( .ip1(i_i2c_ic_fs_lcnt[14]), .ip2(n10719), .op(n10716) );
  nand2_1 U12582 ( .ip1(i_i2c_ic_lcnt[14]), .ip2(n10720), .op(n10715) );
  inv_1 U12583 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[14]), .op(n10732) );
  nand2_2 U12584 ( .ip1(n10835), .ip2(n10732), .op(n10728) );
  nand2_1 U12585 ( .ip1(i_i2c_ic_fs_lcnt[15]), .ip2(n10719), .op(n10722) );
  nand2_1 U12586 ( .ip1(i_i2c_ic_lcnt[15]), .ip2(n10720), .op(n10721) );
  xor2_1 U12587 ( .ip1(n10726), .ip2(n10725), .op(n10917) );
  inv_1 U12588 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[15]), .op(n10727) );
  nand2_1 U12589 ( .ip1(n10728), .ip2(n10730), .op(n10778) );
  nor2_1 U12590 ( .ip1(n10729), .ip2(n10778), .op(n10799) );
  inv_1 U12591 ( .ip(n10730), .op(n10731) );
  nor2_2 U12592 ( .ip1(n10917), .ip2(n10727), .op(n10914) );
  xor2_1 U12593 ( .ip1(n10734), .ip2(n10733), .op(n10887) );
  inv_2 U12594 ( .ip(n10887), .op(n10783) );
  nor2_1 U12595 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[9]), .ip2(
        n10783), .op(n10781) );
  xor2_1 U12596 ( .ip1(n10736), .ip2(n10735), .op(n10875) );
  inv_1 U12597 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[6]), .op(n10765)
         );
  xor2_1 U12598 ( .ip1(n10738), .ip2(n10737), .op(n10870) );
  nor2_1 U12599 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[7]), .ip2(
        n5276), .op(n10763) );
  xor2_1 U12600 ( .ip1(n10740), .ip2(n10739), .op(n10865) );
  inv_1 U12601 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[4]), .op(n10759)
         );
  nor2_1 U12602 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[5]), .ip2(
        n10762), .op(n10758) );
  xor2_1 U12603 ( .ip1(n10742), .ip2(n10741), .op(n10859) );
  nor3_1 U12604 ( .ip1(n10759), .ip2(n10758), .ip3(n10859), .op(n10761) );
  xor2_1 U12605 ( .ip1(n10744), .ip2(n10743), .op(n10854) );
  xor2_1 U12606 ( .ip1(n10746), .ip2(n10745), .op(n10848) );
  inv_1 U12607 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[2]), .op(n10754)
         );
  and2_1 U12608 ( .ip1(n10848), .ip2(n10754), .op(n10752) );
  nor2_1 U12609 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[3]), .ip2(
        n5280), .op(n10753) );
  xor2_1 U12610 ( .ip1(n10747), .ip2(n10748), .op(n10843) );
  inv_1 U12611 ( .ip(n10748), .op(n10841) );
  not_ab_or_c_or_d U12612 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[1]), 
        .ip2(n10749), .ip3(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[0]), .ip4(
        n10748), .op(n10751) );
  nor2_1 U12613 ( .ip1(n10749), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[1]), .op(n10750) );
  nor4_1 U12614 ( .ip1(n10752), .ip2(n10753), .ip3(n10751), .ip4(n10750), .op(
        n10756) );
  nor3_1 U12615 ( .ip1(n10754), .ip2(n10753), .ip3(n10848), .op(n10755) );
  not_ab_or_c_or_d U12616 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[3]), 
        .ip2(n5280), .ip3(n10756), .ip4(n10755), .op(n10757) );
  not_ab_or_c_or_d U12617 ( .ip1(n10859), .ip2(n10759), .ip3(n10758), .ip4(
        n10757), .op(n10760) );
  not_ab_or_c_or_d U12618 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[5]), 
        .ip2(n10762), .ip3(n10761), .ip4(n10760), .op(n10764) );
  not_ab_or_c_or_d U12619 ( .ip1(n10870), .ip2(n10765), .ip3(n10764), .ip4(
        n10763), .op(n10766) );
  not_ab_or_c_or_d U12620 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[7]), 
        .ip2(n5276), .ip3(n10767), .ip4(n10766), .op(n10776) );
  xor2_1 U12621 ( .ip1(n10769), .ip2(n10768), .op(n10881) );
  inv_1 U12622 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[8]), .op(n10782)
         );
  xor2_1 U12623 ( .ip1(n10771), .ip2(n10770), .op(n10891) );
  inv_1 U12624 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[10]), .op(n10890) );
  nand2_1 U12625 ( .ip1(n10891), .ip2(n10890), .op(n10894) );
  xor2_1 U12626 ( .ip1(n10773), .ip2(n10772), .op(n10899) );
  nor2_1 U12627 ( .ip1(n10792), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[11]), .op(n10789) );
  inv_1 U12628 ( .ip(n10789), .op(n10774) );
  or4_1 U12629 ( .ip1(n10781), .ip2(n10776), .ip3(n10775), .ip4(n10787), .op(
        n10780) );
  ab_or_c_or_d U12630 ( .ip1(n10837), .ip2(n10779), .ip3(n10778), .ip4(n10777), 
        .op(n10793) );
  nor2_1 U12631 ( .ip1(n10780), .ip2(n10793), .op(n10796) );
  nor2_1 U12632 ( .ip1(n10783), .ip2(n10784), .op(n10786) );
  nor2_1 U12633 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[9]), .ip2(
        n10784), .op(n10785) );
  or2_1 U12634 ( .ip1(n10786), .ip2(n10785), .op(n10788) );
  nor2_1 U12635 ( .ip1(n10788), .ip2(n10787), .op(n10791) );
  nor3_2 U12636 ( .ip1(n10890), .ip2(n10891), .ip3(n10789), .op(n10790) );
  not_ab_or_c_or_d U12637 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[11]), 
        .ip2(n10792), .ip3(n10791), .ip4(n10790), .op(n10794) );
  nor2_1 U12638 ( .ip1(n10794), .ip2(n10793), .op(n10795) );
  or2_1 U12639 ( .ip1(n10796), .ip2(n10795), .op(n10797) );
  inv_1 U12640 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[3]), .op(n10853)
         );
  inv_1 U12641 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[5]), .op(n10864)
         );
  inv_1 U12642 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[7]), .op(n10838)
         );
  inv_1 U12643 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[9]), .op(n10886)
         );
  inv_1 U12644 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[11]), .op(n10898) );
  inv_1 U12645 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[13]), .op(n10906) );
  inv_1 U12646 ( .ip(n10808), .op(n10805) );
  nor2_1 U12647 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[15]), .ip2(
        n10804), .op(n10803) );
  nand3_1 U12648 ( .ip1(i_i2c_ic_enable_sync), .ip2(n10802), .ip3(n10801), 
        .op(n10833) );
  nor2_1 U12649 ( .ip1(n10803), .ip2(n10833), .op(
        i_i2c_U_DW_apb_i2c_clk_gen_N77) );
  not_ab_or_c_or_d U12650 ( .ip1(n10805), .ip2(n10732), .ip3(n10804), .ip4(
        n10833), .op(i_i2c_U_DW_apb_i2c_clk_gen_N76) );
  inv_1 U12651 ( .ip(n10810), .op(n10807) );
  inv_1 U12652 ( .ip(n10809), .op(n10806) );
  not_ab_or_c_or_d U12653 ( .ip1(n10807), .ip2(n10779), .ip3(n10833), .ip4(
        n10806), .op(i_i2c_U_DW_apb_i2c_clk_gen_N74) );
  not_ab_or_c_or_d U12654 ( .ip1(n10809), .ip2(n10906), .ip3(n10808), .ip4(
        n10833), .op(i_i2c_U_DW_apb_i2c_clk_gen_N75) );
  not_ab_or_c_or_d U12655 ( .ip1(n10812), .ip2(n10898), .ip3(n10810), .ip4(
        n10833), .op(i_i2c_U_DW_apb_i2c_clk_gen_N73) );
  not_ab_or_c_or_d U12656 ( .ip1(n10816), .ip2(n10886), .ip3(n10811), .ip4(
        n10833), .op(i_i2c_U_DW_apb_i2c_clk_gen_N71) );
  not_ab_or_c_or_d U12657 ( .ip1(n10820), .ip2(n10838), .ip3(n10815), .ip4(
        n10833), .op(i_i2c_U_DW_apb_i2c_clk_gen_N69) );
  not_ab_or_c_or_d U12658 ( .ip1(n10824), .ip2(n10864), .ip3(n10819), .ip4(
        n10833), .op(i_i2c_U_DW_apb_i2c_clk_gen_N67) );
  not_ab_or_c_or_d U12659 ( .ip1(n10831), .ip2(n10853), .ip3(n10823), .ip4(
        n10833), .op(i_i2c_U_DW_apb_i2c_clk_gen_N65) );
  inv_1 U12660 ( .ip(n10811), .op(n10814) );
  inv_1 U12661 ( .ip(n10812), .op(n10813) );
  not_ab_or_c_or_d U12662 ( .ip1(n10814), .ip2(n10890), .ip3(n10833), .ip4(
        n10813), .op(i_i2c_U_DW_apb_i2c_clk_gen_N72) );
  inv_1 U12663 ( .ip(n10815), .op(n10818) );
  inv_1 U12664 ( .ip(n10816), .op(n10817) );
  not_ab_or_c_or_d U12665 ( .ip1(n10818), .ip2(n10782), .ip3(n10833), .ip4(
        n10817), .op(i_i2c_U_DW_apb_i2c_clk_gen_N70) );
  inv_1 U12666 ( .ip(n10819), .op(n10822) );
  inv_1 U12667 ( .ip(n10820), .op(n10821) );
  not_ab_or_c_or_d U12668 ( .ip1(n10822), .ip2(n10765), .ip3(n10833), .ip4(
        n10821), .op(i_i2c_U_DW_apb_i2c_clk_gen_N68) );
  inv_1 U12669 ( .ip(n10823), .op(n10826) );
  inv_1 U12670 ( .ip(n10824), .op(n10825) );
  not_ab_or_c_or_d U12671 ( .ip1(n10826), .ip2(n10759), .ip3(n10833), .ip4(
        n10825), .op(i_i2c_U_DW_apb_i2c_clk_gen_N66) );
  inv_1 U12672 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[0]), .op(n10840)
         );
  nand2_1 U12673 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_count_en), .ip2(n5450), 
        .op(n10827) );
  not_ab_or_c_or_d U12674 ( .ip1(n10840), .ip2(n10827), .ip3(n10828), .ip4(
        n10833), .op(i_i2c_U_DW_apb_i2c_clk_gen_N62) );
  inv_1 U12675 ( .ip(n10828), .op(n10829) );
  inv_1 U12676 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[1]), .op(n10842)
         );
  not_ab_or_c_or_d U12677 ( .ip1(n10829), .ip2(n10842), .ip3(n10830), .ip4(
        n10833), .op(i_i2c_U_DW_apb_i2c_clk_gen_N63) );
  inv_1 U12678 ( .ip(n10830), .op(n10834) );
  inv_1 U12679 ( .ip(n10831), .op(n10832) );
  not_ab_or_c_or_d U12680 ( .ip1(n10834), .ip2(n10754), .ip3(n10833), .ip4(
        n10832), .op(i_i2c_U_DW_apb_i2c_clk_gen_N64) );
  nor2_1 U12681 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[14]), .ip2(
        n10910), .op(n10912) );
  nor2_1 U12682 ( .ip1(n10907), .ip2(n10906), .op(n10909) );
  inv_1 U12683 ( .ip(n10837), .op(n10836) );
  nor2_1 U12684 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[12]), .ip2(
        n10836), .op(n10905) );
  nor2_1 U12685 ( .ip1(n10837), .ip2(n10779), .op(n10903) );
  or2_1 U12686 ( .ip1(n10899), .ip2(n10898), .op(n10897) );
  or2_1 U12687 ( .ip1(n10887), .ip2(n10886), .op(n10885) );
  nor2_1 U12688 ( .ip1(n10875), .ip2(n10838), .op(n10874) );
  or2_1 U12689 ( .ip1(n10865), .ip2(n10864), .op(n10863) );
  nand2_1 U12690 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[3]), .ip2(
        n5280), .op(n10852) );
  or2_1 U12691 ( .ip1(n10848), .ip2(n10754), .op(n10847) );
  nand2_1 U12692 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[1]), .ip2(
        n10749), .op(n10839) );
  nand3_1 U12693 ( .ip1(n10841), .ip2(n10840), .ip3(n10839), .op(n10845) );
  nand2_1 U12694 ( .ip1(n10843), .ip2(n10842), .op(n10844) );
  nand2_1 U12695 ( .ip1(n10845), .ip2(n10844), .op(n10846) );
  nand2_1 U12696 ( .ip1(n10847), .ip2(n10846), .op(n10850) );
  nand2_1 U12697 ( .ip1(n10848), .ip2(n10754), .op(n10849) );
  nand2_1 U12698 ( .ip1(n10850), .ip2(n10849), .op(n10851) );
  nand2_1 U12699 ( .ip1(n10852), .ip2(n10851), .op(n10856) );
  nand2_1 U12700 ( .ip1(n10854), .ip2(n10853), .op(n10855) );
  nand2_1 U12701 ( .ip1(n10856), .ip2(n10855), .op(n10858) );
  or2_1 U12702 ( .ip1(n10859), .ip2(n10759), .op(n10857) );
  nand2_1 U12703 ( .ip1(n10858), .ip2(n10857), .op(n10861) );
  nand2_1 U12704 ( .ip1(n10859), .ip2(n10759), .op(n10860) );
  nand2_1 U12705 ( .ip1(n10861), .ip2(n10860), .op(n10862) );
  nand2_1 U12706 ( .ip1(n10863), .ip2(n10862), .op(n10867) );
  nand2_1 U12707 ( .ip1(n10865), .ip2(n10864), .op(n10866) );
  nand2_1 U12708 ( .ip1(n10867), .ip2(n10866), .op(n10869) );
  or2_1 U12709 ( .ip1(n10870), .ip2(n10765), .op(n10868) );
  nand2_1 U12710 ( .ip1(n10869), .ip2(n10868), .op(n10872) );
  nand2_1 U12711 ( .ip1(n10870), .ip2(n10765), .op(n10871) );
  and2_1 U12712 ( .ip1(n10872), .ip2(n10871), .op(n10873) );
  nor2_1 U12713 ( .ip1(n10874), .ip2(n10873), .op(n10877) );
  nor2_1 U12714 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[7]), .ip2(
        n5276), .op(n10876) );
  or2_1 U12715 ( .ip1(n10877), .ip2(n10876), .op(n10880) );
  inv_1 U12716 ( .ip(n10881), .op(n10878) );
  nand2_1 U12717 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[8]), .ip2(
        n10878), .op(n10879) );
  nand2_1 U12718 ( .ip1(n10880), .ip2(n10879), .op(n10883) );
  nand2_1 U12719 ( .ip1(n10881), .ip2(n10782), .op(n10882) );
  nand2_1 U12720 ( .ip1(n10883), .ip2(n10882), .op(n10884) );
  nand2_1 U12721 ( .ip1(n10885), .ip2(n10884), .op(n10889) );
  nand2_1 U12722 ( .ip1(n10887), .ip2(n10886), .op(n10888) );
  nand2_1 U12723 ( .ip1(n10889), .ip2(n10888), .op(n10893) );
  or2_1 U12724 ( .ip1(n10891), .ip2(n10890), .op(n10892) );
  nand2_1 U12725 ( .ip1(n10893), .ip2(n10892), .op(n10895) );
  nand2_1 U12726 ( .ip1(n10895), .ip2(n10894), .op(n10896) );
  nand2_1 U12727 ( .ip1(n10897), .ip2(n10896), .op(n10901) );
  nand2_1 U12728 ( .ip1(n10899), .ip2(n10898), .op(n10900) );
  and2_1 U12729 ( .ip1(n10901), .ip2(n10900), .op(n10902) );
  nor2_1 U12730 ( .ip1(n10903), .ip2(n10902), .op(n10904) );
  not_ab_or_c_or_d U12731 ( .ip1(n10907), .ip2(n10906), .ip3(n10905), .ip4(
        n10904), .op(n10908) );
  not_ab_or_c_or_d U12732 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[14]), 
        .ip2(n10910), .ip3(n10909), .ip4(n10908), .op(n10911) );
  not_ab_or_c_or_d U12733 ( .ip1(n10917), .ip2(n10727), .ip3(n10916), .ip4(
        n10915), .op(i_i2c_U_DW_apb_i2c_clk_gen_N51) );
  inv_1 U12734 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[0]), .op(n10919)
         );
  and2_1 U12735 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[0]), .ip2(
        n10918), .op(n10921) );
  not_ab_or_c_or_d U12736 ( .ip1(n10920), .ip2(n10919), .ip3(n10921), .ip4(
        n10955), .op(n5134) );
  inv_1 U12737 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[1]), .op(n10924)
         );
  inv_1 U12738 ( .ip(n10921), .op(n10923) );
  nand2_1 U12739 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[1]), .ip2(
        n10921), .op(n10925) );
  inv_1 U12740 ( .ip(n10925), .op(n10922) );
  not_ab_or_c_or_d U12741 ( .ip1(n10924), .ip2(n10923), .ip3(n10922), .ip4(
        n10955), .op(n5133) );
  not_ab_or_c_or_d U12742 ( .ip1(n7951), .ip2(n10925), .ip3(n10926), .ip4(
        n10955), .op(n5132) );
  inv_1 U12743 ( .ip(n10926), .op(n10929) );
  inv_1 U12744 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[3]), .op(n10928)
         );
  inv_1 U12745 ( .ip(n10930), .op(n10927) );
  not_ab_or_c_or_d U12746 ( .ip1(n10929), .ip2(n10928), .ip3(n10927), .ip4(
        n10955), .op(n5131) );
  not_ab_or_c_or_d U12747 ( .ip1(n10930), .ip2(n7957), .ip3(n10931), .ip4(
        n10955), .op(n5130) );
  inv_1 U12748 ( .ip(n10931), .op(n10934) );
  inv_1 U12749 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[5]), .op(n10933)
         );
  inv_1 U12750 ( .ip(n10935), .op(n10932) );
  not_ab_or_c_or_d U12751 ( .ip1(n10934), .ip2(n10933), .ip3(n10932), .ip4(
        n10955), .op(n5129) );
  not_ab_or_c_or_d U12752 ( .ip1(n10935), .ip2(n7964), .ip3(n10936), .ip4(
        n10955), .op(n5128) );
  inv_1 U12753 ( .ip(n10936), .op(n10939) );
  inv_1 U12754 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[7]), .op(n10938)
         );
  inv_1 U12755 ( .ip(n10940), .op(n10937) );
  not_ab_or_c_or_d U12756 ( .ip1(n10939), .ip2(n10938), .ip3(n10937), .ip4(
        n10955), .op(n5127) );
  not_ab_or_c_or_d U12757 ( .ip1(n10940), .ip2(n7981), .ip3(n10941), .ip4(
        n10955), .op(n5126) );
  inv_1 U12758 ( .ip(n10941), .op(n10944) );
  inv_1 U12759 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[9]), .op(n10943)
         );
  inv_1 U12760 ( .ip(n10945), .op(n10942) );
  not_ab_or_c_or_d U12761 ( .ip1(n10944), .ip2(n10943), .ip3(n10942), .ip4(
        n10955), .op(n5125) );
  not_ab_or_c_or_d U12762 ( .ip1(n10945), .ip2(n7990), .ip3(n10946), .ip4(
        n10955), .op(n5124) );
  inv_1 U12763 ( .ip(n10946), .op(n10949) );
  inv_1 U12764 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[11]), .op(n10948)
         );
  inv_1 U12765 ( .ip(n10950), .op(n10947) );
  not_ab_or_c_or_d U12766 ( .ip1(n10949), .ip2(n10948), .ip3(n10947), .ip4(
        n10955), .op(n5123) );
  not_ab_or_c_or_d U12767 ( .ip1(n10950), .ip2(n7976), .ip3(n10951), .ip4(
        n10955), .op(n5122) );
  inv_1 U12768 ( .ip(n10951), .op(n10954) );
  inv_1 U12769 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[13]), .op(n10953)
         );
  inv_1 U12770 ( .ip(n10957), .op(n10952) );
  not_ab_or_c_or_d U12771 ( .ip1(n10954), .ip2(n10953), .ip3(n10952), .ip4(
        n10955), .op(n5121) );
  not_ab_or_c_or_d U12772 ( .ip1(n10957), .ip2(n7935), .ip3(n10956), .ip4(
        n10955), .op(n5120) );
  and2_1 U12773 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[0]), .ip2(
        n10958), .op(n10961) );
  not_ab_or_c_or_d U12774 ( .ip1(n10960), .ip2(n10959), .ip3(n10961), .ip4(
        n10994), .op(n5153) );
  inv_1 U12775 ( .ip(n10961), .op(n10963) );
  nand2_1 U12776 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[1]), .ip2(
        n10961), .op(n10967) );
  inv_1 U12777 ( .ip(n10967), .op(n10962) );
  not_ab_or_c_or_d U12778 ( .ip1(n10964), .ip2(n10963), .ip3(n10962), .ip4(
        n10994), .op(n5152) );
  inv_1 U12779 ( .ip(n10965), .op(n10966) );
  not_ab_or_c_or_d U12780 ( .ip1(n10968), .ip2(n10967), .ip3(n10966), .ip4(
        n10994), .op(n5151) );
  inv_1 U12781 ( .ip(n10969), .op(n10972) );
  inv_1 U12782 ( .ip(n10974), .op(n10970) );
  not_ab_or_c_or_d U12783 ( .ip1(n10972), .ip2(n10971), .ip3(n10970), .ip4(
        n10994), .op(n5149) );
  not_ab_or_c_or_d U12784 ( .ip1(n10974), .ip2(n10973), .ip3(n10975), .ip4(
        n10994), .op(n5148) );
  inv_1 U12785 ( .ip(n10975), .op(n10978) );
  inv_1 U12786 ( .ip(n10980), .op(n10976) );
  not_ab_or_c_or_d U12787 ( .ip1(n10978), .ip2(n10977), .ip3(n10976), .ip4(
        n10994), .op(n5147) );
  not_ab_or_c_or_d U12788 ( .ip1(n10980), .ip2(n10979), .ip3(n10981), .ip4(
        n10994), .op(n5146) );
  inv_1 U12789 ( .ip(n10981), .op(n10982) );
  not_ab_or_c_or_d U12790 ( .ip1(n10982), .ip2(n9021), .ip3(n10994), .ip4(
        n10986), .op(n5145) );
  not_ab_or_c_or_d U12791 ( .ip1(n10984), .ip2(n9012), .ip3(n10983), .ip4(
        n10994), .op(n5144) );
  inv_1 U12792 ( .ip(n10983), .op(n10988) );
  inv_1 U12793 ( .ip(n10989), .op(n10987) );
  not_ab_or_c_or_d U12794 ( .ip1(n10988), .ip2(n9010), .ip3(n10987), .ip4(
        n10994), .op(n5143) );
  not_ab_or_c_or_d U12795 ( .ip1(n10989), .ip2(n9029), .ip3(n10990), .ip4(
        n10994), .op(n5142) );
  inv_1 U12796 ( .ip(n10990), .op(n10992) );
  not_ab_or_c_or_d U12797 ( .ip1(n10992), .ip2(n10991), .ip3(n10993), .ip4(
        n10994), .op(n5141) );
  inv_1 U12798 ( .ip(n10993), .op(n10996) );
  not_ab_or_c_or_d U12799 ( .ip1(n10996), .ip2(n8968), .ip3(n10995), .ip4(
        n10994), .op(n5140) );
  inv_1 U12800 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[0]), .op(n10998) );
  and2_1 U12801 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[0]), .ip2(
        n10997), .op(n11000) );
  not_ab_or_c_or_d U12802 ( .ip1(n10999), .ip2(n10998), .ip3(n11041), .ip4(
        n11000), .op(n5169) );
  inv_1 U12803 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[1]), .op(n11003) );
  inv_1 U12804 ( .ip(n11000), .op(n11002) );
  nand2_1 U12805 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[1]), .ip2(
        n11000), .op(n11004) );
  inv_1 U12806 ( .ip(n11004), .op(n11001) );
  not_ab_or_c_or_d U12807 ( .ip1(n11003), .ip2(n11002), .ip3(n11041), .ip4(
        n11001), .op(n5168) );
  inv_1 U12808 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[2]), .op(n11005) );
  not_ab_or_c_or_d U12809 ( .ip1(n11005), .ip2(n11004), .ip3(n11041), .ip4(
        n11006), .op(n5167) );
  inv_1 U12810 ( .ip(n11006), .op(n11009) );
  inv_1 U12811 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[3]), .op(n11008) );
  inv_1 U12812 ( .ip(n11011), .op(n11007) );
  not_ab_or_c_or_d U12813 ( .ip1(n11009), .ip2(n11008), .ip3(n11041), .ip4(
        n11007), .op(n5166) );
  not_ab_or_c_or_d U12814 ( .ip1(n11011), .ip2(n11010), .ip3(n11041), .ip4(
        n11012), .op(n5165) );
  inv_1 U12815 ( .ip(n11012), .op(n11015) );
  inv_1 U12816 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[5]), .op(n11014) );
  inv_1 U12817 ( .ip(n11017), .op(n11013) );
  not_ab_or_c_or_d U12818 ( .ip1(n11015), .ip2(n11014), .ip3(n11041), .ip4(
        n11013), .op(n5164) );
  not_ab_or_c_or_d U12819 ( .ip1(n11017), .ip2(n11016), .ip3(n11041), .ip4(
        n11018), .op(n5163) );
  inv_1 U12820 ( .ip(n11018), .op(n11021) );
  inv_1 U12821 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[7]), .op(n11020) );
  inv_1 U12822 ( .ip(n11023), .op(n11019) );
  not_ab_or_c_or_d U12823 ( .ip1(n11021), .ip2(n11020), .ip3(n11041), .ip4(
        n11019), .op(n5162) );
  not_ab_or_c_or_d U12824 ( .ip1(n11023), .ip2(n11022), .ip3(n11041), .ip4(
        n11024), .op(n5161) );
  inv_1 U12825 ( .ip(n11024), .op(n11027) );
  inv_1 U12826 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[9]), .op(n11026) );
  inv_1 U12827 ( .ip(n11029), .op(n11025) );
  not_ab_or_c_or_d U12828 ( .ip1(n11027), .ip2(n11026), .ip3(n11041), .ip4(
        n11025), .op(n5160) );
  not_ab_or_c_or_d U12829 ( .ip1(n11029), .ip2(n11028), .ip3(n11041), .ip4(
        n11030), .op(n5159) );
  inv_1 U12830 ( .ip(n11030), .op(n11033) );
  inv_1 U12831 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[11]), .op(
        n11032) );
  inv_1 U12832 ( .ip(n11035), .op(n11031) );
  not_ab_or_c_or_d U12833 ( .ip1(n11033), .ip2(n11032), .ip3(n11041), .ip4(
        n11031), .op(n5158) );
  not_ab_or_c_or_d U12834 ( .ip1(n11035), .ip2(n11034), .ip3(n11041), .ip4(
        n11036), .op(n5157) );
  inv_1 U12835 ( .ip(n11036), .op(n11039) );
  inv_1 U12836 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[13]), .op(
        n11038) );
  inv_1 U12837 ( .ip(n11043), .op(n11037) );
  not_ab_or_c_or_d U12838 ( .ip1(n11039), .ip2(n11038), .ip3(n11041), .ip4(
        n11037), .op(n5156) );
  not_ab_or_c_or_d U12839 ( .ip1(n11043), .ip2(n11042), .ip3(n11041), .ip4(
        n11040), .op(n5155) );
  inv_1 U12840 ( .ip(n11044), .op(n11046) );
  and4_1 U12841 ( .ip1(n11305), .ip2(n11047), .ip3(n11046), .ip4(n11045), .op(
        n11055) );
  nor2_1 U12842 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(n11048), .op(n11049) );
  nor3_1 U12843 ( .ip1(n11051), .ip2(n11050), .ip3(n11049), .op(n11054) );
  nor2_1 U12844 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_byte_waiting_q), .ip2(n11055), 
        .op(n11052) );
  not_ab_or_c_or_d U12845 ( .ip1(n11055), .ip2(n11054), .ip3(n11053), .ip4(
        n11052), .op(n5191) );
  not_ab_or_c_or_d U12846 ( .ip1(n11058), .ip2(n11057), .ip3(n11059), .ip4(
        n11099), .op(n4956) );
  inv_1 U12847 ( .ip(n11059), .op(n11061) );
  nand2_1 U12848 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[2]), 
        .ip2(n11059), .op(n11066) );
  inv_1 U12849 ( .ip(n11066), .op(n11060) );
  not_ab_or_c_or_d U12850 ( .ip1(n11062), .ip2(n11061), .ip3(n11060), .ip4(
        n11099), .op(n4955) );
  inv_1 U12851 ( .ip(n11063), .op(n11064) );
  nor2_1 U12852 ( .ip1(n11065), .ip2(n11064), .op(n11068) );
  not_ab_or_c_or_d U12853 ( .ip1(n11067), .ip2(n11066), .ip3(n11068), .ip4(
        n11099), .op(n4954) );
  inv_1 U12854 ( .ip(n11068), .op(n11069) );
  and2_1 U12855 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[4]), .ip2(
        n11068), .op(n11071) );
  not_ab_or_c_or_d U12856 ( .ip1(n11070), .ip2(n11069), .ip3(n11071), .ip4(
        n11099), .op(n4953) );
  inv_1 U12857 ( .ip(n11071), .op(n11073) );
  nand2_1 U12858 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[5]), 
        .ip2(n11071), .op(n11075) );
  inv_1 U12859 ( .ip(n11075), .op(n11072) );
  not_ab_or_c_or_d U12860 ( .ip1(n11074), .ip2(n11073), .ip3(n11072), .ip4(
        n11099), .op(n4952) );
  not_ab_or_c_or_d U12861 ( .ip1(n11076), .ip2(n11075), .ip3(n11077), .ip4(
        n11099), .op(n4951) );
  inv_1 U12862 ( .ip(n11077), .op(n11079) );
  inv_1 U12863 ( .ip(n11081), .op(n11078) );
  not_ab_or_c_or_d U12864 ( .ip1(n11080), .ip2(n11079), .ip3(n11078), .ip4(
        n11099), .op(n4950) );
  not_ab_or_c_or_d U12865 ( .ip1(n11082), .ip2(n11081), .ip3(n11083), .ip4(
        n11099), .op(n4949) );
  inv_1 U12866 ( .ip(n11083), .op(n11085) );
  not_ab_or_c_or_d U12867 ( .ip1(n11086), .ip2(n11085), .ip3(n11084), .ip4(
        n11099), .op(n4948) );
  or2_1 U12868 ( .ip1(n11089), .ip2(n11088), .op(n11091) );
  inv_1 U12869 ( .ip(n11091), .op(n11087) );
  not_ab_or_c_or_d U12870 ( .ip1(n11089), .ip2(n11088), .ip3(n11087), .ip4(
        n11099), .op(n4947) );
  inv_1 U12871 ( .ip(n11093), .op(n11090) );
  not_ab_or_c_or_d U12872 ( .ip1(n11092), .ip2(n11091), .ip3(n11099), .ip4(
        n11090), .op(n4946) );
  nor2_2 U12873 ( .ip1(n11094), .ip2(n11093), .op(n11095) );
  not_ab_or_c_or_d U12874 ( .ip1(n11094), .ip2(n11093), .ip3(n11095), .ip4(
        n11099), .op(n4945) );
  inv_1 U12875 ( .ip(n11095), .op(n11097) );
  nand2_1 U12876 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[13]), 
        .ip2(n11095), .op(n11101) );
  inv_1 U12877 ( .ip(n11101), .op(n11096) );
  not_ab_or_c_or_d U12878 ( .ip1(n11098), .ip2(n11097), .ip3(n11099), .ip4(
        n11096), .op(n4944) );
  nor2_1 U12879 ( .ip1(n11102), .ip2(n11101), .op(n11100) );
  not_ab_or_c_or_d U12880 ( .ip1(n11102), .ip2(n11101), .ip3(n11100), .ip4(
        n11099), .op(n4943) );
  nand3_1 U12881 ( .ip1(n11104), .ip2(i_i2c_U_DW_apb_i2c_tx_shift_N281), .ip3(
        n11103), .op(n11107) );
  and2_1 U12882 ( .ip1(n11106), .ip2(n11105), .op(n11108) );
  nor2_1 U12883 ( .ip1(n11107), .ip2(n11108), .op(n11112) );
  inv_1 U12884 ( .ip(n11108), .op(n11109) );
  nor2_1 U12885 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_ic_data_oe_early), .ip2(
        n11109), .op(n11111) );
  not_ab_or_c_or_d U12886 ( .ip1(n4941), .ip2(n11112), .ip3(n11111), .ip4(
        n11110), .op(i_i2c_U_DW_apb_i2c_tx_shift_N85) );
  not_ab_or_c_or_d U12887 ( .ip1(n11115), .ip2(n11114), .ip3(n11721), .ip4(
        n11113), .op(n5087) );
  nor2_1 U12888 ( .ip1(i_i2c_mst_rx_bit_count[3]), .ip2(n11116), .op(n11120)
         );
  nor3_1 U12889 ( .ip1(i_i2c_mst_rx_bit_count[3]), .ip2(n11116), .ip3(n11167), 
        .op(n11117) );
  nor2_1 U12890 ( .ip1(i_i2c_rx_current_src_en), .ip2(n11117), .op(n11118) );
  not_ab_or_c_or_d U12891 ( .ip1(n11120), .ip2(n11119), .ip3(n11118), .ip4(
        n11170), .op(n5070) );
  nand2_1 U12892 ( .ip1(i_ssi_rx_rd_addr[0]), .ip2(n11164), .op(n11127) );
  inv_1 U12893 ( .ip(n11127), .op(n11122) );
  nand2_1 U12894 ( .ip1(i_ssi_U_fifo_U_rx_fifo_rd_addr_at_max), .ip2(n11164), 
        .op(n11121) );
  nand2_1 U12895 ( .ip1(n11219), .ip2(n11121), .op(n11128) );
  not_ab_or_c_or_d U12896 ( .ip1(n11124), .ip2(n11123), .ip3(n11122), .ip4(
        n11128), .op(n11768) );
  nor2_1 U12897 ( .ip1(n11125), .ip2(n11124), .op(n11130) );
  not_ab_or_c_or_d U12898 ( .ip1(n11127), .ip2(n11126), .ip3(n11130), .ip4(
        n11128), .op(i_ssi_U_fifo_U_rx_fifo_N45) );
  nor2_1 U12899 ( .ip1(i_ssi_rx_rd_addr[2]), .ip2(n11130), .op(n11129) );
  not_ab_or_c_or_d U12900 ( .ip1(n11130), .ip2(i_ssi_rx_rd_addr[2]), .ip3(
        n11129), .ip4(n11128), .op(i_ssi_U_fifo_U_rx_fifo_N46) );
  inv_1 U12901 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[1]), .op(
        n11132) );
  inv_1 U12902 ( .ip(n11140), .op(n11131) );
  not_ab_or_c_or_d U12903 ( .ip1(n11133), .ip2(n11132), .ip3(n11144), .ip4(
        n11131), .op(n5102) );
  inv_1 U12904 ( .ip(n11138), .op(n11136) );
  inv_1 U12905 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[3]), .op(
        n11135) );
  inv_1 U12906 ( .ip(n11143), .op(n11134) );
  not_ab_or_c_or_d U12907 ( .ip1(n11136), .ip2(n11135), .ip3(n11144), .ip4(
        n11134), .op(n5100) );
  nor2_1 U12908 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[6]), 
        .ip2(n11145), .op(n11137) );
  not_ab_or_c_or_d U12909 ( .ip1(n11145), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[6]), .ip3(n11137), 
        .ip4(n11144), .op(n5097) );
  not_ab_or_c_or_d U12910 ( .ip1(n11140), .ip2(n11139), .ip3(n11138), .ip4(
        n11144), .op(n5101) );
  not_ab_or_c_or_d U12911 ( .ip1(n11143), .ip2(n11142), .ip3(n11141), .ip4(
        n11144), .op(n5099) );
  not_ab_or_c_or_d U12912 ( .ip1(n11147), .ip2(n11146), .ip3(n11145), .ip4(
        n11144), .op(n5098) );
  inv_1 U12913 ( .ip(i_ssi_rxftlr[0]), .op(n11234) );
  nor3_1 U12914 ( .ip1(n11234), .ip2(n11228), .ip3(n11229), .op(n11150) );
  nor2_1 U12915 ( .ip1(i_ssi_U_fifo_switch_almost_full), .ip2(n11150), .op(
        n11149) );
  not_ab_or_c_or_d U12916 ( .ip1(n11151), .ip2(n11150), .ip3(n11149), .ip4(
        n11148), .op(i_ssi_U_intctl_N33) );
  nor2_1 U12917 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[3]), .ip2(
        n11152), .op(n11153) );
  nor2_1 U12918 ( .ip1(n11154), .ip2(n11153), .op(n11155) );
  nor2_1 U12919 ( .ip1(n11156), .ip2(n11155), .op(n11163) );
  nand2_1 U12920 ( .ip1(n11158), .ip2(n11157), .op(n11162) );
  inv_1 U12921 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_data_scl), .op(n11159) );
  nor2_1 U12922 ( .ip1(n11163), .ip2(n11159), .op(n11161) );
  ab_or_c_or_d U12923 ( .ip1(n11163), .ip2(n11162), .ip3(n11161), .ip4(n11160), 
        .op(n4124) );
  not_ab_or_c_or_d U12924 ( .ip1(n11166), .ip2(n11165), .ip3(n11227), .ip4(
        n11164), .op(i_ssi_U_fifo_U_rx_fifo_N38) );
  nor3_1 U12925 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[3]), .ip2(
        n11168), .ip3(n11167), .op(n11169) );
  nor2_1 U12926 ( .ip1(i_i2c_tx_current_src_en), .ip2(n11169), .op(n11171) );
  not_ab_or_c_or_d U12927 ( .ip1(n11173), .ip2(n11172), .ip3(n11171), .ip4(
        n11170), .op(n5069) );
  and4_1 U12929 ( .ip1(i_i2c_slv_tx_ready_unconn), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly1), .ip3(n11175), .ip4(
        n11174), .op(n11312) );
  nor2_1 U12930 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[0]), .ip2(
        n11312), .op(n11176) );
  not_ab_or_c_or_d U12931 ( .ip1(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[0]), .ip2(n11312), .ip3(
        n11176), .ip4(n11316), .op(n5108) );
  inv_1 U12932 ( .ip(i_apb_U_DW_apb_ahbsif_use_saved_c), .op(n11360) );
  nor2_1 U12933 ( .ip1(i_apb_pclk_en), .ip2(n11360), .op(
        i_apb_U_DW_apb_ahbsif_N727) );
  or2_1 U12934 ( .ip1(i_i2c_rx_current_src_en), .ip2(i_i2c_tx_current_src_en), 
        .op(i_i2c_U_DW_apb_i2c_toggle_N29) );
  and2_1 U12935 ( .ip1(i_i2c_ic_raw_intr_stat[0]), .ip2(i_i2c_ic_intr_mask[0]), 
        .op(i_i2c_ic_intr_stat[0]) );
  and2_1 U12936 ( .ip1(i_i2c_ic_raw_intr_stat[1]), .ip2(i_i2c_ic_intr_mask[1]), 
        .op(i_i2c_ic_intr_stat[1]) );
  inv_1 U12937 ( .ip(n11177), .op(n11181) );
  nor2_1 U12938 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_i_rx_almost_full), .ip2(n11181), 
        .op(n11179) );
  not_ab_or_c_or_d U12939 ( .ip1(n11181), .ip2(n11180), .ip3(n11179), .ip4(
        n11178), .op(i_i2c_ic_raw_intr_stat[2]) );
  and2_1 U12940 ( .ip1(i_i2c_ic_raw_intr_stat[2]), .ip2(i_i2c_ic_intr_mask[2]), 
        .op(i_i2c_ic_intr_stat[2]) );
  and2_1 U12941 ( .ip1(i_i2c_ic_raw_intr_stat[3]), .ip2(i_i2c_ic_intr_mask[3]), 
        .op(i_i2c_ic_intr_stat[3]) );
  and2_1 U12942 ( .ip1(i_i2c_ic_raw_intr_stat[4]), .ip2(i_i2c_ic_intr_mask[4]), 
        .op(i_i2c_ic_intr_stat[4]) );
  and2_1 U12943 ( .ip1(i_i2c_ic_raw_intr_stat[5]), .ip2(i_i2c_ic_intr_mask[5]), 
        .op(i_i2c_ic_intr_stat[5]) );
  and2_1 U12944 ( .ip1(i_i2c_ic_raw_intr_stat[6]), .ip2(i_i2c_ic_intr_mask[6]), 
        .op(i_i2c_ic_intr_stat[6]) );
  and2_1 U12945 ( .ip1(i_i2c_ic_raw_intr_stat[7]), .ip2(i_i2c_ic_intr_mask[7]), 
        .op(i_i2c_ic_intr_stat[7]) );
  and2_1 U12946 ( .ip1(i_i2c_ic_raw_intr_stat[8]), .ip2(i_i2c_ic_intr_mask[8]), 
        .op(i_i2c_ic_intr_stat[8]) );
  and2_1 U12947 ( .ip1(i_i2c_ic_raw_intr_stat[9]), .ip2(i_i2c_ic_intr_mask[9]), 
        .op(i_i2c_ic_intr_stat[9]) );
  and2_1 U12948 ( .ip1(i_i2c_ic_raw_intr_stat[10]), .ip2(
        i_i2c_ic_intr_mask[10]), .op(i_i2c_ic_intr_stat[10]) );
  and2_1 U12949 ( .ip1(i_i2c_ic_raw_intr_stat[11]), .ip2(
        i_i2c_ic_intr_mask[11]), .op(i_i2c_ic_intr_stat[11]) );
  or2_1 U12950 ( .ip1(i_i2c_ic_enable[0]), .ip2(i_i2c_activity), .op(
        i_i2c_U_DW_apb_i2c_intctl_N4) );
  xor2_1 U12951 ( .ip1(i_i2c_U_DW_apb_i2c_intctl_slv_clr_leftover_flg_sync), 
        .ip2(i_i2c_U_DW_apb_i2c_intctl_slv_clr_leftover_flg_sync_q), .op(
        i_i2c_slv_clr_leftover_flg_edg) );
  or2_1 U12952 ( .ip1(i_i2c_re_start_en), .ip2(i_i2c_split_start_en), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_N207) );
  nor2_1 U12953 ( .ip1(n11182), .ip2(i_ahb_U_dfltslv_current_state), .op(
        i_ahb_U_dfltslv_next_state) );
  nor2_1 U12954 ( .ip1(n11205), .ip2(n11203), .op(n11202) );
  inv_1 U12955 ( .ip(n11202), .op(n11185) );
  nor2_1 U12956 ( .ip1(n11205), .ip2(n11183), .op(n11187) );
  nand2_1 U12957 ( .ip1(n11189), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_rd_addr_at_max), .op(n11184) );
  not_ab_or_c_or_d U12958 ( .ip1(n11186), .ip2(n11185), .ip3(n11187), .ip4(
        n11201), .op(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N45) );
  nor2_1 U12959 ( .ip1(i_i2c_rx_rd_addr[2]), .ip2(n11187), .op(n11188) );
  not_ab_or_c_or_d U12960 ( .ip1(n11190), .ip2(n11189), .ip3(n11188), .ip4(
        n11201), .op(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N46) );
  nand3_1 U12961 ( .ip1(n11191), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_wr_addr_at_max), .ip3(
        i_i2c_rx_push_sync), .op(n11192) );
  nor2_1 U12962 ( .ip1(n11194), .ip2(n11193), .op(n11196) );
  not_ab_or_c_or_d U12963 ( .ip1(n11194), .ip2(n11193), .ip3(n11198), .ip4(
        n11196), .op(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N42) );
  nor2_1 U12964 ( .ip1(i_i2c_rx_wr_addr[2]), .ip2(n11196), .op(n11195) );
  not_ab_or_c_or_d U12965 ( .ip1(i_i2c_rx_wr_addr[2]), .ip2(n11196), .ip3(
        n11198), .ip4(n11195), .op(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N43) );
  inv_1 U12966 ( .ip(n11197), .op(n11200) );
  nor2_1 U12967 ( .ip1(i_i2c_rx_wr_addr[0]), .ip2(n11200), .op(n11199) );
  not_ab_or_c_or_d U12968 ( .ip1(i_i2c_rx_wr_addr[0]), .ip2(n11200), .ip3(
        n11199), .ip4(n11198), .op(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N41) );
  and3_1 U12969 ( .ip1(i_i2c_rx_wr_addr[1]), .ip2(i_i2c_rx_wr_addr[2]), .ip3(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N41), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N40) );
  not_ab_or_c_or_d U12970 ( .ip1(n11205), .ip2(n11203), .ip3(n11202), .ip4(
        n11201), .op(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N44) );
  and3_1 U12971 ( .ip1(i_i2c_rx_rd_addr[2]), .ip2(i_i2c_rx_rd_addr[1]), .ip3(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N44), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N39) );
  inv_1 U12972 ( .ip(i_i2c_rx_push_sync), .op(n11208) );
  nand2_1 U12973 ( .ip1(n11205), .ip2(n11204), .op(n11206) );
  not_ab_or_c_or_d U12974 ( .ip1(n11209), .ip2(n11208), .ip3(n11207), .ip4(
        n11206), .op(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N38) );
  nand2_1 U12975 ( .ip1(n11217), .ip2(i_ssi_U_fifo_U_tx_fifo_wr_addr_at_max), 
        .op(n11210) );
  nand2_1 U12976 ( .ip1(n11210), .ip2(n11219), .op(n11215) );
  not_ab_or_c_or_d U12977 ( .ip1(n11212), .ip2(n11211), .ip3(n11214), .ip4(
        n11215), .op(i_ssi_U_fifo_U_tx_fifo_N42) );
  nor2_1 U12978 ( .ip1(i_ssi_tx_wr_addr[2]), .ip2(n11214), .op(n11213) );
  not_ab_or_c_or_d U12979 ( .ip1(i_ssi_tx_wr_addr[2]), .ip2(n11214), .ip3(
        n11213), .ip4(n11215), .op(i_ssi_U_fifo_U_tx_fifo_N43) );
  nor2_1 U12980 ( .ip1(n11217), .ip2(i_ssi_tx_wr_addr[0]), .op(n11216) );
  not_ab_or_c_or_d U12981 ( .ip1(n11217), .ip2(i_ssi_tx_wr_addr[0]), .ip3(
        n11216), .ip4(n11215), .op(i_ssi_U_fifo_U_tx_fifo_N41) );
  and3_1 U12982 ( .ip1(i_ssi_tx_wr_addr[2]), .ip2(i_ssi_tx_wr_addr[1]), .ip3(
        i_ssi_U_fifo_U_tx_fifo_N41), .op(i_ssi_U_fifo_U_tx_fifo_N40) );
  nand2_1 U12983 ( .ip1(n11226), .ip2(i_ssi_U_fifo_U_rx_fifo_wr_addr_at_max), 
        .op(n11218) );
  nand2_1 U12984 ( .ip1(n11219), .ip2(n11218), .op(n11224) );
  not_ab_or_c_or_d U12985 ( .ip1(n11222), .ip2(n11221), .ip3(n11220), .ip4(
        n11224), .op(i_ssi_U_fifo_U_rx_fifo_N42) );
  not_ab_or_c_or_d U12986 ( .ip1(n5323), .ip2(n11223), .ip3(n5275), .ip4(
        n11224), .op(i_ssi_U_fifo_U_rx_fifo_N43) );
  nor2_1 U12987 ( .ip1(i_ssi_rx_wr_addr[0]), .ip2(n11226), .op(n11225) );
  not_ab_or_c_or_d U12988 ( .ip1(i_ssi_rx_wr_addr[0]), .ip2(n11226), .ip3(
        n11225), .ip4(n11224), .op(i_ssi_U_fifo_U_rx_fifo_N41) );
  and3_1 U12989 ( .ip1(i_ssi_rx_wr_addr[2]), .ip2(i_ssi_rx_wr_addr[1]), .ip3(
        i_ssi_U_fifo_U_rx_fifo_N41), .op(i_ssi_U_fifo_U_rx_fifo_N40) );
  and3_1 U12990 ( .ip1(i_ssi_rx_rd_addr[2]), .ip2(i_ssi_rx_rd_addr[1]), .ip3(
        n11768), .op(i_ssi_U_fifo_U_rx_fifo_N39) );
  not_ab_or_c_or_d U12991 ( .ip1(i_ssi_rxftlr[0]), .ip2(i_ssi_rxftlr[1]), 
        .ip3(i_ssi_rxftlr[2]), .ip4(n11227), .op(n11245) );
  or2_1 U12992 ( .ip1(i_ssi_rxftlr[0]), .ip2(n11228), .op(n11231) );
  or2_1 U12993 ( .ip1(n11229), .ip2(n11228), .op(n11230) );
  nand2_1 U12994 ( .ip1(n11231), .ip2(n11230), .op(n11239) );
  nand2_4 U12995 ( .ip1(n11233), .ip2(n11232), .op(n11242) );
  or2_1 U12996 ( .ip1(n11234), .ip2(i_ssi_rxftlr[1]), .op(n11238) );
  or2_1 U12997 ( .ip1(n11236), .ip2(i_ssi_rxftlr[1]), .op(n11237) );
  not_ab_or_c_or_d U12998 ( .ip1(n11244), .ip2(n11245), .ip3(n11777), .ip4(
        n11243), .op(n11247) );
  nor3_1 U12999 ( .ip1(n11245), .ip2(i_ssi_U_fifo_U_rx_fifo_N49), .ip3(n11777), 
        .op(n11246) );
  nor2_1 U13000 ( .ip1(n11247), .ip2(n11246), .op(i_ssi_U_fifo_U_rx_fifo_N36)
         );
  or4_1 U13001 ( .ip1(i_ssi_U_fifo_U_rx_fifo_N49), .ip2(n11777), .ip3(
        i_ssi_U_fifo_U_rx_fifo_N48), .ip4(i_ssi_U_fifo_U_rx_fifo_N47), .op(
        i_ssi_U_fifo_U_rx_fifo_N33) );
  and2_1 U13002 ( .ip1(n5109), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly2), .op(
        i_i2c_U_DW_apb_i2c_tx_shift_N402) );
  nor2_1 U13003 ( .ip1(i_i2c_tx_rd_addr[2]), .ip2(n11250), .op(n11248) );
  not_ab_or_c_or_d U13004 ( .ip1(i_i2c_tx_rd_addr[2]), .ip2(n11250), .ip3(
        n11249), .ip4(n11248), .op(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N46) );
  not_ab_or_c_or_d U13005 ( .ip1(n11253), .ip2(n11252), .ip3(n11251), .ip4(
        n11254), .op(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N42) );
  not_ab_or_c_or_d U13006 ( .ip1(n11257), .ip2(n11256), .ip3(n11255), .ip4(
        n11254), .op(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N43) );
  not_ab_or_c_or_d U13007 ( .ip1(n11261), .ip2(n11260), .ip3(n11259), .ip4(
        n11258), .op(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N38) );
  inv_1 U13008 ( .ip(i_i2c_ic_10bit_mst), .op(
        i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_mst_1_sync_N2) );
  inv_1 U13009 ( .ip(i_i2c_ic_rstrt_en), .op(
        i_i2c_U_DW_apb_i2c_sync_U_ic_rstrt_en_1_sync_N2) );
  inv_1 U13010 ( .ip(i_i2c_ic_data_in_a), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_U_SYNC_N2) );
  nor2_1 U13011 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[0]), 
        .ip2(n11277), .op(i_i2c_U_DW_apb_i2c_rx_filter_N123) );
  nand2_1 U13012 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[0]), 
        .ip2(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[1]), .op(n11265)
         );
  inv_1 U13013 ( .ip(n11265), .op(n11267) );
  not_ab_or_c_or_d U13014 ( .ip1(n11263), .ip2(n11262), .ip3(n11267), .ip4(
        n11277), .op(i_i2c_U_DW_apb_i2c_rx_filter_N124) );
  not_ab_or_c_or_d U13015 ( .ip1(n11266), .ip2(n11265), .ip3(n11264), .ip4(
        n11277), .op(i_i2c_U_DW_apb_i2c_rx_filter_N125) );
  nand3_1 U13016 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[3]), 
        .ip2(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[2]), .ip3(n11267), 
        .op(n11271) );
  inv_1 U13017 ( .ip(n11271), .op(n11273) );
  not_ab_or_c_or_d U13018 ( .ip1(n11269), .ip2(n11268), .ip3(n11273), .ip4(
        n11277), .op(i_i2c_U_DW_apb_i2c_rx_filter_N126) );
  inv_1 U13019 ( .ip(n11275), .op(n11270) );
  not_ab_or_c_or_d U13020 ( .ip1(n11272), .ip2(n11271), .ip3(n11270), .ip4(
        n11277), .op(i_i2c_U_DW_apb_i2c_rx_filter_N127) );
  nand3_1 U13021 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[5]), 
        .ip2(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[4]), .ip3(n11273), 
        .op(n11279) );
  inv_1 U13022 ( .ip(n11279), .op(n11274) );
  not_ab_or_c_or_d U13023 ( .ip1(n11276), .ip2(n11275), .ip3(n11274), .ip4(
        n11277), .op(i_i2c_U_DW_apb_i2c_rx_filter_N128) );
  not_ab_or_c_or_d U13024 ( .ip1(n11280), .ip2(n11279), .ip3(n11278), .ip4(
        n11277), .op(i_i2c_U_DW_apb_i2c_rx_filter_N129) );
  inv_1 U13025 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt[1]), .op(n11281) );
  nor2_1 U13026 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt[0]), .ip2(n11281), 
        .op(n5234) );
  not_ab_or_c_or_d U13027 ( .ip1(i_i2c_tx_fifo_data_buf[8]), .ip2(n11284), 
        .ip3(n11283), .ip4(n11282), .op(n11285) );
  xor2_1 U13028 ( .ip1(i_i2c_tx_abrt_source[14]), .ip2(n11285), .op(n5220) );
  nor4_1 U13029 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[2]), .ip2(
        n11287), .ip3(n11293), .ip4(n11286), .op(n11288) );
  ab_or_c_or_d U13030 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[2]), 
        .ip2(n11289), .ip3(n11299), .ip4(n11288), .op(n5216) );
  nor2_1 U13031 ( .ip1(n11290), .ip2(n11293), .op(n11291) );
  or2_1 U13032 ( .ip1(n11292), .ip2(n11291), .op(n11300) );
  nor3_1 U13033 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[6]), .ip2(
        n11297), .ip3(n11293), .op(n11294) );
  ab_or_c_or_d U13034 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[6]), 
        .ip2(n11300), .ip3(n11299), .ip4(n11294), .op(n5212) );
  nor3_1 U13035 ( .ip1(n11297), .ip2(n11296), .ip3(n11295), .op(n11298) );
  ab_or_c_or_d U13036 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[7]), 
        .ip2(n11300), .ip3(n11299), .ip4(n11298), .op(n5211) );
  nor3_1 U13037 ( .ip1(i_i2c_slv_rx_aborted), .ip2(n11302), .ip3(n11301), .op(
        n11303) );
  nor2_1 U13038 ( .ip1(i_i2c_ic_enable_sync), .ip2(n11303), .op(n5210) );
  nor2_1 U13039 ( .ip1(i_i2c_re_start_en), .ip2(n11308), .op(n11307) );
  not_ab_or_c_or_d U13040 ( .ip1(n11308), .ip2(i_i2c_byte_wait_scl), .ip3(
        n11307), .ip4(n11306), .op(n5199) );
  ab_or_c_or_d U13041 ( .ip1(i_i2c_mst_rx_bit_count[2]), .ip2(n11311), .ip3(
        n11310), .ip4(n11309), .op(n5114) );
  inv_1 U13042 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[1]), .op(
        n11315) );
  nand2_1 U13043 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[0]), 
        .ip2(n11312), .op(n11314) );
  nand3_1 U13044 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[1]), 
        .ip2(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[0]), .ip3(n11312), 
        .op(n11318) );
  inv_1 U13045 ( .ip(n11318), .op(n11313) );
  not_ab_or_c_or_d U13046 ( .ip1(n11315), .ip2(n11314), .ip3(n11313), .ip4(
        n11316), .op(n5107) );
  not_ab_or_c_or_d U13047 ( .ip1(n11319), .ip2(n11318), .ip3(n11317), .ip4(
        n11316), .op(n5106) );
  or2_1 U13048 ( .ip1(n11320), .ip2(i_i2c_slv_fifo_filled_and_flushed), .op(
        n11322) );
  or2_1 U13049 ( .ip1(i_i2c_slv_rxbyte_rdy), .ip2(
        i_i2c_slv_fifo_filled_and_flushed), .op(n11321) );
  nand2_1 U13050 ( .ip1(n11322), .ip2(n11321), .op(n11323) );
  nor2_1 U13051 ( .ip1(i_i2c_ic_enable_sync), .ip2(n11323), .op(n5086) );
  inv_1 U13052 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[0]), 
        .op(n11324) );
  nand3_1 U13053 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[2]), 
        .ip2(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[1]), .ip3(
        n11344), .op(n11327) );
  nor2_1 U13054 ( .ip1(i_i2c_sda_int), .ip2(n11327), .op(n11325) );
  not_ab_or_c_or_d U13055 ( .ip1(n11327), .ip2(n11326), .ip3(n11721), .ip4(
        n11325), .op(n5080) );
  nor2_1 U13056 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[0]), 
        .ip2(n11328), .op(n11350) );
  nand3_1 U13057 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[2]), 
        .ip2(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[1]), .ip3(
        n11350), .op(n11331) );
  nor2_1 U13058 ( .ip1(i_i2c_sda_int), .ip2(n11331), .op(n11329) );
  not_ab_or_c_or_d U13059 ( .ip1(n11331), .ip2(n11330), .ip3(n11721), .ip4(
        n11329), .op(n5079) );
  inv_1 U13060 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[1]), 
        .op(n11348) );
  nand3_1 U13061 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[2]), 
        .ip2(n11344), .ip3(n11348), .op(n11334) );
  nor2_1 U13062 ( .ip1(i_i2c_sda_int), .ip2(n11334), .op(n11332) );
  not_ab_or_c_or_d U13063 ( .ip1(n11334), .ip2(n11333), .ip3(n11721), .ip4(
        n11332), .op(n5078) );
  nand3_1 U13064 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[2]), 
        .ip2(n11350), .ip3(n11348), .op(n11337) );
  nor2_1 U13065 ( .ip1(i_i2c_sda_int), .ip2(n11337), .op(n11335) );
  not_ab_or_c_or_d U13066 ( .ip1(n11337), .ip2(n11336), .ip3(n11721), .ip4(
        n11335), .op(n5077) );
  inv_1 U13067 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[2]), 
        .op(n11349) );
  nand3_1 U13068 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[1]), 
        .ip2(n11344), .ip3(n11349), .op(n11340) );
  nor2_1 U13069 ( .ip1(i_i2c_sda_int), .ip2(n11340), .op(n11338) );
  not_ab_or_c_or_d U13070 ( .ip1(n11340), .ip2(n11339), .ip3(n11721), .ip4(
        n11338), .op(n5076) );
  nand3_1 U13071 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[1]), 
        .ip2(n11350), .ip3(n11349), .op(n11343) );
  nor2_1 U13072 ( .ip1(i_i2c_sda_int), .ip2(n11343), .op(n11341) );
  not_ab_or_c_or_d U13073 ( .ip1(n11343), .ip2(n11342), .ip3(n11721), .ip4(
        n11341), .op(n5075) );
  nor2_1 U13074 ( .ip1(i_i2c_sda_int), .ip2(n11347), .op(n11345) );
  not_ab_or_c_or_d U13075 ( .ip1(n11347), .ip2(n11346), .ip3(n11721), .ip4(
        n11345), .op(n5074) );
  nor2_1 U13076 ( .ip1(i_i2c_sda_int), .ip2(n11353), .op(n11351) );
  not_ab_or_c_or_d U13077 ( .ip1(n11353), .ip2(n11352), .ip3(n11721), .ip4(
        n11351), .op(n5073) );
  xor2_1 U13078 ( .ip1(i_i2c_tx_abrt_source[13]), .ip2(n11354), .op(n5039) );
  nor2_1 U13079 ( .ip1(n11356), .ip2(n11355), .op(n11357) );
  or2_1 U13080 ( .ip1(n11358), .ip2(n11357), .op(n4857) );
  or2_1 U13081 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[17]), .ip2(n11359), 
        .op(n4841) );
  or2_1 U13082 ( .ip1(n11361), .ip2(n11360), .op(n11362) );
  nand2_1 U13083 ( .ip1(n11363), .ip2(n11362), .op(n11364) );
  or2_1 U13084 ( .ip1(n11365), .ip2(n11364), .op(n4826) );
  nand2_1 U13085 ( .ip1(i_apb_pwrite), .ip2(n11473), .op(n11366) );
  nand2_1 U13086 ( .ip1(n11427), .ip2(n11366), .op(n4825) );
  nand2_1 U13087 ( .ip1(n11427), .ip2(i_apb_pwdata_int[0]), .op(n11373) );
  inv_1 U13088 ( .ip(n11369), .op(n11368) );
  nand2_1 U13089 ( .ip1(n11367), .ip2(i_apb_U_DW_apb_ahbsif_use_saved_data), 
        .op(n11370) );
  nand2_1 U13090 ( .ip1(n5271), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[0]), .op(n11372) );
  nand2_1 U13091 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[0]), 
        .op(n11371) );
  nand3_1 U13092 ( .ip1(n11373), .ip2(n11372), .ip3(n11371), .op(n4791) );
  nand2_1 U13093 ( .ip1(n11427), .ip2(i_apb_pwdata_int[1]), .op(n11376) );
  nand2_1 U13094 ( .ip1(n5271), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[1]), .op(n11375) );
  nand2_1 U13095 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[1]), 
        .op(n11374) );
  nand3_1 U13096 ( .ip1(n11376), .ip2(n11375), .ip3(n11374), .op(n4790) );
  nand2_1 U13097 ( .ip1(n11427), .ip2(i_apb_pwdata_int[2]), .op(n11379) );
  nand2_1 U13098 ( .ip1(n5271), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[2]), .op(n11378) );
  nand2_1 U13099 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[2]), 
        .op(n11377) );
  nand3_1 U13100 ( .ip1(n11379), .ip2(n11378), .ip3(n11377), .op(n4789) );
  nand2_1 U13101 ( .ip1(n11427), .ip2(i_apb_pwdata_int[3]), .op(n11382) );
  nand2_1 U13102 ( .ip1(n5271), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[3]), .op(n11381) );
  nand2_1 U13103 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[3]), 
        .op(n11380) );
  nand3_1 U13104 ( .ip1(n11382), .ip2(n11381), .ip3(n11380), .op(n4788) );
  nand2_1 U13105 ( .ip1(n11427), .ip2(i_apb_pwdata_int[4]), .op(n11385) );
  nand2_1 U13106 ( .ip1(n5271), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[4]), .op(n11384) );
  nand2_1 U13107 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[4]), 
        .op(n11383) );
  nand3_1 U13108 ( .ip1(n11385), .ip2(n11384), .ip3(n11383), .op(n4787) );
  nand2_1 U13109 ( .ip1(n11427), .ip2(i_apb_pwdata_int[5]), .op(n11388) );
  nand2_1 U13110 ( .ip1(n5271), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[5]), .op(n11387) );
  nand2_1 U13111 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[5]), 
        .op(n11386) );
  nand3_1 U13112 ( .ip1(n11388), .ip2(n11387), .ip3(n11386), .op(n4786) );
  nand2_1 U13113 ( .ip1(n11427), .ip2(i_apb_pwdata_int[6]), .op(n11391) );
  nand2_1 U13114 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[6]), 
        .op(n11390) );
  nand2_1 U13115 ( .ip1(n5271), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[6]), .op(n11389) );
  nand3_1 U13116 ( .ip1(n11391), .ip2(n11390), .ip3(n11389), .op(n4785) );
  nand2_1 U13117 ( .ip1(n11427), .ip2(i_apb_pwdata_int[7]), .op(n11394) );
  nand2_1 U13118 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[7]), 
        .op(n11393) );
  nand2_1 U13119 ( .ip1(n5271), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[7]), .op(n11392) );
  nand3_1 U13120 ( .ip1(n11394), .ip2(n11393), .ip3(n11392), .op(n4784) );
  nand2_1 U13121 ( .ip1(n11427), .ip2(i_apb_pwdata_int[8]), .op(n11397) );
  nand2_1 U13122 ( .ip1(n5271), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[8]), .op(n11396) );
  nand2_1 U13123 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[8]), 
        .op(n11395) );
  nand3_1 U13124 ( .ip1(n11397), .ip2(n11396), .ip3(n11395), .op(n4783) );
  nand2_1 U13125 ( .ip1(n11427), .ip2(i_apb_pwdata_int[9]), .op(n11400) );
  nand2_1 U13126 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[9]), 
        .op(n11399) );
  nand2_1 U13127 ( .ip1(n5271), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[9]), .op(n11398) );
  nand3_1 U13128 ( .ip1(n11400), .ip2(n11399), .ip3(n11398), .op(n4782) );
  nand2_1 U13129 ( .ip1(n11427), .ip2(i_apb_pwdata_int[10]), .op(n11403) );
  nand2_1 U13130 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[10]), 
        .op(n11402) );
  nand2_1 U13131 ( .ip1(n5271), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[10]), .op(n11401) );
  nand3_1 U13132 ( .ip1(n11403), .ip2(n11402), .ip3(n11401), .op(n4781) );
  nand2_1 U13133 ( .ip1(n11427), .ip2(i_apb_pwdata_int[11]), .op(n11406) );
  nand2_1 U13134 ( .ip1(n5271), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[11]), .op(n11405) );
  nand2_1 U13135 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[11]), 
        .op(n11404) );
  nand3_1 U13136 ( .ip1(n11406), .ip2(n11405), .ip3(n11404), .op(n4780) );
  nand2_1 U13137 ( .ip1(n11427), .ip2(i_apb_pwdata_int[12]), .op(n11411) );
  nand2_1 U13138 ( .ip1(n5271), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[12]), .op(n11410) );
  nand2_1 U13139 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[12]), 
        .op(n11409) );
  nand3_1 U13140 ( .ip1(n11411), .ip2(n11410), .ip3(n11409), .op(n4779) );
  nand2_1 U13141 ( .ip1(n11427), .ip2(i_apb_pwdata_int[13]), .op(n11414) );
  nand2_1 U13142 ( .ip1(n5271), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[13]), .op(n11413) );
  nand2_1 U13143 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[13]), 
        .op(n11412) );
  nand3_1 U13144 ( .ip1(n11414), .ip2(n11413), .ip3(n11412), .op(n4778) );
  nand2_1 U13145 ( .ip1(n11427), .ip2(i_apb_pwdata_int[14]), .op(n11417) );
  nand2_1 U13146 ( .ip1(n5271), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[14]), .op(n11416) );
  nand2_1 U13147 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[14]), 
        .op(n11415) );
  nand3_1 U13148 ( .ip1(n11417), .ip2(n11416), .ip3(n11415), .op(n4777) );
  nand2_1 U13149 ( .ip1(n11427), .ip2(i_apb_pwdata_int[15]), .op(n11420) );
  nand2_1 U13150 ( .ip1(n5271), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[15]), .op(n11419) );
  nand2_1 U13151 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[15]), 
        .op(n11418) );
  nand3_1 U13152 ( .ip1(n11420), .ip2(n11419), .ip3(n11418), .op(n4776) );
  nand2_1 U13153 ( .ip1(n11427), .ip2(i_apb_pwdata_int[16]), .op(n11423) );
  nand2_1 U13154 ( .ip1(n5271), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[16]), .op(n11422) );
  nand2_1 U13155 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[16]), 
        .op(n11421) );
  nand3_1 U13156 ( .ip1(n11423), .ip2(n11422), .ip3(n11421), .op(n4775) );
  nand2_1 U13157 ( .ip1(n11427), .ip2(i_apb_pwdata_int[17]), .op(n11426) );
  nand2_1 U13158 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[17]), 
        .op(n11425) );
  nand2_1 U13159 ( .ip1(n5271), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[17]), .op(n11424) );
  nand3_1 U13160 ( .ip1(n11426), .ip2(n11425), .ip3(n11424), .op(n4774) );
  nand2_1 U13161 ( .ip1(n11427), .ip2(i_apb_pwdata_int[18]), .op(n11430) );
  nand2_1 U13162 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[18]), 
        .op(n11429) );
  nand2_1 U13163 ( .ip1(n5271), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[18]), .op(n11428) );
  nand3_1 U13164 ( .ip1(n11430), .ip2(n11429), .ip3(n11428), .op(n4773) );
  nand2_1 U13165 ( .ip1(n11427), .ip2(i_apb_pwdata_int[19]), .op(n11433) );
  nand2_1 U13166 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[19]), 
        .op(n11432) );
  nand2_1 U13167 ( .ip1(n5271), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[19]), .op(n11431) );
  nand3_1 U13168 ( .ip1(n11433), .ip2(n11432), .ip3(n11431), .op(n4772) );
  nand2_1 U13169 ( .ip1(n11427), .ip2(i_apb_pwdata_int[20]), .op(n11436) );
  nand2_1 U13170 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[20]), 
        .op(n11435) );
  nand2_1 U13171 ( .ip1(n5271), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[20]), .op(n11434) );
  nand3_1 U13172 ( .ip1(n11436), .ip2(n11435), .ip3(n11434), .op(n4771) );
  nand2_1 U13173 ( .ip1(n11427), .ip2(i_apb_pwdata_int[21]), .op(n11439) );
  nand2_1 U13174 ( .ip1(n5271), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[21]), .op(n11438) );
  nand2_1 U13175 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[21]), 
        .op(n11437) );
  nand3_1 U13176 ( .ip1(n11439), .ip2(n11438), .ip3(n11437), .op(n4770) );
  nand2_1 U13177 ( .ip1(n11427), .ip2(i_apb_pwdata_int[22]), .op(n11442) );
  nand2_1 U13178 ( .ip1(n5271), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[22]), .op(n11441) );
  nand2_1 U13179 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[22]), 
        .op(n11440) );
  nand3_1 U13180 ( .ip1(n11442), .ip2(n11441), .ip3(n11440), .op(n4769) );
  nand2_1 U13181 ( .ip1(n11427), .ip2(i_apb_pwdata_int[23]), .op(n11445) );
  nand2_1 U13182 ( .ip1(n5271), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[23]), .op(n11444) );
  nand2_1 U13183 ( .ip1(n11408), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[23]), 
        .op(n11443) );
  nand3_1 U13184 ( .ip1(n11445), .ip2(n11444), .ip3(n11443), .op(n4768) );
  nand2_1 U13185 ( .ip1(n11466), .ip2(i_apb_U_DW_apb_ahbsif_piped_haddr_c[2]), 
        .op(n11448) );
  nand2_1 U13186 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[2]), .ip2(n5270), 
        .op(n11447) );
  nand2_1 U13187 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[2]), .ip2(n11465), 
        .op(n11446) );
  nand3_1 U13188 ( .ip1(n11448), .ip2(n11447), .ip3(n11446), .op(n4759) );
  nand2_1 U13189 ( .ip1(n5270), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[4]), 
        .op(n11451) );
  nand2_1 U13190 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[4]), .ip2(n11466), 
        .op(n11450) );
  nand2_1 U13191 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[4]), .ip2(n11461), 
        .op(n11449) );
  nand3_1 U13192 ( .ip1(n11451), .ip2(n11450), .ip3(n11449), .op(n4757) );
  nand2_1 U13193 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[5]), .ip2(n11466), 
        .op(n11454) );
  nand2_1 U13194 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[5]), .ip2(n11461), 
        .op(n11453) );
  nand2_1 U13195 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[5]), .ip2(n5270), 
        .op(n11452) );
  nand3_1 U13196 ( .ip1(n11454), .ip2(n11453), .ip3(n11452), .op(n4756) );
  nand2_1 U13197 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[6]), .ip2(n11461), 
        .op(n11457) );
  nand2_1 U13198 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[6]), .ip2(n11466), 
        .op(n11456) );
  nand2_1 U13199 ( .ip1(n5270), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[6]), 
        .op(n11455) );
  nand3_1 U13200 ( .ip1(n11457), .ip2(n11456), .ip3(n11455), .op(n4755) );
  nand2_1 U13201 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[7]), .ip2(n11466), 
        .op(n11460) );
  nand2_1 U13202 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[7]), .ip2(n11465), 
        .op(n11459) );
  nand2_1 U13203 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[7]), .ip2(n5270), 
        .op(n11458) );
  nand3_1 U13204 ( .ip1(n11460), .ip2(n11459), .ip3(n11458), .op(n4754) );
  nand2_1 U13205 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[12]), .ip2(n11466), 
        .op(n11464) );
  nand2_1 U13206 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[12]), .ip2(n11461), 
        .op(n11463) );
  nand2_1 U13207 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[12]), .ip2(n5270), 
        .op(n11462) );
  nand3_1 U13208 ( .ip1(n11464), .ip2(n11463), .ip3(n11462), .op(n4753) );
  nand2_1 U13209 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[17]), .ip2(n11465), 
        .op(n11469) );
  nand2_1 U13210 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[17]), .ip2(n11466), 
        .op(n11468) );
  nand2_1 U13211 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[17]), .ip2(n5270), 
        .op(n11467) );
  nand3_1 U13212 ( .ip1(n11469), .ip2(n11468), .ip3(n11467), .op(n4748) );
  or2_1 U13213 ( .ip1(n11471), .ip2(n11470), .op(n11472) );
  nand2_1 U13214 ( .ip1(n11472), .ip2(i_apb_U_DW_apb_ahbsif_pipeline_c), .op(
        n11474) );
  nor2_1 U13215 ( .ip1(n11474), .ip2(n11473), .op(n11475) );
  nand2_1 U13216 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[2]), .ip2(n11506), 
        .op(n11480) );
  nand2_1 U13217 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[2]), .ip2(n5269), 
        .op(n11479) );
  nand2_1 U13218 ( .ip1(n11507), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[2]), 
        .op(n11478) );
  nand2_1 U13219 ( .ip1(i_ssi_reg_addr[0]), .ip2(n11497), .op(n11477) );
  nand4_1 U13220 ( .ip1(n11480), .ip2(n11479), .ip3(n11478), .ip4(n11477), 
        .op(n4733) );
  nand2_1 U13221 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[3]), .ip2(n5269), 
        .op(n11484) );
  nand2_1 U13222 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[3]), .ip2(n11506), 
        .op(n11483) );
  nand2_1 U13223 ( .ip1(i_ssi_reg_addr[1]), .ip2(n11497), .op(n11482) );
  nand2_1 U13224 ( .ip1(n11507), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[3]), 
        .op(n11481) );
  nand4_1 U13225 ( .ip1(n11484), .ip2(n11483), .ip3(n11482), .ip4(n11481), 
        .op(n4732) );
  nand2_1 U13226 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[4]), .ip2(n5269), 
        .op(n11488) );
  nand2_1 U13227 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[4]), .ip2(n11506), 
        .op(n11487) );
  nand2_1 U13228 ( .ip1(i_ssi_reg_addr[2]), .ip2(n11497), .op(n11486) );
  nand2_1 U13229 ( .ip1(n11507), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[4]), 
        .op(n11485) );
  nand4_1 U13230 ( .ip1(n11488), .ip2(n11487), .ip3(n11486), .ip4(n11485), 
        .op(n4731) );
  nand2_1 U13231 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[5]), .ip2(n11506), 
        .op(n11492) );
  nand2_1 U13232 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[5]), .ip2(n5269), 
        .op(n11491) );
  nand2_1 U13233 ( .ip1(i_ssi_reg_addr[3]), .ip2(n11497), .op(n11490) );
  nand2_1 U13234 ( .ip1(n11507), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[5]), 
        .op(n11489) );
  nand4_1 U13235 ( .ip1(n11492), .ip2(n11491), .ip3(n11490), .ip4(n11489), 
        .op(n4730) );
  nand2_1 U13236 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[6]), .ip2(n5269), 
        .op(n11496) );
  nand2_1 U13237 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[6]), .ip2(n11506), 
        .op(n11495) );
  nand2_1 U13238 ( .ip1(n11507), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[6]), 
        .op(n11494) );
  nand2_1 U13239 ( .ip1(i_ssi_reg_addr[4]), .ip2(n11497), .op(n11493) );
  nand4_1 U13240 ( .ip1(n11496), .ip2(n11495), .ip3(n11494), .ip4(n11493), 
        .op(n4729) );
  nand2_1 U13241 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[7]), .ip2(n11506), 
        .op(n11501) );
  nand2_1 U13242 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[7]), .ip2(n5269), 
        .op(n11500) );
  nand2_1 U13243 ( .ip1(n11507), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[7]), 
        .op(n11499) );
  nand2_1 U13244 ( .ip1(i_ssi_reg_addr[5]), .ip2(n11497), .op(n11498) );
  nand4_1 U13245 ( .ip1(n11501), .ip2(n11500), .ip3(n11499), .ip4(n11498), 
        .op(n4728) );
  nand2_1 U13246 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[12]), .ip2(n11506), 
        .op(n11505) );
  nand2_1 U13247 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[12]), .ip2(n5269), 
        .op(n11504) );
  nand2_1 U13248 ( .ip1(i_apb_paddr[12]), .ip2(n11497), .op(n11503) );
  nand2_1 U13249 ( .ip1(n11507), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[12]), 
        .op(n11502) );
  nand4_1 U13250 ( .ip1(n11505), .ip2(n11504), .ip3(n11503), .ip4(n11502), 
        .op(n4727) );
  nand2_1 U13251 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[17]), .ip2(n11506), 
        .op(n11511) );
  nand2_1 U13252 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_haddr_c[17]), .ip2(n5269), 
        .op(n11510) );
  nand2_1 U13253 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[17]), .ip2(n11507), 
        .op(n11509) );
  nand2_1 U13254 ( .ip1(i_apb_paddr[17]), .ip2(n11497), .op(n11508) );
  nand4_1 U13255 ( .ip1(n11511), .ip2(n11510), .ip3(n11509), .ip4(n11508), 
        .op(n4722) );
  nand2_1 U13256 ( .ip1(n11513), .ip2(i_ssi_U_regfile_txflr[3]), .op(n11515)
         );
  nor2_1 U13257 ( .ip1(n11519), .ip2(n11518), .op(n11520) );
  or2_1 U13258 ( .ip1(n11521), .ip2(n11520), .op(n4455) );
  nand2_1 U13259 ( .ip1(n11522), .ip2(i_ssi_U_regfile_rxflr[3]), .op(n11523)
         );
  nand2_1 U13260 ( .ip1(n11524), .ip2(n11523), .op(n11525) );
  nand2_1 U13261 ( .ip1(i_ssi_U_regfile_rxflr[2]), .ip2(n11525), .op(n11528)
         );
  nand2_1 U13262 ( .ip1(i_ssi_U_regfile_rxflr[3]), .ip2(n11526), .op(n11527)
         );
  nand2_1 U13263 ( .ip1(n11528), .ip2(n11527), .op(n4448) );
  or2_1 U13264 ( .ip1(n11530), .ip2(n11529), .op(n11534) );
  or2_1 U13265 ( .ip1(n11532), .ip2(n11531), .op(n11533) );
  nand3_1 U13266 ( .ip1(n11535), .ip2(n11534), .ip3(n11533), .op(n4446) );
  inv_1 U13267 ( .ip(n11536), .op(n11550) );
  nand2_1 U13268 ( .ip1(n11550), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[8]), .op(n11538) );
  nand2_1 U13269 ( .ip1(n6655), .ip2(i_ssi_rx_push_data[8]), .op(n11537) );
  nand2_1 U13270 ( .ip1(n11538), .ip2(n11537), .op(n4437) );
  nand2_1 U13271 ( .ip1(n6655), .ip2(i_ssi_rx_push_data[9]), .op(n11542) );
  inv_1 U13272 ( .ip(n11555), .op(n11539) );
  nand2_1 U13273 ( .ip1(n11539), .ip2(n11547), .op(n11540) );
  nand3_1 U13274 ( .ip1(n11550), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[9]), .ip3(n11540), .op(n11541)
         );
  nand2_1 U13275 ( .ip1(n11542), .ip2(n11541), .op(n4436) );
  nand2_1 U13276 ( .ip1(n6655), .ip2(i_ssi_rx_push_data[10]), .op(n11546) );
  nand2_1 U13277 ( .ip1(n11543), .ip2(n11547), .op(n11544) );
  nand3_1 U13278 ( .ip1(n11550), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[10]), .ip3(n11544), .op(n11545) );
  nand2_1 U13279 ( .ip1(n11546), .ip2(n11545), .op(n4435) );
  nand2_1 U13280 ( .ip1(n6655), .ip2(i_ssi_rx_push_data[11]), .op(n11552) );
  inv_1 U13281 ( .ip(n11558), .op(n11548) );
  nand2_1 U13282 ( .ip1(n11548), .ip2(n11547), .op(n11549) );
  nand3_1 U13283 ( .ip1(n11550), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[11]), .ip3(n11549), .op(n11551) );
  nand2_1 U13284 ( .ip1(n11552), .ip2(n11551), .op(n4434) );
  nand2_1 U13285 ( .ip1(n11559), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[12]), .op(n11554) );
  nand2_1 U13286 ( .ip1(n6655), .ip2(i_ssi_rx_push_data[12]), .op(n11553) );
  nand2_1 U13287 ( .ip1(n11554), .ip2(n11553), .op(n4433) );
  nand3_1 U13288 ( .ip1(n11559), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[13]), .ip3(n11555), .op(n11557) );
  nand2_1 U13289 ( .ip1(n6655), .ip2(i_ssi_rx_push_data[13]), .op(n11556) );
  nand2_1 U13290 ( .ip1(n11557), .ip2(n11556), .op(n4432) );
  nand3_1 U13291 ( .ip1(n11559), .ip2(n11558), .ip3(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[15]), .op(n11561) );
  nand2_1 U13292 ( .ip1(n6655), .ip2(i_ssi_rx_push_data[15]), .op(n11560) );
  nand2_1 U13293 ( .ip1(n11561), .ip2(n11560), .op(n4430) );
  nand2_1 U13294 ( .ip1(i_ssi_dfs[0]), .ip2(n11692), .op(n11566) );
  nand2_1 U13295 ( .ip1(i_ssi_ser_0_), .ip2(n11563), .op(n11565) );
  nand2_1 U13296 ( .ip1(i_ssi_U_regfile_ctrlr1_int[0]), .ip2(n11693), .op(
        n11564) );
  nand3_1 U13297 ( .ip1(n11566), .ip2(n11565), .ip3(n11564), .op(n11570) );
  mux3_2 U13298 ( .ip1(n11570), .ip2(n5282), .ip3(n11569), .s0(n11568), .s1(
        n11567), .op(n11572) );
  mux2_1 U13299 ( .ip1(i_ssi_txftlr[0]), .ip2(n11572), .s(n11571), .op(n11575)
         );
  inv_1 U13300 ( .ip(n11573), .op(n11574) );
  mux2_1 U13301 ( .ip1(i_ssi_rxftlr[0]), .ip2(n11575), .s(n11574), .op(n11577)
         );
  nor2_1 U13302 ( .ip1(n11584), .ip2(i_ssi_ssi_txe_intr_n), .op(n11585) );
  not_ab_or_c_or_d U13303 ( .ip1(n11587), .ip2(i_ssi_risr[0]), .ip3(n11586), 
        .ip4(n11585), .op(n11604) );
  nand2_1 U13304 ( .ip1(n11674), .ip2(i_ssi_U_dff_rx_mem[112]), .op(n11596) );
  and2_1 U13305 ( .ip1(n11675), .ip2(i_ssi_U_dff_rx_mem[0]), .op(n11593) );
  nand2_1 U13306 ( .ip1(n11687), .ip2(i_ssi_U_dff_rx_mem[96]), .op(n11591) );
  nand2_1 U13307 ( .ip1(n11678), .ip2(i_ssi_U_dff_rx_mem[80]), .op(n11590) );
  nand2_1 U13308 ( .ip1(n11677), .ip2(i_ssi_U_dff_rx_mem[48]), .op(n11589) );
  nand2_1 U13309 ( .ip1(n11679), .ip2(i_ssi_U_dff_rx_mem[32]), .op(n11588) );
  nand4_1 U13310 ( .ip1(n11591), .ip2(n11590), .ip3(n11589), .ip4(n11588), 
        .op(n11592) );
  not_ab_or_c_or_d U13311 ( .ip1(i_ssi_U_dff_rx_mem[64]), .ip2(n11686), .ip3(
        n11593), .ip4(n11592), .op(n11595) );
  nand2_1 U13312 ( .ip1(n11676), .ip2(i_ssi_U_dff_rx_mem[16]), .op(n11594) );
  nand3_1 U13313 ( .ip1(n11596), .ip2(n11595), .ip3(n11594), .op(n11597) );
  nand2_1 U13314 ( .ip1(n11598), .ip2(n11597), .op(n11603) );
  nand2_1 U13315 ( .ip1(n11599), .ip2(i_ssi_U_regfile_rxflr[0]), .op(n11602)
         );
  nand2_1 U13316 ( .ip1(n11600), .ip2(i_ssi_imr[0]), .op(n11601) );
  or2_1 U13317 ( .ip1(n11605), .ip2(n11606), .op(n11609) );
  or2_1 U13318 ( .ip1(n11607), .ip2(n11606), .op(n11608) );
  nand2_1 U13319 ( .ip1(n11609), .ip2(n11608), .op(n11610) );
  nor2_1 U13320 ( .ip1(i_ssi_reg_addr[0]), .ip2(n11610), .op(n11611) );
  nand3_1 U13321 ( .ip1(i_ssi_ssi_rxo_intr_n), .ip2(i_ssi_ssi_rxu_intr_n), 
        .ip3(i_ssi_ssi_txo_intr_n), .op(n11619) );
  nor2_1 U13322 ( .ip1(n11614), .ip2(i_ssi_ssi_mst_intr_n), .op(n11618) );
  nor3_1 U13323 ( .ip1(n11616), .ip2(n11615), .ip3(i_ssi_ssi_rxo_intr_n), .op(
        n11617) );
  not_ab_or_c_or_d U13324 ( .ip1(n11620), .ip2(n11619), .ip3(n11618), .ip4(
        n11617), .op(n11621) );
  nand2_1 U13325 ( .ip1(i_ssi_prdata[0]), .ip2(n11697), .op(n11625) );
  nand2_1 U13326 ( .ip1(n11626), .ip2(n11625), .op(n4244) );
  nand2_1 U13327 ( .ip1(n11687), .ip2(i_ssi_U_dff_rx_mem[104]), .op(n11635) );
  and2_1 U13328 ( .ip1(n11675), .ip2(i_ssi_U_dff_rx_mem[8]), .op(n11632) );
  nand2_1 U13329 ( .ip1(n11678), .ip2(i_ssi_U_dff_rx_mem[88]), .op(n11630) );
  nand2_1 U13330 ( .ip1(n11674), .ip2(i_ssi_U_dff_rx_mem[120]), .op(n11629) );
  nand2_1 U13331 ( .ip1(n11676), .ip2(i_ssi_U_dff_rx_mem[24]), .op(n11628) );
  nand2_1 U13332 ( .ip1(n11686), .ip2(i_ssi_U_dff_rx_mem[72]), .op(n11627) );
  nand4_1 U13333 ( .ip1(n11630), .ip2(n11629), .ip3(n11628), .ip4(n11627), 
        .op(n11631) );
  not_ab_or_c_or_d U13334 ( .ip1(i_ssi_U_dff_rx_mem[56]), .ip2(n11677), .ip3(
        n11632), .ip4(n11631), .op(n11634) );
  nand2_1 U13335 ( .ip1(n11679), .ip2(i_ssi_U_dff_rx_mem[40]), .op(n11633) );
  nand3_1 U13336 ( .ip1(n11635), .ip2(n11634), .ip3(n11633), .op(n11642) );
  inv_1 U13337 ( .ip(n11636), .op(n11700) );
  nand2_1 U13338 ( .ip1(i_ssi_baudr[8]), .ip2(n11691), .op(n11639) );
  nand2_1 U13339 ( .ip1(i_ssi_tmod[0]), .ip2(n11692), .op(n11638) );
  nand2_1 U13340 ( .ip1(n5393), .ip2(n11693), .op(n11637) );
  nand3_1 U13341 ( .ip1(n11639), .ip2(n11638), .ip3(n11637), .op(n11640) );
  mux2_1 U13342 ( .ip1(n11640), .ip2(i_ssi_prdata[8]), .s(n11697), .op(n11641)
         );
  ab_or_c_or_d U13343 ( .ip1(n11782), .ip2(n11642), .ip3(n11700), .ip4(n11641), 
        .op(n4236) );
  nand2_1 U13344 ( .ip1(n11674), .ip2(i_ssi_U_dff_rx_mem[121]), .op(n11651) );
  and2_1 U13345 ( .ip1(n11675), .ip2(i_ssi_U_dff_rx_mem[9]), .op(n11648) );
  nand2_1 U13346 ( .ip1(n11679), .ip2(i_ssi_U_dff_rx_mem[41]), .op(n11646) );
  nand2_1 U13347 ( .ip1(n11677), .ip2(i_ssi_U_dff_rx_mem[57]), .op(n11645) );
  nand2_1 U13348 ( .ip1(n11676), .ip2(i_ssi_U_dff_rx_mem[25]), .op(n11644) );
  nand2_1 U13349 ( .ip1(n11687), .ip2(i_ssi_U_dff_rx_mem[105]), .op(n11643) );
  nand4_1 U13350 ( .ip1(n11646), .ip2(n11645), .ip3(n11644), .ip4(n11643), 
        .op(n11647) );
  not_ab_or_c_or_d U13351 ( .ip1(i_ssi_U_dff_rx_mem[89]), .ip2(n11678), .ip3(
        n11648), .ip4(n11647), .op(n11650) );
  nand2_1 U13352 ( .ip1(n11686), .ip2(i_ssi_U_dff_rx_mem[73]), .op(n11649) );
  nand3_1 U13353 ( .ip1(n11651), .ip2(n11650), .ip3(n11649), .op(n11658) );
  nand2_1 U13354 ( .ip1(i_ssi_U_regfile_ctrlr1_int[9]), .ip2(n11693), .op(
        n11653) );
  nand3_1 U13355 ( .ip1(n11655), .ip2(n11654), .ip3(n11653), .op(n11656) );
  mux2_1 U13356 ( .ip1(n11656), .ip2(i_ssi_prdata[9]), .s(n11697), .op(n11657)
         );
  ab_or_c_or_d U13357 ( .ip1(n11782), .ip2(n11658), .ip3(n11700), .ip4(n11657), 
        .op(n4235) );
  nand2_1 U13358 ( .ip1(n11674), .ip2(i_ssi_U_dff_rx_mem[124]), .op(n11667) );
  and2_1 U13359 ( .ip1(n11675), .ip2(i_ssi_U_dff_rx_mem[12]), .op(n11664) );
  nand2_1 U13360 ( .ip1(n11676), .ip2(i_ssi_U_dff_rx_mem[28]), .op(n11662) );
  nand2_1 U13361 ( .ip1(n11677), .ip2(i_ssi_U_dff_rx_mem[60]), .op(n11661) );
  nand2_1 U13362 ( .ip1(n11678), .ip2(i_ssi_U_dff_rx_mem[92]), .op(n11660) );
  nand2_1 U13363 ( .ip1(n11679), .ip2(i_ssi_U_dff_rx_mem[44]), .op(n11659) );
  nand4_1 U13364 ( .ip1(n11662), .ip2(n11661), .ip3(n11660), .ip4(n11659), 
        .op(n11663) );
  not_ab_or_c_or_d U13365 ( .ip1(i_ssi_U_dff_rx_mem[108]), .ip2(n11687), .ip3(
        n11664), .ip4(n11663), .op(n11666) );
  nand2_1 U13366 ( .ip1(n11686), .ip2(i_ssi_U_dff_rx_mem[76]), .op(n11665) );
  nand3_1 U13367 ( .ip1(n11667), .ip2(n11666), .ip3(n11665), .op(n11673) );
  nand2_1 U13368 ( .ip1(i_ssi_baudr[12]), .ip2(n11691), .op(n11670) );
  nand2_1 U13369 ( .ip1(i_ssi_cfs[0]), .ip2(n11692), .op(n11669) );
  nand2_1 U13370 ( .ip1(i_ssi_U_regfile_ctrlr1_int[12]), .ip2(n11693), .op(
        n11668) );
  nand3_1 U13371 ( .ip1(n11670), .ip2(n11669), .ip3(n11668), .op(n11671) );
  mux2_1 U13372 ( .ip1(n11671), .ip2(i_ssi_prdata[12]), .s(n11697), .op(n11672) );
  ab_or_c_or_d U13373 ( .ip1(n11782), .ip2(n11673), .ip3(n11700), .ip4(n11672), 
        .op(n4232) );
  nand2_1 U13374 ( .ip1(n11674), .ip2(i_ssi_U_dff_rx_mem[125]), .op(n11690) );
  and2_1 U13375 ( .ip1(n11675), .ip2(i_ssi_U_dff_rx_mem[13]), .op(n11685) );
  nand2_1 U13376 ( .ip1(n11676), .ip2(i_ssi_U_dff_rx_mem[29]), .op(n11683) );
  nand2_1 U13377 ( .ip1(n11677), .ip2(i_ssi_U_dff_rx_mem[61]), .op(n11682) );
  nand2_1 U13378 ( .ip1(n11678), .ip2(i_ssi_U_dff_rx_mem[93]), .op(n11681) );
  nand2_1 U13379 ( .ip1(n11679), .ip2(i_ssi_U_dff_rx_mem[45]), .op(n11680) );
  nand4_1 U13380 ( .ip1(n11683), .ip2(n11682), .ip3(n11681), .ip4(n11680), 
        .op(n11684) );
  not_ab_or_c_or_d U13381 ( .ip1(i_ssi_U_dff_rx_mem[77]), .ip2(n11686), .ip3(
        n11685), .ip4(n11684), .op(n11689) );
  nand2_1 U13382 ( .ip1(n11687), .ip2(i_ssi_U_dff_rx_mem[109]), .op(n11688) );
  nand3_1 U13383 ( .ip1(n11690), .ip2(n11689), .ip3(n11688), .op(n11701) );
  nand2_1 U13384 ( .ip1(i_ssi_baudr[13]), .ip2(n11691), .op(n11696) );
  nand2_1 U13385 ( .ip1(i_ssi_cfs[1]), .ip2(n11692), .op(n11695) );
  nand2_1 U13386 ( .ip1(i_ssi_U_regfile_ctrlr1_int[13]), .ip2(n11693), .op(
        n11694) );
  nand3_1 U13387 ( .ip1(n11696), .ip2(n11695), .ip3(n11694), .op(n11698) );
  mux2_1 U13388 ( .ip1(n11698), .ip2(i_ssi_prdata[13]), .s(n11697), .op(n11699) );
  ab_or_c_or_d U13389 ( .ip1(n11782), .ip2(n11701), .ip3(n11700), .ip4(n11699), 
        .op(n4231) );
  nand3_1 U13390 ( .ip1(n11702), .ip2(i_ssi_U_mstfsm_ctrl_cnt[0]), .ip3(
        i_ssi_U_mstfsm_ctrl_cnt[1]), .op(n11707) );
  inv_1 U13391 ( .ip(n11707), .op(n11703) );
  not_ab_or_c_or_d U13392 ( .ip1(n11705), .ip2(n11704), .ip3(n11703), .ip4(
        n11708), .op(n4204) );
  nor2_1 U13393 ( .ip1(n11707), .ip2(n11706), .op(n11710) );
  not_ab_or_c_or_d U13394 ( .ip1(n11707), .ip2(n11706), .ip3(n11710), .ip4(
        n11708), .op(n4203) );
  nor2_1 U13395 ( .ip1(i_ssi_U_mstfsm_ctrl_cnt[3]), .ip2(n11710), .op(n11709)
         );
  not_ab_or_c_or_d U13396 ( .ip1(i_ssi_U_mstfsm_ctrl_cnt[3]), .ip2(n11710), 
        .ip3(n11709), .ip4(n11708), .op(n4202) );
  nand2_1 U13397 ( .ip1(n11711), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[0]), .op(n11716) );
  inv_1 U13398 ( .ip(n11716), .op(n11712) );
  not_ab_or_c_or_d U13399 ( .ip1(n11714), .ip2(n11713), .ip3(n11721), .ip4(
        n11712), .op(n4176) );
  not_ab_or_c_or_d U13400 ( .ip1(n11716), .ip2(n11715), .ip3(n11721), .ip4(
        n11717), .op(n4175) );
  not_ab_or_c_or_d U13401 ( .ip1(n11719), .ip2(n11718), .ip3(n11721), .ip4(
        n11722), .op(n4174) );
  nor2_1 U13402 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[3]), .ip2(
        n11722), .op(n11720) );
  not_ab_or_c_or_d U13403 ( .ip1(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[3]), .ip2(n11722), .ip3(
        n11721), .ip4(n11720), .op(n4173) );
  nor2_1 U13404 ( .ip1(i_i2c_p_det), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_count_en), 
        .op(n11723) );
  nor2_1 U13405 ( .ip1(i_i2c_s_det), .ip2(n11723), .op(n4125) );
endmodule

