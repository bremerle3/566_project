
module system_top ( HCLK_top, HRESETn_top, SYSRESETREQ_top_out, LOCKUP_top_out, 
        TXEV_top_out );
  input HCLK_top, HRESETn_top;
  output SYSRESETREQ_top_out, LOCKUP_top_out, TXEV_top_out;
  wire   HREADY_top, PID_hmastlock_top, \PID_htrans_top[1] , PID_hwrite_top,
         RAM_hready_resp_top, \RAM_hresp_top[0] , RAM_hsel_top,
         i_ssi_ssi_clk_top, i_ssi_ssi_rst_n_top, i_ssi_sclk_out_top,
         i_ssi_ss_0_n_top, i_ssi_ssi_mst_intr_n_top, i_ssi_ssi_oe_n_top,
         i_ssi_ssi_rxf_intr_n_top, i_ssi_ssi_rxo_intr_n_top,
         i_ssi_ssi_rxu_intr_n_top, i_ssi_ssi_sleep_top,
         i_ssi_ssi_txe_intr_n_top, i_ssi_ssi_intr_n_top, i_ssi_txd_top,
         \interconnect_ip_inst/n5991 , \interconnect_ip_inst/n6491 ,
         \interconnect_ip_inst/i_apb_hready_resp ,
         \interconnect_ip_inst/n4829 , \interconnect_ip_inst/i_ssi_fsm_sleep ,
         \interconnect_ip_inst/i_ssi_U_mstfsm_c_state[3] ,
         \interconnect_ip_inst/n4860 , \interconnect_ip_inst/n4861 ,
         \interconnect_ip_inst/n4862 , \interconnect_ip_inst/n4863 ,
         \interconnect_ip_inst/n4864 ,
         \interconnect_ip_inst/i_ahb_hresp_none_0_ ,
         \interconnect_ip_inst/i_ahb_U_dfltslv_N4 ,
         \interconnect_ip_inst/i_ahb_U_dfltslv_current_state ,
         \interconnect_ip_inst/n10765 , \interconnect_ip_inst/n11572 ,
         \CORTEXM0DS_INST/cm0_primask[0] , \CORTEXM0DS_INST/cm0_control[1] ,
         \CORTEXM0DS_INST/cm0_xpsr[24] , \CORTEXM0DS_INST/u_logic/N4816 ,
         \CORTEXM0DS_INST/u_logic/N4767 , \CORTEXM0DS_INST/u_logic/N4751 ,
         \CORTEXM0DS_INST/u_logic/N4674 , \CORTEXM0DS_INST/u_logic/N4518 ,
         \CORTEXM0DS_INST/u_logic/N4439 , \CORTEXM0DS_INST/u_logic/N4422 ,
         \CORTEXM0DS_INST/u_logic/N4421 , \CORTEXM0DS_INST/u_logic/N4396 ,
         \CORTEXM0DS_INST/u_logic/N4359 , \CORTEXM0DS_INST/u_logic/N4282 ,
         \CORTEXM0DS_INST/u_logic/N4227 , \CORTEXM0DS_INST/u_logic/N4170 ,
         \CORTEXM0DS_INST/u_logic/N4116 , \CORTEXM0DS_INST/u_logic/N4005 ,
         \CORTEXM0DS_INST/u_logic/N3967 , \CORTEXM0DS_INST/u_logic/N3966 ,
         \CORTEXM0DS_INST/u_logic/N3946 , \CORTEXM0DS_INST/u_logic/N3783 ,
         \CORTEXM0DS_INST/u_logic/N2678 , \CORTEXM0DS_INST/u_logic/N1447 ,
         \CORTEXM0DS_INST/u_logic/N586 , \CORTEXM0DS_INST/u_logic/E562z4 ,
         \CORTEXM0DS_INST/u_logic/Q462z4 , \CORTEXM0DS_INST/u_logic/A362z4 ,
         \CORTEXM0DS_INST/u_logic/Oq42z4 , \CORTEXM0DS_INST/u_logic/Xmywx4 ,
         \CORTEXM0DS_INST/u_logic/Ldhvx4 , \CORTEXM0DS_INST/u_logic/Sdhvx4 ,
         \CORTEXM0DS_INST/u_logic/Zdhvx4 , \CORTEXM0DS_INST/u_logic/Gehvx4 ,
         \CORTEXM0DS_INST/u_logic/Nehvx4 , \CORTEXM0DS_INST/u_logic/Uehvx4 ,
         \CORTEXM0DS_INST/u_logic/Bfhvx4 , \CORTEXM0DS_INST/u_logic/Ifhvx4 ,
         \CORTEXM0DS_INST/u_logic/Pfhvx4 , \CORTEXM0DS_INST/u_logic/Wfhvx4 ,
         \CORTEXM0DS_INST/u_logic/Dghvx4 , \CORTEXM0DS_INST/u_logic/Rghvx4 ,
         \CORTEXM0DS_INST/u_logic/Mhhvx4 , \CORTEXM0DS_INST/u_logic/Thhvx4 ,
         \CORTEXM0DS_INST/u_logic/Aihvx4 , \CORTEXM0DS_INST/u_logic/Hihvx4 ,
         \CORTEXM0DS_INST/u_logic/Oihvx4 , \CORTEXM0DS_INST/u_logic/Vihvx4 ,
         \CORTEXM0DS_INST/u_logic/Cjhvx4 , \CORTEXM0DS_INST/u_logic/Jjhvx4 ,
         \CORTEXM0DS_INST/u_logic/Qjhvx4 , \CORTEXM0DS_INST/u_logic/Xjhvx4 ,
         \CORTEXM0DS_INST/u_logic/Ekhvx4 , \CORTEXM0DS_INST/u_logic/Lkhvx4 ,
         \CORTEXM0DS_INST/u_logic/Skhvx4 , \CORTEXM0DS_INST/u_logic/Zkhvx4 ,
         \CORTEXM0DS_INST/u_logic/Glhvx4 , \CORTEXM0DS_INST/u_logic/Nlhvx4 ,
         \CORTEXM0DS_INST/u_logic/Ulhvx4 , \CORTEXM0DS_INST/u_logic/Bmhvx4 ,
         \CORTEXM0DS_INST/u_logic/Imhvx4 , \CORTEXM0DS_INST/u_logic/Lrhvx4 ,
         \CORTEXM0DS_INST/u_logic/Ithvx4 , \CORTEXM0DS_INST/u_logic/Pthvx4 ,
         \CORTEXM0DS_INST/u_logic/Wthvx4 , \CORTEXM0DS_INST/u_logic/Duhvx4 ,
         \CORTEXM0DS_INST/u_logic/Kuhvx4 , \CORTEXM0DS_INST/u_logic/Ruhvx4 ,
         \CORTEXM0DS_INST/u_logic/Yuhvx4 , \CORTEXM0DS_INST/u_logic/Fvhvx4 ,
         \CORTEXM0DS_INST/u_logic/Mvhvx4 , \CORTEXM0DS_INST/u_logic/Tvhvx4 ,
         \CORTEXM0DS_INST/u_logic/Awhvx4 , \CORTEXM0DS_INST/u_logic/Hwhvx4 ,
         \CORTEXM0DS_INST/u_logic/Owhvx4 , \CORTEXM0DS_INST/u_logic/Vwhvx4 ,
         \CORTEXM0DS_INST/u_logic/Cxhvx4 , \CORTEXM0DS_INST/u_logic/Jxhvx4 ,
         \CORTEXM0DS_INST/u_logic/Qxhvx4 , \CORTEXM0DS_INST/u_logic/Xxhvx4 ,
         \CORTEXM0DS_INST/u_logic/Eyhvx4 , \CORTEXM0DS_INST/u_logic/Lyhvx4 ,
         \CORTEXM0DS_INST/u_logic/Bq5wx4 , \CORTEXM0DS_INST/u_logic/Owgvx4 ,
         \CORTEXM0DS_INST/u_logic/T2ivx4 , \CORTEXM0DS_INST/u_logic/F2ivx4 ,
         \CORTEXM0DS_INST/u_logic/Y1ivx4 , \CORTEXM0DS_INST/u_logic/M2ivx4 ,
         \CORTEXM0DS_INST/u_logic/K1ivx4 , \CORTEXM0DS_INST/u_logic/D1ivx4 ,
         \CORTEXM0DS_INST/u_logic/R1ivx4 , \CORTEXM0DS_INST/u_logic/P0ivx4 ,
         \CORTEXM0DS_INST/u_logic/I0ivx4 , \CORTEXM0DS_INST/u_logic/W0ivx4 ,
         \CORTEXM0DS_INST/u_logic/B0ivx4 , \CORTEXM0DS_INST/u_logic/Uzhvx4 ,
         \CORTEXM0DS_INST/u_logic/Gzhvx4 , \CORTEXM0DS_INST/u_logic/Zyhvx4 ,
         \CORTEXM0DS_INST/u_logic/Nzhvx4 , \CORTEXM0DS_INST/u_logic/Syhvx4 ,
         \CORTEXM0DS_INST/u_logic/O24wx4 , \CORTEXM0DS_INST/u_logic/Sx3wx4 ,
         \CORTEXM0DS_INST/u_logic/H3ivx4 , \CORTEXM0DS_INST/u_logic/V3ivx4 ,
         \CORTEXM0DS_INST/u_logic/C4ivx4 , \CORTEXM0DS_INST/u_logic/J4ivx4 ,
         \CORTEXM0DS_INST/u_logic/Q4ivx4 , \CORTEXM0DS_INST/u_logic/X4ivx4 ,
         \CORTEXM0DS_INST/u_logic/E5ivx4 , \CORTEXM0DS_INST/u_logic/L5ivx4 ,
         \CORTEXM0DS_INST/u_logic/S5ivx4 , \CORTEXM0DS_INST/u_logic/Z5ivx4 ,
         \CORTEXM0DS_INST/u_logic/G6ivx4 , \CORTEXM0DS_INST/u_logic/N6ivx4 ,
         \CORTEXM0DS_INST/u_logic/U6ivx4 , \CORTEXM0DS_INST/u_logic/B7ivx4 ,
         \CORTEXM0DS_INST/u_logic/I7ivx4 , \CORTEXM0DS_INST/u_logic/P7ivx4 ,
         \CORTEXM0DS_INST/u_logic/W7ivx4 , \CORTEXM0DS_INST/u_logic/D8ivx4 ,
         \CORTEXM0DS_INST/u_logic/Y92wx4 , \CORTEXM0DS_INST/u_logic/R8ivx4 ,
         \CORTEXM0DS_INST/u_logic/Y8ivx4 , \CORTEXM0DS_INST/u_logic/F9ivx4 ,
         \CORTEXM0DS_INST/u_logic/M9ivx4 , \CORTEXM0DS_INST/u_logic/T9ivx4 ,
         \CORTEXM0DS_INST/u_logic/Aaivx4 , \CORTEXM0DS_INST/u_logic/Haivx4 ,
         \CORTEXM0DS_INST/u_logic/Oaivx4 , \CORTEXM0DS_INST/u_logic/Vaivx4 ,
         \CORTEXM0DS_INST/u_logic/Cbivx4 , \CORTEXM0DS_INST/u_logic/Jbivx4 ,
         \CORTEXM0DS_INST/u_logic/Qbivx4 , \CORTEXM0DS_INST/u_logic/Xbivx4 ,
         \CORTEXM0DS_INST/u_logic/Ecivx4 , \CORTEXM0DS_INST/u_logic/Lcivx4 ,
         \CORTEXM0DS_INST/u_logic/Scivx4 , \CORTEXM0DS_INST/u_logic/Gdivx4 ,
         \CORTEXM0DS_INST/u_logic/Ndivx4 , \CORTEXM0DS_INST/u_logic/Udivx4 ,
         \CORTEXM0DS_INST/u_logic/Beivx4 , \CORTEXM0DS_INST/u_logic/Ieivx4 ,
         \CORTEXM0DS_INST/u_logic/Peivx4 , \CORTEXM0DS_INST/u_logic/Weivx4 ,
         \CORTEXM0DS_INST/u_logic/Dfivx4 , \CORTEXM0DS_INST/u_logic/Kfivx4 ,
         \CORTEXM0DS_INST/u_logic/Rfivx4 , \CORTEXM0DS_INST/u_logic/Yfivx4 ,
         \CORTEXM0DS_INST/u_logic/Fgivx4 , \CORTEXM0DS_INST/u_logic/Mgivx4 ,
         \CORTEXM0DS_INST/u_logic/Tgivx4 , \CORTEXM0DS_INST/u_logic/Ahivx4 ,
         \CORTEXM0DS_INST/u_logic/Hhivx4 , \CORTEXM0DS_INST/u_logic/Vhivx4 ,
         \CORTEXM0DS_INST/u_logic/Ciivx4 , \CORTEXM0DS_INST/u_logic/Jiivx4 ,
         \CORTEXM0DS_INST/u_logic/Qiivx4 , \CORTEXM0DS_INST/u_logic/Xiivx4 ,
         \CORTEXM0DS_INST/u_logic/Ejivx4 , \CORTEXM0DS_INST/u_logic/Ljivx4 ,
         \CORTEXM0DS_INST/u_logic/Sjivx4 , \CORTEXM0DS_INST/u_logic/Zjivx4 ,
         \CORTEXM0DS_INST/u_logic/Gkivx4 , \CORTEXM0DS_INST/u_logic/Nkivx4 ,
         \CORTEXM0DS_INST/u_logic/Ukivx4 , \CORTEXM0DS_INST/u_logic/Blivx4 ,
         \CORTEXM0DS_INST/u_logic/Ilivx4 , \CORTEXM0DS_INST/u_logic/Plivx4 ,
         \CORTEXM0DS_INST/u_logic/Wlivx4 , \CORTEXM0DS_INST/u_logic/Kmivx4 ,
         \CORTEXM0DS_INST/u_logic/Rmivx4 , \CORTEXM0DS_INST/u_logic/Ymivx4 ,
         \CORTEXM0DS_INST/u_logic/Fnivx4 , \CORTEXM0DS_INST/u_logic/Mnivx4 ,
         \CORTEXM0DS_INST/u_logic/Tnivx4 , \CORTEXM0DS_INST/u_logic/Aoivx4 ,
         \CORTEXM0DS_INST/u_logic/Hoivx4 , \CORTEXM0DS_INST/u_logic/Ooivx4 ,
         \CORTEXM0DS_INST/u_logic/Voivx4 , \CORTEXM0DS_INST/u_logic/Cpivx4 ,
         \CORTEXM0DS_INST/u_logic/Jpivx4 , \CORTEXM0DS_INST/u_logic/Qpivx4 ,
         \CORTEXM0DS_INST/u_logic/Xpivx4 , \CORTEXM0DS_INST/u_logic/Eqivx4 ,
         \CORTEXM0DS_INST/u_logic/Lqivx4 , \CORTEXM0DS_INST/u_logic/Sqivx4 ,
         \CORTEXM0DS_INST/u_logic/Zqivx4 , \CORTEXM0DS_INST/u_logic/Grivx4 ,
         \CORTEXM0DS_INST/u_logic/Nrivx4 , \CORTEXM0DS_INST/u_logic/Urivx4 ,
         \CORTEXM0DS_INST/u_logic/Bsivx4 , \CORTEXM0DS_INST/u_logic/Isivx4 ,
         \CORTEXM0DS_INST/u_logic/Psivx4 , \CORTEXM0DS_INST/u_logic/Wsivx4 ,
         \CORTEXM0DS_INST/u_logic/Dtivx4 , \CORTEXM0DS_INST/u_logic/Ktivx4 ,
         \CORTEXM0DS_INST/u_logic/Rtivx4 , \CORTEXM0DS_INST/u_logic/Ytivx4 ,
         \CORTEXM0DS_INST/u_logic/Fuivx4 , \CORTEXM0DS_INST/u_logic/Muivx4 ,
         \CORTEXM0DS_INST/u_logic/Tuivx4 , \CORTEXM0DS_INST/u_logic/Avivx4 ,
         \CORTEXM0DS_INST/u_logic/Ovivx4 , \CORTEXM0DS_INST/u_logic/Vvivx4 ,
         \CORTEXM0DS_INST/u_logic/Cwivx4 , \CORTEXM0DS_INST/u_logic/Jwivx4 ,
         \CORTEXM0DS_INST/u_logic/Qwivx4 , \CORTEXM0DS_INST/u_logic/Xwivx4 ,
         \CORTEXM0DS_INST/u_logic/Exivx4 , \CORTEXM0DS_INST/u_logic/Lxivx4 ,
         \CORTEXM0DS_INST/u_logic/Sxivx4 , \CORTEXM0DS_INST/u_logic/Zxivx4 ,
         \CORTEXM0DS_INST/u_logic/Gyivx4 , \CORTEXM0DS_INST/u_logic/Nyivx4 ,
         \CORTEXM0DS_INST/u_logic/Uyivx4 , \CORTEXM0DS_INST/u_logic/Bzivx4 ,
         \CORTEXM0DS_INST/u_logic/Izivx4 , \CORTEXM0DS_INST/u_logic/Pzivx4 ,
         \CORTEXM0DS_INST/u_logic/D0jvx4 , \CORTEXM0DS_INST/u_logic/K0jvx4 ,
         \CORTEXM0DS_INST/u_logic/R0jvx4 , \CORTEXM0DS_INST/u_logic/Y0jvx4 ,
         \CORTEXM0DS_INST/u_logic/F1jvx4 , \CORTEXM0DS_INST/u_logic/M1jvx4 ,
         \CORTEXM0DS_INST/u_logic/T1jvx4 , \CORTEXM0DS_INST/u_logic/A2jvx4 ,
         \CORTEXM0DS_INST/u_logic/H2jvx4 , \CORTEXM0DS_INST/u_logic/O2jvx4 ,
         \CORTEXM0DS_INST/u_logic/V2jvx4 , \CORTEXM0DS_INST/u_logic/C3jvx4 ,
         \CORTEXM0DS_INST/u_logic/J3jvx4 , \CORTEXM0DS_INST/u_logic/Q3jvx4 ,
         \CORTEXM0DS_INST/u_logic/X3jvx4 , \CORTEXM0DS_INST/u_logic/E4jvx4 ,
         \CORTEXM0DS_INST/u_logic/S4jvx4 , \CORTEXM0DS_INST/u_logic/Z4jvx4 ,
         \CORTEXM0DS_INST/u_logic/G5jvx4 , \CORTEXM0DS_INST/u_logic/N5jvx4 ,
         \CORTEXM0DS_INST/u_logic/U5jvx4 , \CORTEXM0DS_INST/u_logic/B6jvx4 ,
         \CORTEXM0DS_INST/u_logic/I6jvx4 , \CORTEXM0DS_INST/u_logic/P6jvx4 ,
         \CORTEXM0DS_INST/u_logic/W6jvx4 , \CORTEXM0DS_INST/u_logic/D7jvx4 ,
         \CORTEXM0DS_INST/u_logic/K7jvx4 , \CORTEXM0DS_INST/u_logic/R7jvx4 ,
         \CORTEXM0DS_INST/u_logic/Y7jvx4 , \CORTEXM0DS_INST/u_logic/F8jvx4 ,
         \CORTEXM0DS_INST/u_logic/M8jvx4 , \CORTEXM0DS_INST/u_logic/T8jvx4 ,
         \CORTEXM0DS_INST/u_logic/H9jvx4 , \CORTEXM0DS_INST/u_logic/O9jvx4 ,
         \CORTEXM0DS_INST/u_logic/V9jvx4 , \CORTEXM0DS_INST/u_logic/Cajvx4 ,
         \CORTEXM0DS_INST/u_logic/Jajvx4 , \CORTEXM0DS_INST/u_logic/Qajvx4 ,
         \CORTEXM0DS_INST/u_logic/Xajvx4 , \CORTEXM0DS_INST/u_logic/Ebjvx4 ,
         \CORTEXM0DS_INST/u_logic/Lbjvx4 , \CORTEXM0DS_INST/u_logic/Sbjvx4 ,
         \CORTEXM0DS_INST/u_logic/Zbjvx4 , \CORTEXM0DS_INST/u_logic/Gcjvx4 ,
         \CORTEXM0DS_INST/u_logic/Ncjvx4 , \CORTEXM0DS_INST/u_logic/Ucjvx4 ,
         \CORTEXM0DS_INST/u_logic/Bdjvx4 , \CORTEXM0DS_INST/u_logic/Idjvx4 ,
         \CORTEXM0DS_INST/u_logic/Wdjvx4 , \CORTEXM0DS_INST/u_logic/Dejvx4 ,
         \CORTEXM0DS_INST/u_logic/Kejvx4 , \CORTEXM0DS_INST/u_logic/Rejvx4 ,
         \CORTEXM0DS_INST/u_logic/Yejvx4 , \CORTEXM0DS_INST/u_logic/Ffjvx4 ,
         \CORTEXM0DS_INST/u_logic/Mfjvx4 , \CORTEXM0DS_INST/u_logic/Tfjvx4 ,
         \CORTEXM0DS_INST/u_logic/Agjvx4 , \CORTEXM0DS_INST/u_logic/Hgjvx4 ,
         \CORTEXM0DS_INST/u_logic/Ogjvx4 , \CORTEXM0DS_INST/u_logic/Vgjvx4 ,
         \CORTEXM0DS_INST/u_logic/Chjvx4 , \CORTEXM0DS_INST/u_logic/Jhjvx4 ,
         \CORTEXM0DS_INST/u_logic/Qhjvx4 , \CORTEXM0DS_INST/u_logic/Xhjvx4 ,
         \CORTEXM0DS_INST/u_logic/Lijvx4 , \CORTEXM0DS_INST/u_logic/Sijvx4 ,
         \CORTEXM0DS_INST/u_logic/Zijvx4 , \CORTEXM0DS_INST/u_logic/Gjjvx4 ,
         \CORTEXM0DS_INST/u_logic/Njjvx4 , \CORTEXM0DS_INST/u_logic/Ujjvx4 ,
         \CORTEXM0DS_INST/u_logic/Bkjvx4 , \CORTEXM0DS_INST/u_logic/Ikjvx4 ,
         \CORTEXM0DS_INST/u_logic/Pkjvx4 , \CORTEXM0DS_INST/u_logic/Wkjvx4 ,
         \CORTEXM0DS_INST/u_logic/Dljvx4 , \CORTEXM0DS_INST/u_logic/Kljvx4 ,
         \CORTEXM0DS_INST/u_logic/Rljvx4 , \CORTEXM0DS_INST/u_logic/Yljvx4 ,
         \CORTEXM0DS_INST/u_logic/Fmjvx4 , \CORTEXM0DS_INST/u_logic/Mmjvx4 ,
         \CORTEXM0DS_INST/u_logic/Bv0wx4 , \CORTEXM0DS_INST/u_logic/Anjvx4 ,
         \CORTEXM0DS_INST/u_logic/Hnjvx4 , \CORTEXM0DS_INST/u_logic/Onjvx4 ,
         \CORTEXM0DS_INST/u_logic/Vnjvx4 , \CORTEXM0DS_INST/u_logic/Cojvx4 ,
         \CORTEXM0DS_INST/u_logic/Jojvx4 , \CORTEXM0DS_INST/u_logic/Qojvx4 ,
         \CORTEXM0DS_INST/u_logic/Xojvx4 , \CORTEXM0DS_INST/u_logic/Epjvx4 ,
         \CORTEXM0DS_INST/u_logic/Lpjvx4 , \CORTEXM0DS_INST/u_logic/Spjvx4 ,
         \CORTEXM0DS_INST/u_logic/Zpjvx4 , \CORTEXM0DS_INST/u_logic/Gqjvx4 ,
         \CORTEXM0DS_INST/u_logic/Nqjvx4 , \CORTEXM0DS_INST/u_logic/Uqjvx4 ,
         \CORTEXM0DS_INST/u_logic/Brjvx4 , \CORTEXM0DS_INST/u_logic/Fq0wx4 ,
         \CORTEXM0DS_INST/u_logic/Prjvx4 , \CORTEXM0DS_INST/u_logic/Wrjvx4 ,
         \CORTEXM0DS_INST/u_logic/Dsjvx4 , \CORTEXM0DS_INST/u_logic/Ksjvx4 ,
         \CORTEXM0DS_INST/u_logic/Rsjvx4 , \CORTEXM0DS_INST/u_logic/Ysjvx4 ,
         \CORTEXM0DS_INST/u_logic/Ftjvx4 , \CORTEXM0DS_INST/u_logic/Mtjvx4 ,
         \CORTEXM0DS_INST/u_logic/Ttjvx4 , \CORTEXM0DS_INST/u_logic/Aujvx4 ,
         \CORTEXM0DS_INST/u_logic/Hujvx4 , \CORTEXM0DS_INST/u_logic/Oujvx4 ,
         \CORTEXM0DS_INST/u_logic/Vujvx4 , \CORTEXM0DS_INST/u_logic/Cvjvx4 ,
         \CORTEXM0DS_INST/u_logic/Jvjvx4 , \CORTEXM0DS_INST/u_logic/Qvjvx4 ,
         \CORTEXM0DS_INST/u_logic/Ql0wx4 , \CORTEXM0DS_INST/u_logic/Ewjvx4 ,
         \CORTEXM0DS_INST/u_logic/Lwjvx4 , \CORTEXM0DS_INST/u_logic/Swjvx4 ,
         \CORTEXM0DS_INST/u_logic/Zwjvx4 , \CORTEXM0DS_INST/u_logic/Gxjvx4 ,
         \CORTEXM0DS_INST/u_logic/Nxjvx4 , \CORTEXM0DS_INST/u_logic/Uxjvx4 ,
         \CORTEXM0DS_INST/u_logic/Byjvx4 , \CORTEXM0DS_INST/u_logic/Iyjvx4 ,
         \CORTEXM0DS_INST/u_logic/Pyjvx4 , \CORTEXM0DS_INST/u_logic/Wyjvx4 ,
         \CORTEXM0DS_INST/u_logic/Dzjvx4 , \CORTEXM0DS_INST/u_logic/Kzjvx4 ,
         \CORTEXM0DS_INST/u_logic/Rzjvx4 , \CORTEXM0DS_INST/u_logic/Yzjvx4 ,
         \CORTEXM0DS_INST/u_logic/F0kvx4 , \CORTEXM0DS_INST/u_logic/Ug0wx4 ,
         \CORTEXM0DS_INST/u_logic/T0kvx4 , \CORTEXM0DS_INST/u_logic/A1kvx4 ,
         \CORTEXM0DS_INST/u_logic/H1kvx4 , \CORTEXM0DS_INST/u_logic/O1kvx4 ,
         \CORTEXM0DS_INST/u_logic/V1kvx4 , \CORTEXM0DS_INST/u_logic/C2kvx4 ,
         \CORTEXM0DS_INST/u_logic/J2kvx4 , \CORTEXM0DS_INST/u_logic/Q2kvx4 ,
         \CORTEXM0DS_INST/u_logic/X2kvx4 , \CORTEXM0DS_INST/u_logic/E3kvx4 ,
         \CORTEXM0DS_INST/u_logic/L3kvx4 , \CORTEXM0DS_INST/u_logic/S3kvx4 ,
         \CORTEXM0DS_INST/u_logic/Z3kvx4 , \CORTEXM0DS_INST/u_logic/G4kvx4 ,
         \CORTEXM0DS_INST/u_logic/N4kvx4 , \CORTEXM0DS_INST/u_logic/U4kvx4 ,
         \CORTEXM0DS_INST/u_logic/Fc0wx4 , \CORTEXM0DS_INST/u_logic/I5kvx4 ,
         \CORTEXM0DS_INST/u_logic/P5kvx4 , \CORTEXM0DS_INST/u_logic/W5kvx4 ,
         \CORTEXM0DS_INST/u_logic/D6kvx4 , \CORTEXM0DS_INST/u_logic/K6kvx4 ,
         \CORTEXM0DS_INST/u_logic/R6kvx4 , \CORTEXM0DS_INST/u_logic/Y6kvx4 ,
         \CORTEXM0DS_INST/u_logic/F7kvx4 , \CORTEXM0DS_INST/u_logic/M7kvx4 ,
         \CORTEXM0DS_INST/u_logic/T7kvx4 , \CORTEXM0DS_INST/u_logic/A8kvx4 ,
         \CORTEXM0DS_INST/u_logic/H8kvx4 , \CORTEXM0DS_INST/u_logic/O8kvx4 ,
         \CORTEXM0DS_INST/u_logic/V8kvx4 , \CORTEXM0DS_INST/u_logic/C9kvx4 ,
         \CORTEXM0DS_INST/u_logic/J9kvx4 , \CORTEXM0DS_INST/u_logic/C70wx4 ,
         \CORTEXM0DS_INST/u_logic/X9kvx4 , \CORTEXM0DS_INST/u_logic/Eakvx4 ,
         \CORTEXM0DS_INST/u_logic/Lakvx4 , \CORTEXM0DS_INST/u_logic/Sakvx4 ,
         \CORTEXM0DS_INST/u_logic/Zakvx4 , \CORTEXM0DS_INST/u_logic/Gbkvx4 ,
         \CORTEXM0DS_INST/u_logic/Nbkvx4 , \CORTEXM0DS_INST/u_logic/Ubkvx4 ,
         \CORTEXM0DS_INST/u_logic/Bckvx4 , \CORTEXM0DS_INST/u_logic/Ickvx4 ,
         \CORTEXM0DS_INST/u_logic/Pckvx4 , \CORTEXM0DS_INST/u_logic/Wckvx4 ,
         \CORTEXM0DS_INST/u_logic/Ddkvx4 , \CORTEXM0DS_INST/u_logic/Kdkvx4 ,
         \CORTEXM0DS_INST/u_logic/Rdkvx4 , \CORTEXM0DS_INST/u_logic/Ydkvx4 ,
         \CORTEXM0DS_INST/u_logic/Fekvx4 , \CORTEXM0DS_INST/u_logic/Tekvx4 ,
         \CORTEXM0DS_INST/u_logic/Afkvx4 , \CORTEXM0DS_INST/u_logic/Hfkvx4 ,
         \CORTEXM0DS_INST/u_logic/Ofkvx4 , \CORTEXM0DS_INST/u_logic/Vfkvx4 ,
         \CORTEXM0DS_INST/u_logic/Cgkvx4 , \CORTEXM0DS_INST/u_logic/Jgkvx4 ,
         \CORTEXM0DS_INST/u_logic/Qgkvx4 , \CORTEXM0DS_INST/u_logic/Xgkvx4 ,
         \CORTEXM0DS_INST/u_logic/Ehkvx4 , \CORTEXM0DS_INST/u_logic/Lhkvx4 ,
         \CORTEXM0DS_INST/u_logic/Shkvx4 , \CORTEXM0DS_INST/u_logic/Zhkvx4 ,
         \CORTEXM0DS_INST/u_logic/Gikvx4 , \CORTEXM0DS_INST/u_logic/Nikvx4 ,
         \CORTEXM0DS_INST/u_logic/Uikvx4 , \CORTEXM0DS_INST/u_logic/Ijkvx4 ,
         \CORTEXM0DS_INST/u_logic/Pjkvx4 , \CORTEXM0DS_INST/u_logic/Wjkvx4 ,
         \CORTEXM0DS_INST/u_logic/Dkkvx4 , \CORTEXM0DS_INST/u_logic/Kkkvx4 ,
         \CORTEXM0DS_INST/u_logic/Rkkvx4 , \CORTEXM0DS_INST/u_logic/Ykkvx4 ,
         \CORTEXM0DS_INST/u_logic/Flkvx4 , \CORTEXM0DS_INST/u_logic/Mlkvx4 ,
         \CORTEXM0DS_INST/u_logic/Tlkvx4 , \CORTEXM0DS_INST/u_logic/Amkvx4 ,
         \CORTEXM0DS_INST/u_logic/Hmkvx4 , \CORTEXM0DS_INST/u_logic/Omkvx4 ,
         \CORTEXM0DS_INST/u_logic/Vmkvx4 , \CORTEXM0DS_INST/u_logic/Cnkvx4 ,
         \CORTEXM0DS_INST/u_logic/Jnkvx4 , \CORTEXM0DS_INST/u_logic/Rxzvx4 ,
         \CORTEXM0DS_INST/u_logic/Xnkvx4 , \CORTEXM0DS_INST/u_logic/Eokvx4 ,
         \CORTEXM0DS_INST/u_logic/Lokvx4 , \CORTEXM0DS_INST/u_logic/Sokvx4 ,
         \CORTEXM0DS_INST/u_logic/Zokvx4 , \CORTEXM0DS_INST/u_logic/Gpkvx4 ,
         \CORTEXM0DS_INST/u_logic/Npkvx4 , \CORTEXM0DS_INST/u_logic/Upkvx4 ,
         \CORTEXM0DS_INST/u_logic/Bqkvx4 , \CORTEXM0DS_INST/u_logic/Iqkvx4 ,
         \CORTEXM0DS_INST/u_logic/Pqkvx4 , \CORTEXM0DS_INST/u_logic/Wqkvx4 ,
         \CORTEXM0DS_INST/u_logic/Drkvx4 , \CORTEXM0DS_INST/u_logic/Krkvx4 ,
         \CORTEXM0DS_INST/u_logic/Rrkvx4 , \CORTEXM0DS_INST/u_logic/Yrkvx4 ,
         \CORTEXM0DS_INST/u_logic/Hszvx4 , \CORTEXM0DS_INST/u_logic/Mskvx4 ,
         \CORTEXM0DS_INST/u_logic/Tskvx4 , \CORTEXM0DS_INST/u_logic/Atkvx4 ,
         \CORTEXM0DS_INST/u_logic/Htkvx4 , \CORTEXM0DS_INST/u_logic/Otkvx4 ,
         \CORTEXM0DS_INST/u_logic/Vtkvx4 , \CORTEXM0DS_INST/u_logic/Cukvx4 ,
         \CORTEXM0DS_INST/u_logic/Jukvx4 , \CORTEXM0DS_INST/u_logic/Qukvx4 ,
         \CORTEXM0DS_INST/u_logic/Xukvx4 , \CORTEXM0DS_INST/u_logic/Evkvx4 ,
         \CORTEXM0DS_INST/u_logic/Lvkvx4 , \CORTEXM0DS_INST/u_logic/Svkvx4 ,
         \CORTEXM0DS_INST/u_logic/Zvkvx4 , \CORTEXM0DS_INST/u_logic/Gwkvx4 ,
         \CORTEXM0DS_INST/u_logic/Nwkvx4 , \CORTEXM0DS_INST/u_logic/Uwkvx4 ,
         \CORTEXM0DS_INST/u_logic/Bxkvx4 , \CORTEXM0DS_INST/u_logic/Ixkvx4 ,
         \CORTEXM0DS_INST/u_logic/Pxkvx4 , \CORTEXM0DS_INST/u_logic/Wxkvx4 ,
         \CORTEXM0DS_INST/u_logic/Dykvx4 , \CORTEXM0DS_INST/u_logic/Kykvx4 ,
         \CORTEXM0DS_INST/u_logic/Rykvx4 , \CORTEXM0DS_INST/u_logic/Yykvx4 ,
         \CORTEXM0DS_INST/u_logic/Fzkvx4 , \CORTEXM0DS_INST/u_logic/Mzkvx4 ,
         \CORTEXM0DS_INST/u_logic/Tzkvx4 , \CORTEXM0DS_INST/u_logic/A0lvx4 ,
         \CORTEXM0DS_INST/u_logic/H0lvx4 , \CORTEXM0DS_INST/u_logic/O0lvx4 ,
         \CORTEXM0DS_INST/u_logic/V0lvx4 , \CORTEXM0DS_INST/u_logic/J1lvx4 ,
         \CORTEXM0DS_INST/u_logic/Q1lvx4 , \CORTEXM0DS_INST/u_logic/X1lvx4 ,
         \CORTEXM0DS_INST/u_logic/E2lvx4 , \CORTEXM0DS_INST/u_logic/L2lvx4 ,
         \CORTEXM0DS_INST/u_logic/S2lvx4 , \CORTEXM0DS_INST/u_logic/Z2lvx4 ,
         \CORTEXM0DS_INST/u_logic/G3lvx4 , \CORTEXM0DS_INST/u_logic/N3lvx4 ,
         \CORTEXM0DS_INST/u_logic/U3lvx4 , \CORTEXM0DS_INST/u_logic/B4lvx4 ,
         \CORTEXM0DS_INST/u_logic/I4lvx4 , \CORTEXM0DS_INST/u_logic/P4lvx4 ,
         \CORTEXM0DS_INST/u_logic/W4lvx4 , \CORTEXM0DS_INST/u_logic/D5lvx4 ,
         \CORTEXM0DS_INST/u_logic/K5lvx4 , \CORTEXM0DS_INST/u_logic/Nhzvx4 ,
         \CORTEXM0DS_INST/u_logic/Y5lvx4 , \CORTEXM0DS_INST/u_logic/F6lvx4 ,
         \CORTEXM0DS_INST/u_logic/M6lvx4 , \CORTEXM0DS_INST/u_logic/T6lvx4 ,
         \CORTEXM0DS_INST/u_logic/A7lvx4 , \CORTEXM0DS_INST/u_logic/H7lvx4 ,
         \CORTEXM0DS_INST/u_logic/O7lvx4 , \CORTEXM0DS_INST/u_logic/V7lvx4 ,
         \CORTEXM0DS_INST/u_logic/C8lvx4 , \CORTEXM0DS_INST/u_logic/J8lvx4 ,
         \CORTEXM0DS_INST/u_logic/Q8lvx4 , \CORTEXM0DS_INST/u_logic/X8lvx4 ,
         \CORTEXM0DS_INST/u_logic/E9lvx4 , \CORTEXM0DS_INST/u_logic/L9lvx4 ,
         \CORTEXM0DS_INST/u_logic/S9lvx4 , \CORTEXM0DS_INST/u_logic/Z9lvx4 ,
         \CORTEXM0DS_INST/u_logic/Vezvx4 , \CORTEXM0DS_INST/u_logic/Nalvx4 ,
         \CORTEXM0DS_INST/u_logic/Ualvx4 , \CORTEXM0DS_INST/u_logic/Bblvx4 ,
         \CORTEXM0DS_INST/u_logic/Iblvx4 , \CORTEXM0DS_INST/u_logic/Pblvx4 ,
         \CORTEXM0DS_INST/u_logic/Wblvx4 , \CORTEXM0DS_INST/u_logic/Dclvx4 ,
         \CORTEXM0DS_INST/u_logic/Kclvx4 , \CORTEXM0DS_INST/u_logic/Rclvx4 ,
         \CORTEXM0DS_INST/u_logic/Yclvx4 , \CORTEXM0DS_INST/u_logic/Fdlvx4 ,
         \CORTEXM0DS_INST/u_logic/Mdlvx4 , \CORTEXM0DS_INST/u_logic/Tdlvx4 ,
         \CORTEXM0DS_INST/u_logic/Aelvx4 , \CORTEXM0DS_INST/u_logic/Helvx4 ,
         \CORTEXM0DS_INST/u_logic/Oelvx4 , \CORTEXM0DS_INST/u_logic/Cflvx4 ,
         \CORTEXM0DS_INST/u_logic/Jflvx4 , \CORTEXM0DS_INST/u_logic/Qflvx4 ,
         \CORTEXM0DS_INST/u_logic/Xflvx4 , \CORTEXM0DS_INST/u_logic/Eglvx4 ,
         \CORTEXM0DS_INST/u_logic/Lglvx4 , \CORTEXM0DS_INST/u_logic/Sglvx4 ,
         \CORTEXM0DS_INST/u_logic/Zglvx4 , \CORTEXM0DS_INST/u_logic/Ghlvx4 ,
         \CORTEXM0DS_INST/u_logic/Nhlvx4 , \CORTEXM0DS_INST/u_logic/Uhlvx4 ,
         \CORTEXM0DS_INST/u_logic/Bilvx4 , \CORTEXM0DS_INST/u_logic/Iilvx4 ,
         \CORTEXM0DS_INST/u_logic/Pilvx4 , \CORTEXM0DS_INST/u_logic/Wilvx4 ,
         \CORTEXM0DS_INST/u_logic/Djlvx4 , \CORTEXM0DS_INST/u_logic/Kjlvx4 ,
         \CORTEXM0DS_INST/u_logic/Rjlvx4 , \CORTEXM0DS_INST/u_logic/Yjlvx4 ,
         \CORTEXM0DS_INST/u_logic/Fklvx4 , \CORTEXM0DS_INST/u_logic/Mklvx4 ,
         \CORTEXM0DS_INST/u_logic/Tklvx4 , \CORTEXM0DS_INST/u_logic/Allvx4 ,
         \CORTEXM0DS_INST/u_logic/Hllvx4 , \CORTEXM0DS_INST/u_logic/Ollvx4 ,
         \CORTEXM0DS_INST/u_logic/Cmlvx4 , \CORTEXM0DS_INST/u_logic/Jmlvx4 ,
         \CORTEXM0DS_INST/u_logic/Qmlvx4 , \CORTEXM0DS_INST/u_logic/Xmlvx4 ,
         \CORTEXM0DS_INST/u_logic/Enlvx4 , \CORTEXM0DS_INST/u_logic/Lnlvx4 ,
         \CORTEXM0DS_INST/u_logic/Snlvx4 , \CORTEXM0DS_INST/u_logic/Znlvx4 ,
         \CORTEXM0DS_INST/u_logic/Golvx4 , \CORTEXM0DS_INST/u_logic/Nolvx4 ,
         \CORTEXM0DS_INST/u_logic/Uolvx4 , \CORTEXM0DS_INST/u_logic/Bplvx4 ,
         \CORTEXM0DS_INST/u_logic/Iplvx4 , \CORTEXM0DS_INST/u_logic/Pplvx4 ,
         \CORTEXM0DS_INST/u_logic/Wplvx4 , \CORTEXM0DS_INST/u_logic/Dqlvx4 ,
         \CORTEXM0DS_INST/u_logic/Kqlvx4 , \CORTEXM0DS_INST/u_logic/Rqlvx4 ,
         \CORTEXM0DS_INST/u_logic/Yqlvx4 , \CORTEXM0DS_INST/u_logic/Frlvx4 ,
         \CORTEXM0DS_INST/u_logic/Mrlvx4 , \CORTEXM0DS_INST/u_logic/Trlvx4 ,
         \CORTEXM0DS_INST/u_logic/Aslvx4 , \CORTEXM0DS_INST/u_logic/Hslvx4 ,
         \CORTEXM0DS_INST/u_logic/Oslvx4 , \CORTEXM0DS_INST/u_logic/Vslvx4 ,
         \CORTEXM0DS_INST/u_logic/Ctlvx4 , \CORTEXM0DS_INST/u_logic/Jtlvx4 ,
         \CORTEXM0DS_INST/u_logic/Qtlvx4 , \CORTEXM0DS_INST/u_logic/Xtlvx4 ,
         \CORTEXM0DS_INST/u_logic/Eulvx4 , \CORTEXM0DS_INST/u_logic/Lulvx4 ,
         \CORTEXM0DS_INST/u_logic/Sulvx4 , \CORTEXM0DS_INST/u_logic/Zulvx4 ,
         \CORTEXM0DS_INST/u_logic/Gvlvx4 , \CORTEXM0DS_INST/u_logic/Nvlvx4 ,
         \CORTEXM0DS_INST/u_logic/Uvlvx4 , \CORTEXM0DS_INST/u_logic/Bwlvx4 ,
         \CORTEXM0DS_INST/u_logic/Iwlvx4 , \CORTEXM0DS_INST/u_logic/Pwlvx4 ,
         \CORTEXM0DS_INST/u_logic/Wwlvx4 , \CORTEXM0DS_INST/u_logic/Dxlvx4 ,
         \CORTEXM0DS_INST/u_logic/Kxlvx4 , \CORTEXM0DS_INST/u_logic/Rxlvx4 ,
         \CORTEXM0DS_INST/u_logic/Yxlvx4 , \CORTEXM0DS_INST/u_logic/Fylvx4 ,
         \CORTEXM0DS_INST/u_logic/Mylvx4 , \CORTEXM0DS_INST/u_logic/Tylvx4 ,
         \CORTEXM0DS_INST/u_logic/Azlvx4 , \CORTEXM0DS_INST/u_logic/Hzlvx4 ,
         \CORTEXM0DS_INST/u_logic/Ozlvx4 , \CORTEXM0DS_INST/u_logic/Vzlvx4 ,
         \CORTEXM0DS_INST/u_logic/C0mvx4 , \CORTEXM0DS_INST/u_logic/J0mvx4 ,
         \CORTEXM0DS_INST/u_logic/Q0mvx4 , \CORTEXM0DS_INST/u_logic/X0mvx4 ,
         \CORTEXM0DS_INST/u_logic/E1mvx4 , \CORTEXM0DS_INST/u_logic/L1mvx4 ,
         \CORTEXM0DS_INST/u_logic/S1mvx4 , \CORTEXM0DS_INST/u_logic/Z1mvx4 ,
         \CORTEXM0DS_INST/u_logic/G2mvx4 , \CORTEXM0DS_INST/u_logic/N2mvx4 ,
         \CORTEXM0DS_INST/u_logic/U2mvx4 , \CORTEXM0DS_INST/u_logic/L8mvx4 ,
         \CORTEXM0DS_INST/u_logic/U9mvx4 , \CORTEXM0DS_INST/u_logic/Pamvx4 ,
         \CORTEXM0DS_INST/u_logic/Wamvx4 , \CORTEXM0DS_INST/u_logic/Jemvx4 ,
         \CORTEXM0DS_INST/u_logic/Qemvx4 , \CORTEXM0DS_INST/u_logic/Xemvx4 ,
         \CORTEXM0DS_INST/u_logic/Efmvx4 , \CORTEXM0DS_INST/u_logic/Lfmvx4 ,
         \CORTEXM0DS_INST/u_logic/Sfmvx4 , \CORTEXM0DS_INST/u_logic/Zfmvx4 ,
         \CORTEXM0DS_INST/u_logic/Ggmvx4 , \CORTEXM0DS_INST/u_logic/Ngmvx4 ,
         \CORTEXM0DS_INST/u_logic/Ugmvx4 , \CORTEXM0DS_INST/u_logic/Bhmvx4 ,
         \CORTEXM0DS_INST/u_logic/Ihmvx4 , \CORTEXM0DS_INST/u_logic/Phmvx4 ,
         \CORTEXM0DS_INST/u_logic/Whmvx4 , \CORTEXM0DS_INST/u_logic/Dimvx4 ,
         \CORTEXM0DS_INST/u_logic/Kimvx4 , \CORTEXM0DS_INST/u_logic/Rimvx4 ,
         \CORTEXM0DS_INST/u_logic/Yimvx4 , \CORTEXM0DS_INST/u_logic/Fjmvx4 ,
         \CORTEXM0DS_INST/u_logic/Mjmvx4 , \CORTEXM0DS_INST/u_logic/Tjmvx4 ,
         \CORTEXM0DS_INST/u_logic/Akmvx4 , \CORTEXM0DS_INST/u_logic/Hkmvx4 ,
         \CORTEXM0DS_INST/u_logic/Okmvx4 , \CORTEXM0DS_INST/u_logic/Vkmvx4 ,
         \CORTEXM0DS_INST/u_logic/Clmvx4 , \CORTEXM0DS_INST/u_logic/Jlmvx4 ,
         \CORTEXM0DS_INST/u_logic/Qlmvx4 , \CORTEXM0DS_INST/u_logic/Xlmvx4 ,
         \CORTEXM0DS_INST/u_logic/Emmvx4 , \CORTEXM0DS_INST/u_logic/Lmmvx4 ,
         \CORTEXM0DS_INST/u_logic/Smmvx4 , \CORTEXM0DS_INST/u_logic/F4nvx4 ,
         \CORTEXM0DS_INST/u_logic/G8nvx4 , \CORTEXM0DS_INST/u_logic/Acnvx4 ,
         \CORTEXM0DS_INST/u_logic/Ocnvx4 , \CORTEXM0DS_INST/u_logic/Jdnvx4 ,
         \CORTEXM0DS_INST/u_logic/Eenvx4 , \CORTEXM0DS_INST/u_logic/Lenvx4 ,
         \CORTEXM0DS_INST/u_logic/Senvx4 , \CORTEXM0DS_INST/u_logic/Zenvx4 ,
         \CORTEXM0DS_INST/u_logic/Gfnvx4 , \CORTEXM0DS_INST/u_logic/Ufnvx4 ,
         \CORTEXM0DS_INST/u_logic/Bgnvx4 , \CORTEXM0DS_INST/u_logic/Ignvx4 ,
         \CORTEXM0DS_INST/u_logic/S4qvx4 , \CORTEXM0DS_INST/u_logic/Wgnvx4 ,
         \CORTEXM0DS_INST/u_logic/Dhnvx4 , \CORTEXM0DS_INST/u_logic/V2qvx4 ,
         \CORTEXM0DS_INST/u_logic/Rhnvx4 , \CORTEXM0DS_INST/u_logic/Finvx4 ,
         \CORTEXM0DS_INST/u_logic/Minvx4 , \CORTEXM0DS_INST/u_logic/Tinvx4 ,
         \CORTEXM0DS_INST/u_logic/Ojnvx4 , \CORTEXM0DS_INST/u_logic/Y1pvx4 ,
         \CORTEXM0DS_INST/u_logic/Xxovx4 , \CORTEXM0DS_INST/u_logic/Jxovx4 ,
         \CORTEXM0DS_INST/u_logic/Owovx4 , \CORTEXM0DS_INST/u_logic/Fvovx4 ,
         \CORTEXM0DS_INST/u_logic/Yuovx4 , \CORTEXM0DS_INST/u_logic/Cqovx4 ,
         \CORTEXM0DS_INST/u_logic/Vpovx4 , \CORTEXM0DS_INST/u_logic/Rnovx4 ,
         \CORTEXM0DS_INST/u_logic/Ekovx4 , \CORTEXM0DS_INST/u_logic/Llnvx4 ,
         \CORTEXM0DS_INST/u_logic/Slnvx4 , \CORTEXM0DS_INST/u_logic/Z6ovx4 ,
         \CORTEXM0DS_INST/u_logic/Pxdvx4 , \CORTEXM0DS_INST/u_logic/H0gvx4 ,
         \CORTEXM0DS_INST/u_logic/W1evx4 , \CORTEXM0DS_INST/u_logic/Itdvx4 ,
         \CORTEXM0DS_INST/u_logic/Mqdvx4 , \CORTEXM0DS_INST/u_logic/Rddvx4 ,
         \CORTEXM0DS_INST/u_logic/Gcdvx4 , \CORTEXM0DS_INST/u_logic/Oy8vx4 ,
         \CORTEXM0DS_INST/u_logic/Fs8vx4 , \CORTEXM0DS_INST/u_logic/Vu8vx4 ,
         \CORTEXM0DS_INST/u_logic/Y3dvx4 , \CORTEXM0DS_INST/u_logic/S0hvx4 ,
         \CORTEXM0DS_INST/u_logic/F2hvx4 , \CORTEXM0DS_INST/u_logic/N6hvx4 ,
         \CORTEXM0DS_INST/u_logic/O2dvx4 , \CORTEXM0DS_INST/u_logic/E1dvx4 ,
         \CORTEXM0DS_INST/u_logic/Ukdvx4 , \CORTEXM0DS_INST/u_logic/C8dvx4 ,
         \CORTEXM0DS_INST/u_logic/S6dvx4 , \CORTEXM0DS_INST/u_logic/Nt8vx4 ,
         \CORTEXM0DS_INST/u_logic/Ks9vx4 , \CORTEXM0DS_INST/u_logic/Gr9vx4 ,
         \CORTEXM0DS_INST/u_logic/Cq9vx4 , \CORTEXM0DS_INST/u_logic/Uzcvx4 ,
         \CORTEXM0DS_INST/u_logic/Bx9vx4 , \CORTEXM0DS_INST/u_logic/Wv9vx4 ,
         \CORTEXM0DS_INST/u_logic/Cf9vx4 , \CORTEXM0DS_INST/u_logic/Ud9vx4 ,
         \CORTEXM0DS_INST/u_logic/Mc9vx4 , \CORTEXM0DS_INST/u_logic/Fb9vx4 ,
         \CORTEXM0DS_INST/u_logic/Y99vx4 , \CORTEXM0DS_INST/u_logic/R89vx4 ,
         \CORTEXM0DS_INST/u_logic/K79vx4 , \CORTEXM0DS_INST/u_logic/D69vx4 ,
         \CORTEXM0DS_INST/u_logic/W49vx4 , \CORTEXM0DS_INST/u_logic/P39vx4 ,
         \CORTEXM0DS_INST/u_logic/I29vx4 , \CORTEXM0DS_INST/u_logic/V8evx4 ,
         \CORTEXM0DS_INST/u_logic/G8fvx4 , \CORTEXM0DS_INST/u_logic/V6fvx4 ,
         \CORTEXM0DS_INST/u_logic/Z3fvx4 , \CORTEXM0DS_INST/u_logic/O2fvx4 ,
         \CORTEXM0DS_INST/u_logic/D1fvx4 , \CORTEXM0DS_INST/u_logic/Tzevx4 ,
         \CORTEXM0DS_INST/u_logic/Jyevx4 , \CORTEXM0DS_INST/u_logic/Zwevx4 ,
         \CORTEXM0DS_INST/u_logic/Pvevx4 , \CORTEXM0DS_INST/u_logic/R9fvx4 ,
         \CORTEXM0DS_INST/u_logic/Fuevx4 , \CORTEXM0DS_INST/u_logic/I4gvx4 ,
         \CORTEXM0DS_INST/u_logic/A3gvx4 , \CORTEXM0DS_INST/u_logic/Mk8vx4 ,
         \CORTEXM0DS_INST/u_logic/Aj9vx4 , \CORTEXM0DS_INST/u_logic/Bwfvx4 ,
         \CORTEXM0DS_INST/u_logic/Qufvx4 , \CORTEXM0DS_INST/u_logic/Ftfvx4 ,
         \CORTEXM0DS_INST/u_logic/Urfvx4 , \CORTEXM0DS_INST/u_logic/Jqfvx4 ,
         \CORTEXM0DS_INST/u_logic/Yofvx4 , \CORTEXM0DS_INST/u_logic/Onfvx4 ,
         \CORTEXM0DS_INST/u_logic/Emfvx4 , \CORTEXM0DS_INST/u_logic/Ukfvx4 ,
         \CORTEXM0DS_INST/u_logic/Kjfvx4 , \CORTEXM0DS_INST/u_logic/Aifvx4 ,
         \CORTEXM0DS_INST/u_logic/Qgfvx4 , \CORTEXM0DS_INST/u_logic/Gffvx4 ,
         \CORTEXM0DS_INST/u_logic/Wdfvx4 , \CORTEXM0DS_INST/u_logic/Mcfvx4 ,
         \CORTEXM0DS_INST/u_logic/Cbfvx4 , \CORTEXM0DS_INST/u_logic/Mxfvx4 ,
         \CORTEXM0DS_INST/u_logic/Xyfvx4 , \CORTEXM0DS_INST/u_logic/Ki8vx4 ,
         \CORTEXM0DS_INST/u_logic/Krgvx4 , \CORTEXM0DS_INST/u_logic/Ul8vx4 ,
         \CORTEXM0DS_INST/u_logic/Rkgvx4 , \CORTEXM0DS_INST/u_logic/Wtgvx4 ,
         \CORTEXM0DS_INST/u_logic/Hx8vx4 , \CORTEXM0DS_INST/u_logic/Vogvx4 ,
         \CORTEXM0DS_INST/u_logic/Nngvx4 , \CORTEXM0DS_INST/u_logic/Pp8vx4 ,
         \CORTEXM0DS_INST/u_logic/Mj8vx4 , \CORTEXM0DS_INST/u_logic/Q5gvx4 ,
         \CORTEXM0DS_INST/u_logic/Fjgvx4 , \CORTEXM0DS_INST/u_logic/Dmgvx4 ,
         \CORTEXM0DS_INST/u_logic/Ot9vx4 , \CORTEXM0DS_INST/u_logic/Eg8vx4 ,
         \CORTEXM0DS_INST/u_logic/Z7hvx4 , \CORTEXM0DS_INST/u_logic/Wadvx4 ,
         \CORTEXM0DS_INST/u_logic/M9dvx4 , \CORTEXM0DS_INST/u_logic/Ngdvx4 ,
         \CORTEXM0DS_INST/u_logic/Cfdvx4 , \CORTEXM0DS_INST/u_logic/Ik9vx4 ,
         \CORTEXM0DS_INST/u_logic/Yo9vx4 , \CORTEXM0DS_INST/u_logic/Vsevx4 ,
         \CORTEXM0DS_INST/u_logic/Xrdvx4 , \CORTEXM0DS_INST/u_logic/Jjdvx4 ,
         \CORTEXM0DS_INST/u_logic/Yhdvx4 , \CORTEXM0DS_INST/u_logic/Kycvx4 ,
         \CORTEXM0DS_INST/u_logic/Un9vx4 , \CORTEXM0DS_INST/u_logic/Lrevx4 ,
         \CORTEXM0DS_INST/u_logic/L9hvx4 , \CORTEXM0DS_INST/u_logic/I5dvx4 ,
         \CORTEXM0DS_INST/u_logic/Bpdvx4 , \CORTEXM0DS_INST/u_logic/Qndvx4 ,
         \CORTEXM0DS_INST/u_logic/Fmdvx4 , \CORTEXM0DS_INST/u_logic/H3evx4 ,
         \CORTEXM0DS_INST/u_logic/Izgvx4 , \CORTEXM0DS_INST/u_logic/Qm9vx4 ,
         \CORTEXM0DS_INST/u_logic/Bqevx4 , \CORTEXM0DS_INST/u_logic/Kg9vx4 ,
         \CORTEXM0DS_INST/u_logic/K5fvx4 , \CORTEXM0DS_INST/u_logic/Xlevx4 ,
         \CORTEXM0DS_INST/u_logic/Ml9vx4 , \CORTEXM0DS_INST/u_logic/B19vx4 ,
         \CORTEXM0DS_INST/u_logic/Roevx4 , \CORTEXM0DS_INST/u_logic/B5hvx4 ,
         \CORTEXM0DS_INST/u_logic/Mf8vx4 , \CORTEXM0DS_INST/u_logic/D6evx4 ,
         \CORTEXM0DS_INST/u_logic/Xq8vx4 , \CORTEXM0DS_INST/u_logic/Su9vx4 ,
         \CORTEXM0DS_INST/u_logic/Vdgvx4 , \CORTEXM0DS_INST/u_logic/Z6gvx4 ,
         \CORTEXM0DS_INST/u_logic/U9gvx4 , \CORTEXM0DS_INST/u_logic/Dbgvx4 ,
         \CORTEXM0DS_INST/u_logic/Qsgvx4 , \CORTEXM0DS_INST/u_logic/L0evx4 ,
         \CORTEXM0DS_INST/u_logic/Azdvx4 , \CORTEXM0DS_INST/u_logic/R3hvx4 ,
         \CORTEXM0DS_INST/u_logic/Mcgvx4 , \CORTEXM0DS_INST/u_logic/Efgvx4 ,
         \CORTEXM0DS_INST/u_logic/Nggvx4 , \CORTEXM0DS_INST/u_logic/Ho8vx4 ,
         \CORTEXM0DS_INST/u_logic/Ewdvx4 , \CORTEXM0DS_INST/u_logic/Tudvx4 ,
         \CORTEXM0DS_INST/u_logic/O7evx4 , \CORTEXM0DS_INST/u_logic/Uz8vx4 ,
         \CORTEXM0DS_INST/u_logic/Hnevx4 , \CORTEXM0DS_INST/u_logic/Eqgvx4 ,
         \CORTEXM0DS_INST/u_logic/Whgvx4 , \CORTEXM0DS_INST/u_logic/Cn8vx4 ,
         \CORTEXM0DS_INST/u_logic/Ih8vx4 , \CORTEXM0DS_INST/u_logic/S4evx4 ,
         \CORTEXM0DS_INST/u_logic/O8gvx4 , \CORTEXM0DS_INST/u_logic/Dw8vx4 ,
         \CORTEXM0DS_INST/u_logic/Sh9vx4 , \CORTEXM0DS_INST/u_logic/Xahvx4 ,
         n1, n2, n450, n488, n489, n1061, n1062, n1063, n1076, n1079, n1081,
         n1084, n1086, n1089, n1091, n1094, n1096, n1101, n1104, n1106, n1109,
         n1111, n1114, n1116, n1119, n1121, n1124, n1126, n1129, n1131, n1134,
         n1136, n1139, n1141, n1144, n1145, n1147, n1148, n1154, n1155, n1157,
         n1160, n1162, n1164, n1166, n1168, n1169, n1172, n1174, n1176, n1178,
         n1180, n1182, n1184, n1186, n1188, n1403, n1473, n1476, n1479, n1482,
         n1485, n1488, n1491, n1495, n1497, n1501, n1505, n1506, n1510, n1515,
         n1521, n1629, n1630, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1670, n1671, n1672, n1675, n1676, n1677, n1678, n1685, n1687, n1691,
         n1709, n1744, n1770, n1789, n1813, n1851, n1870, n1944, n2057, n2060,
         n2065, n2069, n2095, n2120, n2122, n2135, n2136, n2140, n2168, n2197,
         n2198, n2205, n2208, n2209, n2212, n2213, n2214, n2215, n2216, n2217,
         n2266, n2267, n2270, n2271, n2326, n2328, n2460, n2463, n2464, n2490,
         n2492, n2500, n2502, n2511, n2512, n2513, n2514, n2528, n2531, n2533,
         n2541, n2543, n2544, n2577, n2620, n2623, n2624, n2626, n2627, n2641,
         n2644, n2645, n2647, n2648, n2683, n2686, n2711, n2713, n2714, n2754,
         n2757, n2774, n2776, n2786, n2790, n2791, n2976, n2984, n3002, n3015,
         n3016, n3024, n3025, n3027, n3048, n3049, n3067, n3081, n3082, n3084,
         n3101, n3127, n3128, n3164, n3178, n3197, n3204, n3217, n3223, n3224,
         n3226, n3227, n3228, n3229, n3230, n3231, n3233, n3317, n3348, n3368,
         n3392, n3419, n3485, n3514, n3554, n3958, n3962, n3977, n3978, n3979,
         n4087, n4092, n4097, n4109, n4110, n4130, n4150, n4175, n4180, n4185,
         n4190, n4203, n4227, n4237, n4241, n4243, n4263, n4348, n4408, n4585,
         n4626, n4627, n4704, n4706, n4708, n4711, n4712, n4814, n4815, n4816,
         n4831, n5021, n5022, n5100, n5428, n5664, n5780, n5822, n5888, n5889,
         n5893, n5894, n5914, n5915, n5916, n5920, n5921, n5924, n5926, n5928,
         n5931, n5932, n5933, n5935, n5937, n5938, n5939, n5940, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6147, n6149, n6153,
         n6156, n6157, n6159, n6162, n6163, n6164, n6166, n6167, n6171, n6172,
         n6173, n6175, n6176, n6177, n6180, n6181, n6182, n6183, n6189, n6190,
         n6192, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751;
  wire   [31:0] PID_haddr_top;
  wire   [3:0] PID_hprot_top;
  wire   [2:0] PID_hsize_top;
  wire   [31:0] PID_hwdata_top;
  wire   [31:0] RAM_hrdata_top;
  wire   [2:0] \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state ;
  wire   [2:0] \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_nextstate ;
  wire   [4:1] \interconnect_ip_inst/i_ahb_U_mux_hsel_prev ;
  wire   [5:0] \CORTEXM0DS_INST/vis_ipsr ;
  wire   [3:0] \CORTEXM0DS_INST/vis_apsr ;
  wire   [30:0] \CORTEXM0DS_INST/vis_pc ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r14 ;
  wire   [29:0] \CORTEXM0DS_INST/vis_psp ;
  wire   [29:0] \CORTEXM0DS_INST/vis_msp ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r12 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r11 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r10 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r09 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r08 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r07 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r06 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r05 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r04 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r03 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r02 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r01 ;
  wire   [31:0] \CORTEXM0DS_INST/cm0_r00 ;
  wire   [15:0] \CORTEXM0DS_INST/u_logic/L0i2z4 ;
  wire   [1:0] \CORTEXM0DS_INST/u_logic/Uth2z4 ;
  wire   [1:0] \CORTEXM0DS_INST/u_logic/Zph2z4 ;
  wire   [1:0] \CORTEXM0DS_INST/u_logic/Txh2z4 ;
  wire   [23:0] \CORTEXM0DS_INST/u_logic/Irh2z4 ;
  wire   [23:0] \CORTEXM0DS_INST/u_logic/Czh2z4 ;
  wire   [31:0] \CORTEXM0DS_INST/u_logic/Zuh2z4 ;
  wire   [15:0] \CORTEXM0DS_INST/u_logic/T1i2z4 ;
  wire   [1:0] \CORTEXM0DS_INST/u_logic/Psh2z4 ;
  wire   [3:0] \CORTEXM0DS_INST/u_logic/Tjh2z4 ;
  wire   UNCONNECTED_0;

  CPU_stub CPU_stub_inst ( .i_ssi_rxd(), .i_ssi_ss_in_n(), .i_ssi_ssi_clk(
        i_ssi_ssi_clk_top), .i_ssi_ssi_rst_n(i_ssi_ssi_rst_n_top), 
        .i_ssi_sclk_out(i_ssi_sclk_out_top), .i_ssi_ss_0_n(i_ssi_ss_0_n_top), 
        .i_ssi_ssi_mst_intr_n(i_ssi_ssi_mst_intr_n_top), .i_ssi_ssi_oe_n(
        i_ssi_ssi_oe_n_top), .i_ssi_ssi_rxf_intr_n(i_ssi_ssi_rxf_intr_n_top), 
        .i_ssi_ssi_rxo_intr_n(i_ssi_ssi_rxo_intr_n_top), 
        .i_ssi_ssi_rxu_intr_n(i_ssi_ssi_rxu_intr_n_top), .i_ssi_ssi_sleep(
        i_ssi_ssi_sleep_top), .i_ssi_ssi_txe_intr_n(i_ssi_ssi_txe_intr_n_top), 
        .i_ssi_ssi_txo_intr_n(i_ssi_ssi_intr_n_top), .i_ssi_txd(i_ssi_txd_top), 
        .HCLK(HCLK_top), .HRESETn(HRESETn_top) );
  cortexM0RAM ram2ahb_wrapper_inst ( .HCLK(HCLK_top), .HRESETn(HRESETn_top), 
        .ex_i_ahb_AHB_Slave_RAM_hrdata(RAM_hrdata_top), 
        .ex_i_ahb_AHB_Slave_RAM_hready_resp(RAM_hready_resp_top), 
        .ex_i_ahb_AHB_Slave_RAM_hresp({UNCONNECTED_0, \RAM_hresp_top[0] }), 
        .ex_i_ahb_AHB_Slave_RAM_haddr(PID_haddr_top), 
        .ex_i_ahb_AHB_Slave_RAM_hburst({1'b0, 1'b0, 1'b0}), 
        .ex_i_ahb_AHB_Slave_RAM_hmastlock(PID_hmastlock_top), 
        .ex_i_ahb_AHB_Slave_RAM_hprot({PID_hprot_top[3:2], 1'b1, 
        PID_hprot_top[0]}), .ex_i_ahb_AHB_Slave_RAM_hready(HREADY_top), 
        .ex_i_ahb_AHB_Slave_RAM_hsel(RAM_hsel_top), 
        .ex_i_ahb_AHB_Slave_RAM_hsize({1'b0, PID_hsize_top[1:0]}), 
        .ex_i_ahb_AHB_Slave_RAM_htrans({\PID_htrans_top[1] , 1'b0}), 
        .ex_i_ahb_AHB_Slave_RAM_hwdata(PID_hwdata_top), 
        .ex_i_ahb_AHB_Slave_RAM_hwrite(PID_hwrite_top) );
  nand2_1 \interconnect_ip_inst/U11942  ( .ip1(1'b0), .ip2(1'b1), .op(
        i_ssi_ssi_rxf_intr_n_top) );
  nand2_1 \interconnect_ip_inst/U11875  ( .ip1(1'b0), .ip2(1'b1), .op(
        i_ssi_ssi_txe_intr_n_top) );
  nand2_1 \interconnect_ip_inst/U11802  ( .ip1(1'b0), .ip2(1'b1), .op(
        i_ssi_ssi_rxo_intr_n_top) );
  nand2_1 \interconnect_ip_inst/U11791  ( .ip1(1'b0), .ip2(1'b1), .op(
        i_ssi_ssi_intr_n_top) );
  nand2_1 \interconnect_ip_inst/U11778  ( .ip1(1'b0), .ip2(1'b1), .op(
        i_ssi_ssi_rxu_intr_n_top) );
  nand2_1 \interconnect_ip_inst/U10788  ( .ip1(1'b0), .ip2(1'b1), .op(
        i_ssi_ssi_mst_intr_n_top) );
  nor2_1 \interconnect_ip_inst/U7231  ( .ip1(PID_haddr_top[17]), .ip2(n6117), 
        .op(RAM_hsel_top) );
  inv_1 \interconnect_ip_inst/U6038  ( .ip(1'b0), .op(i_ssi_ss_0_n_top) );
  nand2_1 \interconnect_ip_inst/U5634  ( .ip1(\interconnect_ip_inst/n6491 ), 
        .ip2(\interconnect_ip_inst/n5991 ), .op(HREADY_top) );
  drsp_1 \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_hready_resp_reg  ( .ip(
        \interconnect_ip_inst/n4829 ), .ck(HCLK_top), .rb(1'b1), .s(n12696), 
        .q(\interconnect_ip_inst/i_apb_hready_resp ) );
  drp_1 \interconnect_ip_inst/i_ssi_U_regfile_ssi_sleep_ir_reg  ( .ip(
        \interconnect_ip_inst/i_ssi_fsm_sleep ), .ck(HCLK_top), .rb(
        HRESETn_top), .q(i_ssi_ssi_sleep_top) );
  drp_1 \interconnect_ip_inst/i_ssi_U_mstfsm_fsm_sleep_reg  ( .ip(
        \interconnect_ip_inst/i_ssi_U_mstfsm_c_state[3] ), .ck(
        i_ssi_ssi_clk_top), .rb(i_ssi_ssi_rst_n_top), .q(
        \interconnect_ip_inst/i_ssi_fsm_sleep ) );
  drp_1 \interconnect_ip_inst/i_ssi_U_sclkgen_sclk_out_reg  ( .ip(1'b0), .ck(
        i_ssi_ssi_clk_top), .rb(i_ssi_ssi_rst_n_top), .q(i_ssi_sclk_out_top)
         );
  drp_1 \interconnect_ip_inst/i_ssi_U_shift_U_tx_shifter_txd_reg  ( .ip(
        i_ssi_txd_top), .ck(i_ssi_ssi_clk_top), .rb(i_ssi_ssi_rst_n_top), .q(
        i_ssi_txd_top) );
  drp_1 \interconnect_ip_inst/i_ssi_U_mstfsm_c_state_reg_3_  ( .ip(1'b1), .ck(
        i_ssi_ssi_clk_top), .rb(i_ssi_ssi_rst_n_top), .q(
        \interconnect_ip_inst/i_ssi_U_mstfsm_c_state[3] ) );
  drp_1 \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state_reg_2_  ( .ip(
        \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_nextstate [2]), .ck(
        HCLK_top), .rb(HRESETn_top), .q(
        \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state [2]) );
  drp_1 \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state_reg_0_  ( .ip(
        \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_nextstate [0]), .ck(
        HCLK_top), .rb(HRESETn_top), .q(
        \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state [0]) );
  drp_1 \interconnect_ip_inst/i_ahb_U_arblite_hmastlock_reg  ( .ip(
        \interconnect_ip_inst/n4860 ), .ck(HCLK_top), .rb(HRESETn_top), .q(
        PID_hmastlock_top) );
  drp_1 \interconnect_ip_inst/i_ahb_U_mux_hsel_prev_reg_1_  ( .ip(
        \interconnect_ip_inst/n4861 ), .ck(HCLK_top), .rb(HRESETn_top), .q(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [1]) );
  drp_1 \interconnect_ip_inst/i_ahb_U_mux_hsel_prev_reg_2_  ( .ip(
        \interconnect_ip_inst/n4862 ), .ck(HCLK_top), .rb(HRESETn_top), .q(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [2]) );
  drp_1 \interconnect_ip_inst/i_ahb_U_mux_hsel_prev_reg_3_  ( .ip(
        \interconnect_ip_inst/n4863 ), .ck(HCLK_top), .rb(HRESETn_top), .q(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [3]) );
  drp_1 \interconnect_ip_inst/i_ahb_U_mux_hsel_prev_reg_4_  ( .ip(
        \interconnect_ip_inst/n4864 ), .ck(HCLK_top), .rb(HRESETn_top), .q(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [4]) );
  drp_1 \interconnect_ip_inst/i_ahb_U_dfltslv_hresp_none_reg_0_  ( .ip(
        \interconnect_ip_inst/i_ahb_U_dfltslv_N4 ), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\interconnect_ip_inst/i_ahb_hresp_none_0_ ) );
  drp_1 \interconnect_ip_inst/i_ahb_U_dfltslv_current_state_reg  ( .ip(
        \interconnect_ip_inst/n10765 ), .ck(HCLK_top), .rb(HRESETn_top), .q(
        \interconnect_ip_inst/i_ahb_U_dfltslv_current_state ) );
  drsp_1 \interconnect_ip_inst/i_ssi_U_mstfsm_ssi_oe_n_reg  ( .ip(1'b1), .ck(
        i_ssi_ssi_clk_top), .rb(1'b1), .s(\interconnect_ip_inst/n11572 ), .q(
        i_ssi_ssi_oe_n_top) );
  drp_1 \CORTEXM0DS_INST/u_logic/J6i2z4_reg  ( .ip(n6067), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Xahvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/A4t2z4_reg  ( .ip(n6015), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Dmgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Pet2z4_reg  ( .ip(n6007), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Hx8vx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Mjl2z4_reg  ( .ip(n6066), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/B5hvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Jhy2z4_reg  ( .ip(n6048), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/V8evx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Emi2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qxhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Whgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Uqi2z4_reg  ( .ip(n6011), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Psh2z4 [1]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Zei2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Finvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/vis_apsr [1]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Gji2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/H3ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Ih8vx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Tki2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xxhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Cn8vx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Hzj2z4_reg  ( .ip(n6119), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/R3hvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Y6t2z4_reg  ( .ip(n6009), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Q5gvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/I6w2z4_reg  ( .ip(n6071), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Ul8vx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Qrp2z4_reg  ( .ip(n6013), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Txh2z4 [1]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Kop2z4_reg  ( .ip(n6068), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L9hvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/P2a3z4_reg  ( .ip(n6014), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Uth2z4 [1]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Vve3z4_reg  ( .ip(n6157), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [9]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Wbk2z4_reg  ( .ip(n6149), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Qsgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/S4w2z4_reg  ( .ip(n6008), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Rkgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/U7w2z4_reg  ( .ip(n6164), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Krgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Fed3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Efmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [4]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Nnc3z4_reg  ( .ip(n6162), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [10]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ble3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uzhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [11]) );
  drp_1 \CORTEXM0DS_INST/u_logic/D4g3z4_reg  ( .ip(n6153), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [13]) );
  drp_1 \CORTEXM0DS_INST/u_logic/T8f3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/P0ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [8]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Sgj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Owhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Efgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Vaw2z4_reg  ( .ip(n6065), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Xyfvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ffj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vwhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Nggvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Aok2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mvhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Dbgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Fij2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hwhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Mcgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/L8t2z4_reg  ( .ip(n6114), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Mj8vx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ark2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yuhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Z6gvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Nsk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ruhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Vdgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Nbm2z4_reg  ( .ip(n6115), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Xlevx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Cam2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/L8mvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/vis_ipsr [3]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Trq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pamvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/vis_ipsr [4]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Tdp2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wamvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/vis_ipsr [5]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Npk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fvhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/U9gvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Y9t2z4_reg  ( .ip(n6006), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Pp8vx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Thm2z4_reg  ( .ip(n6064), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/cm0_primask[0] ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Wxp2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/X9kvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zph2z4 [1]) );
  drp_1 \CORTEXM0DS_INST/u_logic/C3w2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ufnvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zph2z4 [0]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Dpc3z4_reg  ( .ip(n6177), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [12]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ffs2z4_reg  ( .ip(n6069), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Z7hvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/U5x2z4_reg  ( .ip(n6072), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Mk8vx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Uaj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/U9mvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/vis_ipsr [2]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Uyv2z4_reg  ( .ip(n6163), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Wtgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Nen2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ollvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/cm0_control[1] ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Idk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rhnvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/vis_apsr [0]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Lz93z4_reg  ( .ip(n6070), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/N6hvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ywi2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Owgvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Eqgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/K3l2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/F4nvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Mf8vx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Cps2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vkmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [31]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Uls2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jlmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [29]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Dks2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qlmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [28]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Tib3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lmmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [25]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Pab3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Smmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [24]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Azs2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rimvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [23]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Svs2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fjmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [21]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Bus2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mjmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [20]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Kkb3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hkmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [17]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Gcb3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Okmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [16]) );
  drp_1 \CORTEXM0DS_INST/u_logic/H8l2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ngmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [15]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Z4l2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bhmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [13]) );
  drp_1 \CORTEXM0DS_INST/u_logic/G8n2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ihmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [12]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Bmb3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dimvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [9]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Xdb3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kimvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [8]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Bjd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jemvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [7]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Vfd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xemvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [5]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Zad3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zfmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [1]) );
  drp_1 \CORTEXM0DS_INST/u_logic/J9d3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ggmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [0]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Gxk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/T2ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [0]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Vac3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/M2ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [1]) );
  drp_1 \CORTEXM0DS_INST/u_logic/F4c3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/D1ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [6]) );
  drp_1 \CORTEXM0DS_INST/u_logic/N7c3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/K1ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [5]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Oar2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nzhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [12]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ipb3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/R1ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [4]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Hub3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Y1ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [3]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Pxb3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/F2ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [2]) );
  drp_1 \CORTEXM0DS_INST/u_logic/X0c3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/W0ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [7]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ipn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/B0ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [10]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Y9l2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/I0ivx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [9]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Wuq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gzhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [13]) );
  drp_1 \CORTEXM0DS_INST/u_logic/V3o2z4_reg  ( .ip(n6145), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Izgvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ztc3z4_reg  ( .ip(n6192), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [0]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Mcc3z4_reg  ( .ip(n6189), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [1]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Jkc3z4_reg  ( .ip(n6182), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [6]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Uic3z4_reg  ( .ip(n6180), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [5]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Fhc3z4_reg  ( .ip(n6175), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [4]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Qfc3z4_reg  ( .ip(n6173), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [3]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Bec3z4_reg  ( .ip(n6171), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [2]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ylc3z4_reg  ( .ip(n6166), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [7]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Lee3z4_reg  ( .ip(n6159), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [11]) );
  drp_1 \CORTEXM0DS_INST/u_logic/H2f3z4_reg  ( .ip(n6156), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [8]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Lns2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Clmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [30]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Jxs2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yimvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [22]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Q6l2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ugmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [14]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Lhd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qemvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [6]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Mis2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Emmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [26]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Kss2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Akmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [18]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Axm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Whmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [10]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Pcd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sfmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [2]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Tqc3z4_reg  ( .ip(n6183), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [14]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Rym2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zyhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [14]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Vgs2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xlmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [27]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Tqs2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tjmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [19]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Usl2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Phmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [11]) );
  drp_1 \CORTEXM0DS_INST/u_logic/T7d3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lfmvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/Zuh2z4 [3]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Lul2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Syhvx4 ), .ck(HCLK_top), .rb(HRESETn_top), 
        .q(\CORTEXM0DS_INST/u_logic/T1i2z4 [15]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Jsc3z4_reg  ( .ip(n6147), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/L0i2z4 [15]) );
  drp_1 \CORTEXM0DS_INST/u_logic/Ypi3z4_reg  ( .ip(n6118), .ck(HCLK_top), .rb(
        HRESETn_top), .q(SYSRESETREQ_top_out) );
  drp_1 \CORTEXM0DS_INST/u_logic/Aqp2z4_reg  ( .ip(n5975), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Txh2z4 [0]) );
  drp_1 \CORTEXM0DS_INST/u_logic/B1a3z4_reg  ( .ip(n5974), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Uth2z4 [0]) );
  drp_1 \CORTEXM0DS_INST/u_logic/X9n2z4_reg  ( .ip(n5973), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Psh2z4 [0]) );
  drp_1 \CORTEXM0DS_INST/u_logic/R0t2z4_reg  ( .ip(n5972), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Eg8vx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Mbt2z4_reg  ( .ip(n5971), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Nngvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Adt2z4_reg  ( .ip(n5970), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/Vogvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/Tna3z4_reg  ( .ip(n5969), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/F2hvx4 ) );
  drp_1 \CORTEXM0DS_INST/u_logic/S5b3z4_reg  ( .ip(n5968), .ck(HCLK_top), .rb(
        HRESETn_top), .q(\CORTEXM0DS_INST/u_logic/S0hvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/H9i2z4_reg  ( .ip(n6016), .ck(HCLK_top), 
        .rb(1'b1), .s(\CORTEXM0DS_INST/u_logic/N586 ), .q(
        \CORTEXM0DS_INST/u_logic/Sh9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hxx2z4_reg  ( .ip(n6010), .ck(HCLK_top), 
        .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/u_logic/A3gvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tyx2z4_reg  ( .ip(n6110), .ck(HCLK_top), 
        .rb(1'b1), .s(\CORTEXM0DS_INST/u_logic/N586 ), .q(
        \CORTEXM0DS_INST/u_logic/I4gvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hyy2z4_reg  ( .ip(n6017), .ck(HCLK_top), 
        .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/u_logic/Cf9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I2t2z4_reg  ( .ip(n6073), .ck(HCLK_top), 
        .rb(1'b1), .s(\CORTEXM0DS_INST/u_logic/N586 ), .q(
        \CORTEXM0DS_INST/u_logic/Ot9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cqo2z4_reg  ( .ip(n6078), .ck(HCLK_top), 
        .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/u_logic/H3evx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Igi2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cflvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/vis_apsr [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rhi2z4_reg  ( .ip(n6084), .ck(HCLK_top), 
        .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/u_logic/S4evx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ft73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xflvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/cm0_r02 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Iwp2z4_reg  ( .ip(n6082), .ck(HCLK_top), 
        .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/u_logic/Kycvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U4z2z4_reg  ( .ip(n6083), .ck(HCLK_top), 
        .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/u_logic/Uzcvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/S3i3z4_reg  ( .ip(n6127), .ck(HCLK_top), 
        .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bdm2z4_reg  ( .ip(n6050), .ck(HCLK_top), 
        .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/u_logic/K5fvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fcj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cxhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/vis_pc [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Swy2z4_reg  ( .ip(n6018), .ck(HCLK_top), 
        .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/u_logic/Ud9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cyq2z4_reg  ( .ip(n6111), .ck(HCLK_top), 
        .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/u_logic/Yo9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Svk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kuhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/u_logic/Xq8vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gci2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/V3ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/vis_apsr [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/V1l2z4_reg  ( .ip(n6108), .ck(HCLK_top), 
        .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/u_logic/D6evx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pdi2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Eyhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/u_logic/O8gvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/C183z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Atkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r02 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Q7j2z4_reg  ( .ip(n6077), .ck(HCLK_top), 
        .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/u_logic/Ewdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ogo2z4_reg  ( .ip(n6123), .ck(HCLK_top), 
        .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F483z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wjkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/cm0_r02 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jca3z4_reg  ( .ip(n6012), .ck(HCLK_top), 
        .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z7i2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ojnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_xpsr[24] ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/T1y2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Slnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/R9fvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jcw2z4_reg  ( .ip(n6005), .ck(HCLK_top), 
        .rb(1'b1), .s(n12739), .q(\CORTEXM0DS_INST/u_logic/Mxfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qdj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Llnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12738), .q(\CORTEXM0DS_INST/u_logic/Ho8vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Auk2z4_reg  ( .ip(n6075), .ck(HCLK_top), 
        .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/u_logic/Su9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yaz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pfhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12737), .q(\CORTEXM0DS_INST/u_logic/Nt8vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wbf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/C4ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r00 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/G6d3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sqivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/Oy8vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/G1s2z4_reg  ( .ip(n6104), .ck(HCLK_top), 
        .rb(1'b1), .s(n12739), .q(\CORTEXM0DS_INST/u_logic/Wadvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kyi2z4_reg  ( .ip(n6063), .ck(HCLK_top), 
        .rb(1'b1), .s(n12739), .q(\CORTEXM0DS_INST/u_logic/Hnevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yzi2z4_reg  ( .ip(n6029), .ck(HCLK_top), 
        .rb(1'b1), .s(n12739), .q(\CORTEXM0DS_INST/u_logic/Uz8vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dq73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/E1mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12739), .q(\CORTEXM0DS_INST/cm0_r02 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/An73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/S1mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12739), .q(\CORTEXM0DS_INST/cm0_r02 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ohh3z4_reg  ( .ip(n6079), .ck(HCLK_top), 
        .rb(1'b1), .s(n12739), .q(\CORTEXM0DS_INST/u_logic/W1evx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/T583z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hfkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12739), .q(\CORTEXM0DS_INST/cm0_r02 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z2h3z4_reg  ( .ip(n6124), .ck(HCLK_top), 
        .rb(1'b1), .s(n12739), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rdg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Swjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12739), .q(\CORTEXM0DS_INST/cm0_r02 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tzg3z4_reg  ( .ip(n6094), .ck(HCLK_top), 
        .rb(1'b1), .s(n12739), .q(\CORTEXM0DS_INST/u_logic/Mqdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Llq2z4_reg  ( .ip(n6093), .ck(HCLK_top), 
        .rb(1'b1), .s(n12739), .q(\CORTEXM0DS_INST/u_logic/Xrdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ka83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/H1kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12739), .q(\CORTEXM0DS_INST/cm0_r02 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/G0w2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Acnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12738), .q(\CORTEXM0DS_INST/vis_ipsr [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/G9w2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lrhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12738), .q(\CORTEXM0DS_INST/u_logic/Ki8vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/H3d3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/G2mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12738), .q(\CORTEXM0DS_INST/u_logic/Fs8vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lbn2z4_reg  ( .ip(n6061), .ck(HCLK_top), 
        .rb(1'b1), .s(n12738), .q(\CORTEXM0DS_INST/u_logic/Bqevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Viy2z4_reg  ( .ip(n6027), .ck(HCLK_top), 
        .rb(1'b1), .s(n12738), .q(\CORTEXM0DS_INST/u_logic/I29vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/K1z2z4_reg  ( .ip(n6076), .ck(HCLK_top), 
        .rb(1'b1), .s(n12738), .q(\CORTEXM0DS_INST/u_logic/Wv9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/An83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nrivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12738), .q(\CORTEXM0DS_INST/cm0_r02 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yx73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/X1lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12738), .q(\CORTEXM0DS_INST/cm0_r02 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/S8k2z4_reg  ( .ip(n6086), .ck(HCLK_top), 
        .rb(1'b1), .s(n12738), .q(\CORTEXM0DS_INST/u_logic/Azdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hak2z4_reg  ( .ip(n6085), .ck(HCLK_top), 
        .rb(1'b1), .s(n12738), .q(\CORTEXM0DS_INST/u_logic/L0evx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jw73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/M6lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12738), .q(\CORTEXM0DS_INST/cm0_r02 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nz73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ixkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12738), .q(\CORTEXM0DS_INST/cm0_r02 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/H783z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sakvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12737), .q(\CORTEXM0DS_INST/cm0_r02 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zb83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dsjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12737), .q(\CORTEXM0DS_INST/cm0_r02 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wj83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/G5jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12737), .q(\CORTEXM0DS_INST/cm0_r02 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dwl2z4_reg  ( .ip(n6062), .ck(HCLK_top), 
        .rb(1'b1), .s(n12737), .q(\CORTEXM0DS_INST/u_logic/Roevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rxl2z4_reg  ( .ip(n6028), .ck(HCLK_top), 
        .rb(1'b1), .s(n12737), .q(\CORTEXM0DS_INST/u_logic/B19vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Po83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ymivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12737), .q(\CORTEXM0DS_INST/cm0_r02 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/O0o2z4_reg  ( .ip(n6126), .ck(HCLK_top), 
        .rb(1'b1), .s(n12737), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Od83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Onjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12737), .q(\CORTEXM0DS_INST/cm0_r02 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/E0d3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/R8ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12737), .q(\CORTEXM0DS_INST/cm0_r00 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Df83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zijvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12737), .q(\CORTEXM0DS_INST/cm0_r02 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qyc3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gdivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12737), .q(\CORTEXM0DS_INST/cm0_r00 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rr73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/X0mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12737), .q(\CORTEXM0DS_INST/cm0_r02 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wqd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cwivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/cm0_r02 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wce3z4_reg  ( .ip(n6102), .ck(HCLK_top), 
        .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/Rddvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ufy2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/G8nvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/G8fvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gtp2z4_reg  ( .ip(n6060), .ck(HCLK_top), 
        .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/Lrevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Owq2z4_reg  ( .ip(n6059), .ck(HCLK_top), 
        .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/Vsevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F0y2z4_reg  ( .ip(n6058), .ck(HCLK_top), 
        .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/Fuevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I3y2z4_reg  ( .ip(n6057), .ck(HCLK_top), 
        .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/Pvevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/W4y2z4_reg  ( .ip(n6056), .ck(HCLK_top), 
        .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/Zwevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/K6y2z4_reg  ( .ip(n6055), .ck(HCLK_top), 
        .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/Jyevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Y7y2z4_reg  ( .ip(n6054), .ck(HCLK_top), 
        .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/Tzevx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M9y2z4_reg  ( .ip(n6053), .ck(HCLK_top), 
        .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/D1fvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bby2z4_reg  ( .ip(n6052), .ck(HCLK_top), 
        .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/u_logic/O2fvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qcy2z4_reg  ( .ip(n6051), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/Z3fvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fey2z4_reg  ( .ip(n6049), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/V6fvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F1x2z4_reg  ( .ip(n6032), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/Bwfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U2x2z4_reg  ( .ip(n6031), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/Aj9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ydw2z4_reg  ( .ip(n6047), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/Cbfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mfw2z4_reg  ( .ip(n6046), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/Mcfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ahw2z4_reg  ( .ip(n6045), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/Wdfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Oiw2z4_reg  ( .ip(n6044), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/Gffvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jky2z4_reg  ( .ip(n6026), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/P39vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ckw2z4_reg  ( .ip(n6043), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/Qgfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xly2z4_reg  ( .ip(n6025), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/W49vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qlw2z4_reg  ( .ip(n6042), .ck(HCLK_top), 
        .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/u_logic/Aifvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lny2z4_reg  ( .ip(n6024), .ck(HCLK_top), 
        .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/u_logic/D69vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Enw2z4_reg  ( .ip(n6041), .ck(HCLK_top), 
        .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/u_logic/Kjfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zoy2z4_reg  ( .ip(n6023), .ck(HCLK_top), 
        .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/u_logic/K79vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sow2z4_reg  ( .ip(n6040), .ck(HCLK_top), 
        .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/u_logic/Ukfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nqy2z4_reg  ( .ip(n6022), .ck(HCLK_top), 
        .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/u_logic/R89vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gqw2z4_reg  ( .ip(n6039), .ck(HCLK_top), 
        .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/u_logic/Emfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bsy2z4_reg  ( .ip(n6021), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/Y99vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Urw2z4_reg  ( .ip(n6038), .ck(HCLK_top), 
        .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/u_logic/Onfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pty2z4_reg  ( .ip(n6020), .ck(HCLK_top), 
        .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/u_logic/Fb9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Itw2z4_reg  ( .ip(n6037), .ck(HCLK_top), 
        .rb(1'b1), .s(n12738), .q(\CORTEXM0DS_INST/u_logic/Yofvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dvy2z4_reg  ( .ip(n6019), .ck(HCLK_top), 
        .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/u_logic/Mc9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xuw2z4_reg  ( .ip(n6036), .ck(HCLK_top), 
        .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/u_logic/Jqfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mww2z4_reg  ( .ip(n6035), .ck(HCLK_top), 
        .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Urfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Byw2z4_reg  ( .ip(n6034), .ck(HCLK_top), 
        .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Ftfvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qem2z4_reg  ( .ip(n6030), .ck(HCLK_top), 
        .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Kg9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/O5t2z4_reg  ( .ip(n6109), .ck(HCLK_top), 
        .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Fjgvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/R1w2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ocnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/vis_ipsr [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fgm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pthvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Tjh2z4 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wzy2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rghvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Tjh2z4 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sjj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Awhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Tjh2z4 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rni2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jxhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Tjh2z4 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/K9z2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wfhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Ks9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/W7z2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dghvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Gr9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I6z2z4_reg  ( .ip(n6112), .ck(HCLK_top), 
        .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Cq9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jwf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sdhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/vis_pc [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tme3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nehvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/vis_pc [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gmd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uehvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/vis_pc [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/V4d3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bfhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/vis_pc [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vvx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mhhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/vis_pc [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jux2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Thhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/vis_pc [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lrx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hihvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/vis_pc [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zpx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Oihvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/vis_pc [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jex2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Skhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/vis_pc [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cax2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nlhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/vis_pc [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/R8x2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ulhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/vis_pc [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/G7x2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bmhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/vis_pc [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J0l2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wthvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/vis_pc [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qzq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tinvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/u_logic/Ik9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fzl2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jdnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/u_logic/Ml9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zcn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/U2mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/u_logic/Qm9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Uup2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/N2mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/u_logic/Un9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lgi3z4_reg  ( .ip(n6087), .ck(HCLK_top), 
        .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/u_logic/Pxdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qzw2z4_reg  ( .ip(n6033), .ck(HCLK_top), 
        .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/u_logic/Qufvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wai2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lyhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/u_logic/Dw8vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/C3z2z4_reg  ( .ip(n6074), .ck(HCLK_top), 
        .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/u_logic/Bx9vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/T1d3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ifhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/u_logic/Vu8vx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ftf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/P7ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r14 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Arh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ecivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r14 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/E913z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tgivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_r14 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Q713z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xpivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/cm0_r14 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/B613z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Muivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r14 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F8e3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bzivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/cm0_r14 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kzf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/F8jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/cm0_r14 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tz03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yljvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/cm0_r14 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ey03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nqjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r14 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ixh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cvjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r14 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Avg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rzjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r14 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/P9h3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/G4kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/cm0_r14 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bv03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rdkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/cm0_r14 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nt03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gikvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r14 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zr03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vmkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r14 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fli3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zvkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r14 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wo03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/H0lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r14 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hn03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/W4lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r14 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Skh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/L9lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r14 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sl03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Aelvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r14 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Y6i3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wilvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r14 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ek03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vslvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r14 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qi03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ctlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r14 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nf03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qtlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r14 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yd03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xtlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r14 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wa03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qpivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r12 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/H903z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fuivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/cm0_r12 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Q6e3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uyivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/cm0_r12 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vxf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Y7jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/cm0_r12 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z203z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rljvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/cm0_r12 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/K103z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gqjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/cm0_r12 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tvh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vujvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/cm0_r12 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ltg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kzjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/cm0_r12 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/A8h3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Z3kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/cm0_r12 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hyz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kdkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/cm0_r12 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Twz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zhkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/cm0_r12 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fvz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Omkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/cm0_r12 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qji3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Svkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12731), .q(\CORTEXM0DS_INST/cm0_r12 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Csz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/A0lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/cm0_r12 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nqz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/P4lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/cm0_r12 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Djh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/E9lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/cm0_r12 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yoz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tdlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/cm0_r12 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J5i3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pilvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/cm0_r12 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Knz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mrlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/cm0_r12 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wlz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Trlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/cm0_r12 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tiz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hslvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/cm0_r12 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ehz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Oslvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/cm0_r12 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qrf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/I7ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/cm0_r12 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lph3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xbivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/cm0_r12 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kc03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mgivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/cm0_r12 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wd23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hoivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/cm0_r11 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hc23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wsivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/cm0_r11 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tyd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lxivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/cm0_r11 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/D923z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/P6jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/cm0_r11 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/K423z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ikjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/cm0_r11 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/V223z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xojvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/cm0_r11 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/G123z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mtjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/cm0_r11 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Olg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Byjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/cm0_r11 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rz13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Q2kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/cm0_r11 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ow13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bckvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/cm0_r11 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Av13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qgkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/cm0_r11 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mt13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Flkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/cm0_r11 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jq13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jukvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r11 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Uo13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rykvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r11 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fn13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/G3lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r11 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ql13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/V7lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r11 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bk13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kclvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r11 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mi13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ghlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r11 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yg13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Eulvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r11 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kf13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lulvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r11 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hc13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zulvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r11 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sa13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gvlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r11 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ilf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Z5ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r11 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mi23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Oaivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r11 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yg23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dfivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r11 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tjf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/S5ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r10 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vr33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Haivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r10 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hq33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Weivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r10 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fn33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Aoivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r10 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ql33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Psivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r10 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Exd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Exivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r10 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mi33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/I6jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r10 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Td33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bkjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r10 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ec33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qojvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r10 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pa33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ftjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r10 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zjg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uxjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/cm0_r10 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/A933z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/J2kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r10 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/X533z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ubkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r10 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J433z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jgkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r10 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/V233z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ykkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r10 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sz23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cukvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r10 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dy23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kykvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r10 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ow23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Z2lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r10 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zu23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/O7lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r10 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kt23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dclvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r10 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vr23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zglvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r10 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hq23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nvlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r10 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/To23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uvlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r10 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ql23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Iwlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r10 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bk23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pwlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r10 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ow43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tnivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r09 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zu43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Isivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r09 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pvd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xwivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r09 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vr43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/B6jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r09 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cn43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ujjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r09 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nl43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jojvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r09 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yj43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ysjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r09 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kig3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nxjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r09 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ji43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/C2kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r09 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gf43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nbkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r09 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sd43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cgkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r09 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ec43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rkkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r09 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/B943z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vtkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r09 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M743z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dykvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r09 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/X543z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/S2lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r09 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I443z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/H7lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r09 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/T243z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wblvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r09 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/E143z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sglvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r09 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qz33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wwlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r09 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cy33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dxlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r09 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zu33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rxlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r09 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kt33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yxlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r09 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Eif3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/L5ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r09 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/E153z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Aaivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r09 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qz43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Peivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r09 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/X563z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mnivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r08 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I463z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bsivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r08 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Aud3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qwivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r08 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/E163z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/U5jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r08 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lw53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Njjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r08 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wu53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cojvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r08 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ht53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rsjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r08 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vgg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gxjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r08 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sr53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/V1kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r08 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Po53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gbkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/cm0_r08 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bn53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vfkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r08 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nl53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kkkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/cm0_r08 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ki53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Otkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/cm0_r08 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vg53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wxkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r08 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gf53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/L2lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r08 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rd53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/A7lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r08 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cc53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pblvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r08 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Na53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lglvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r08 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z853z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fylvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r08 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/L753z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mylvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12739), .q(\CORTEXM0DS_INST/cm0_r08 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I453z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Azlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_r08 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/T253z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hzlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r08 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pgf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/E5ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r08 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Na63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/T9ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r08 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z863z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ieivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r08 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ajn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jpivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r07 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Oas2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ytivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r07 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/B5e3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nyivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r07 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lqr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/R7jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r07 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ozo2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kljvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r07 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Eun2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zpjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r07 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ecp2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Oujvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r07 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wrg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dzjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r07 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Eqq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/S3kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r07 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/V3m2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ddkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r07 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/G4r2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Shkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r07 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ujp2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hmkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r07 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F9j2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lvkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r07 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tel2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tzkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r07 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z3k2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/I4lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r07 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kiq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/X8lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r07 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jlo2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mdlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r07 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vuo2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Iilvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r07 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Skm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dqlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r07 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ruj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kqlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r07 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vhk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yqlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r07 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Isi2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Frlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r07 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fpi2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/B7ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r07 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rdq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qbivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r07 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cvr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fgivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r07 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bqf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/U6ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r06 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wnu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jbivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r06 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Imu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yfivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r06 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gju2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cpivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r06 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rhu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rtivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r06 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M3e3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gyivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r06 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Neu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/K7jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r06 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U9u2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dljvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r06 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F8u2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Spjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r06 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Q6u2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hujvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r06 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hqg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wyjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r06 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/B5u2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/L3kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r06 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Y1u2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wckvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r06 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/K0u2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lhkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r06 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wyt2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Amkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r06 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tvt2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Evkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r06 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Eut2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mzkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r06 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pst2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/B4lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r06 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Art2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Q8lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r06 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lpt2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fdlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r06 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wnt2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bilvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r06 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Imt2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uolvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r06 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ukt2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bplvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r06 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rht2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pplvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r06 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cgt2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wplvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r06 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mhn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Voivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r05 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z8s2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ktivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r05 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/X1e3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zxivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r05 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wor2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/D7jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r05 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zxo2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wkjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r05 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Psn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lpjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r05 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pap2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Aujvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/cm0_r05 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sog3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pyjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/cm0_r05 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Poq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/E3kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r05 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/H2m2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pckvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/cm0_r05 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/S2r2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ehkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r05 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gip2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tlkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/cm0_r05 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vmj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xukvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12739), .q(\CORTEXM0DS_INST/cm0_r05 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Edl2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fzkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/cm0_r05 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/K2k2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/U3lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/cm0_r05 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vgq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/J8lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/cm0_r05 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ujo2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yclvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/cm0_r05 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gto2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uhlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/cm0_r05 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ejm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lnlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r05 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dtj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Snlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r05 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ggk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Golvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r05 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Glj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nolvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r05 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mof3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/N6ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r05 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ccq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cbivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r05 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Otr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rfivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r05 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Psv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ooivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r04 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Arv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dtivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r04 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I0e3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sxivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r04 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wnv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/W6jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r04 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Djv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pkjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r04 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ohv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Epjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r04 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zfv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ttjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r04 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dng3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Iyjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r04 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kev2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/X2kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r04 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hbv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ickvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r04 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/T9v2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xgkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r04 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F8v2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mlkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r04 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/C5v2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qukvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r04 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/N3v2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yykvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r04 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Y1v2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/N3lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r04 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J0v2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/C8lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r04 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Uyu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rclvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r04 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fxu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nhlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r04 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rvu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cmlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r04 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Duu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jmlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r04 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Aru2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xmlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r04 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lpu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Enlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r04 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xmf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/G6ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r04 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fxv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vaivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r04 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rvv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kfivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r04 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gf73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fnivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r03 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rd73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Urivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r03 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lsd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jwivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r03 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Na73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/N5jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r03 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U573z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gjjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12737), .q(\CORTEXM0DS_INST/cm0_r03 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F473z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vnjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/cm0_r03 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Q273z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ksjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(
        \CORTEXM0DS_INST/u_logic/N586 ), .q(\CORTEXM0DS_INST/cm0_r03 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gfg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zwjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r03 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/B173z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/O1kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/cm0_r03 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yx63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zakvx4 ), .ck(HCLK_top), .rb(1'b1), .s(
        \CORTEXM0DS_INST/u_logic/N586 ), .q(\CORTEXM0DS_INST/cm0_r03 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kw63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ofkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/cm0_r03 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wu63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dkkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/cm0_r03 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tr63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Htkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(
        \CORTEXM0DS_INST/u_logic/N586 ), .q(\CORTEXM0DS_INST/cm0_r03 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Eq63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pxkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r03 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Po63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/E2lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/cm0_r03 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/An63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/T6lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(
        \CORTEXM0DS_INST/u_logic/N586 ), .q(\CORTEXM0DS_INST/cm0_r03 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ll63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Iblvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r03 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wj63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Eglvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r03 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ii63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ozlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r03 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ug63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vzlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r03 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rd63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/J0mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r03 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cc63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Q0mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r03 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Aff3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/X4ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r03 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wj73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/M9ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r03 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ii73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Beivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r03 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ldf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Q4ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r02 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ft83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/F9ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r02 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rr83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Udivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/cm0_r02 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Uu73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bblvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/cm0_r02 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ll73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Z1mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12738), .q(\CORTEXM0DS_INST/cm0_r02 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yfn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rmivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/cm0_r01 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/K7s2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Grivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_r01 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hpd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vvivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/cm0_r01 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hnr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Z4jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12737), .q(\CORTEXM0DS_INST/cm0_r01 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kwo2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sijvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r01 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Arn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hnjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/cm0_r01 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/A9p2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wrjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/cm0_r01 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ccg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lwjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r01 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Anq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/A1kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r01 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/T0m2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lakvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r01 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/E1r2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Afkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r01 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sgp2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pjkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r01 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zpj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tskvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r01 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pbl2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bxkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r01 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/V0k2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Q1lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r01 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gfq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/F6lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r01 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fio2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ualvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r01 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rro2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qflvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r01 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gmm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Eenvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r01 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fwj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lenvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r01 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kjk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zenvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r01 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Koj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gfnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r01 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Orj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/J4ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r01 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Naq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Y8ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r01 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Asr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ndivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r01 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vu93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kmivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r00 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gt93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zqivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r00 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Snd3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ovivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r00 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cq93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/S4jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r00 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Uj93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lijvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r00 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fi93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Anjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r00 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qg93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Prjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r00 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nag3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ewjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r00 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bf93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/T0kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/cm0_r00 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yb93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Eakvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r00 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ka93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tekvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r00 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/W893z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ijkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r00 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/R293z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mskvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r00 [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/C193z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uwkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r00 [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nz83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/J1lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r00 [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yx83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Y5lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/cm0_r00 [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jw83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nalvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r00 [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Uu83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jflvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r00 [30]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Unm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bgnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12738), .q(\CORTEXM0DS_INST/cm0_r00 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xti2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wgnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/cm0_r00 [31]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zkk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dhnvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r00 [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Txj2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Minvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r00 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/B9g3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ldhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/vis_pc [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bnx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cjhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/vis_pc [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Plx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jjhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/vis_pc [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zjq2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ithvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/vis_pc [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fhx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ekhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/vis_pc [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dkr2z4_reg  ( .ip(n6101), .ck(HCLK_top), 
        .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/u_logic/Cfdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/S703z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/J3jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r12 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kfr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/C3jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r07 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vdr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/O2jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r05 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lpv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/H2jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r04 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sa23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/A2jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r11 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kt43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/M1jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r09 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/T263z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/F1jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r08 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cc73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Y0jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r03 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gcr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/K0jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r01 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rr93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/D0jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r00 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M413z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Q3jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r14 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cgu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/V2jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r06 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bk33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/T1jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r10 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ll83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/R0jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r02 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ycx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zkhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/vis_pc [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ikz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Aslvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r12 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Eol2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rqlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r07 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qml2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Znlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r05 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Psu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qmlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r04 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wd13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sulvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r11 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ow33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kxlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r09 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/X553z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tylvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r08 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gf63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/C0mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r03 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Spl2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Senvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r01 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Grl2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ignvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r00 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ch03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jtlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r14 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gjt2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Iplvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r06 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fn23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bwlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r10 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Po73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/L1mvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12709), .q(\CORTEXM0DS_INST/cm0_r02 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I793z4_reg  ( .ip(n6080), .ck(HCLK_top), 
        .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/u_logic/C8dvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Szr2z4_reg  ( .ip(n6105), .ck(HCLK_top), 
        .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/u_logic/M9dvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rpe3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Blivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r12 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/W5s2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ukivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r07 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I4s2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gkivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r05 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Duv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zjivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r04 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kf23z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sjivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r11 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cy43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ejivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r09 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/L763z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xiivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r08 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ug73z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qiivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r03 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U2s2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ciivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r01 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cxc3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vhivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r00 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Fre3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ilivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/cm0_r14 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Uku2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nkivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/cm0_r06 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/To33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ljivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/cm0_r10 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dq83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jiivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/cm0_r02 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ufx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lkhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/vis_pc [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rkd3z4_reg  ( .ip(n6103), .ck(HCLK_top), 
        .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/u_logic/Gcdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J4x2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Imhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/vis_pc [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M1j2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hllvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/u_logic/O7evx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Eyr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hhivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/vis_psp [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hue3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wlivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/vis_psp [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cmn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lqivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/vis_psp [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rds2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Avivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/vis_psp [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ibe3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pzivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/vis_psp [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Oir2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/E4jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/vis_psp [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/O2g3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/T8jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/vis_psp [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/S2p2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mmjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/vis_psp [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ixn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Brjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/vis_psp [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M0i3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qvjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/vis_psp [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Eyg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/F0kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/vis_psp [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tch3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/U4kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/vis_psp [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/X6m2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fekvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/vis_psp [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I7r2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uikvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/vis_psp [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wmp2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jnkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/vis_psp [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Joi3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nwkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/vis_psp [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xhl2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/V0lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/vis_psp [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/D7k2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/K5lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/vis_psp [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wnh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Z9lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/vis_psp [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Noo2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Oelvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/vis_psp [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cai3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kjlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/vis_psp [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pfz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mklvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/vis_psp [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Aez2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tklvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/vis_psp [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mcz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Allvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/vis_psp [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Uuf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/D8ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/vis_psp [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Euh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Scivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/vis_psp [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tse3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Plivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/vis_msp [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Okn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Eqivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12705), .q(\CORTEXM0DS_INST/vis_msp [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dcs2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tuivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/vis_msp [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U9e3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Izivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/vis_msp [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zgr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/X3jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/vis_msp [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z0g3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/M8jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/vis_msp [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/D1p2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fmjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/vis_msp [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Tvn2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Uqjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/vis_msp [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xyh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jvjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/vis_msp [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pwg3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yzjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/vis_msp [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ebh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/N4kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/vis_msp [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J5m2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ydkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/vis_msp [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U5r2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Nikvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/vis_msp [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ilp2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cnkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/vis_msp [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Umi3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gwkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_msp [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Igl2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/O0lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_msp [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/O5k2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/D5lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_msp [24]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hmh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/S9lvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_msp [25]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ymo2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Helvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_msp [27]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/N8i3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Djlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_msp [28]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/X2j2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rjlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_msp [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rek2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yjlvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_msp [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cll2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Fklvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_msp [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M4j2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/W7ivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_msp [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Psh3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lcivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_msp [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qwr2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ahivx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12703), .q(\CORTEXM0DS_INST/vis_msp [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Slr2z4_reg  ( .ip(n6100), .ck(HCLK_top), 
        .rb(1'b1), .s(n12719), .q(\CORTEXM0DS_INST/u_logic/Ngdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rbi3z4_reg  ( .ip(n6113), .ck(HCLK_top), 
        .rb(1'b1), .s(n12712), .q(\CORTEXM0DS_INST/u_logic/H0gvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jw93z4_reg  ( .ip(n6081), .ck(HCLK_top), 
        .rb(1'b1), .s(n12723), .q(\CORTEXM0DS_INST/u_logic/E1dvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xx93z4_reg  ( .ip(n6091), .ck(HCLK_top), 
        .rb(1'b1), .s(n12714), .q(\CORTEXM0DS_INST/u_logic/O2dvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ovc3z4_reg  ( .ip(n6090), .ck(HCLK_top), 
        .rb(1'b1), .s(n12718), .q(\CORTEXM0DS_INST/u_logic/Y3dvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Efp2z4_reg  ( .ip(n6089), .ck(HCLK_top), 
        .rb(1'b1), .s(n12739), .q(\CORTEXM0DS_INST/u_logic/I5dvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F2o2z4_reg  ( .ip(n6144), .ck(HCLK_top), 
        .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/C4b3z4_reg  ( .ip(n6143), .ck(HCLK_top), 
        .rb(1'b1), .s(n12734), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M2b3z4_reg  ( .ip(n6142), .ck(HCLK_top), 
        .rb(1'b1), .s(n12704), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/W0b3z4_reg  ( .ip(n6141), .ck(HCLK_top), 
        .rb(1'b1), .s(n12706), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gza3z4_reg  ( .ip(n6140), .ck(HCLK_top), 
        .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qxa3z4_reg  ( .ip(n6139), .ck(HCLK_top), 
        .rb(1'b1), .s(n12721), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z8b3z4_reg  ( .ip(n6138), .ck(HCLK_top), 
        .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dhb3z4_reg  ( .ip(n6137), .ck(HCLK_top), 
        .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M5f3z4_reg  ( .ip(n6136), .ck(HCLK_top), 
        .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Aze3z4_reg  ( .ip(n6135), .ck(HCLK_top), 
        .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zva3z4_reg  ( .ip(n6134), .ck(HCLK_top), 
        .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/She3z4_reg  ( .ip(n6133), .ck(HCLK_top), 
        .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Iua3z4_reg  ( .ip(n6132), .ck(HCLK_top), 
        .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/K7g3z4_reg  ( .ip(n6131), .ck(HCLK_top), 
        .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ddi3z4_reg  ( .ip(n6122), .ck(HCLK_top), 
        .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Uei3z4_reg  ( .ip(n6121), .ck(HCLK_top), 
        .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nbx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Glhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/vis_pc [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ytm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rrkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/vis_msp [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rtz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Drkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r12 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ksm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wqkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r07 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wqm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Iqkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r05 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/R6v2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bqkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r04 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Yr13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Upkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r11 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qa43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gpkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/cm0_r09 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zj53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zokvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12736), .q(\CORTEXM0DS_INST/cm0_r08 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/It63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sokvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12707), .q(\CORTEXM0DS_INST/cm0_r03 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ipm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Eokvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12715), .q(\CORTEXM0DS_INST/cm0_r01 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/G493z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xnkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12713), .q(\CORTEXM0DS_INST/cm0_r00 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mvm2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yrkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(
        \CORTEXM0DS_INST/u_logic/N586 ), .q(\CORTEXM0DS_INST/vis_psp [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Lq03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Krkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12730), .q(\CORTEXM0DS_INST/cm0_r14 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ixt2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Pqkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/cm0_r06 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/H133z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Npkvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/cm0_r10 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/R283z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lokvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/cm0_r02 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dkx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qjhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/vis_pc [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cao2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qhjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/vis_msp [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/O403z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Chjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/cm0_r12 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/N8o2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vgjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/cm0_r07 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Y6o2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Hgjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/cm0_r05 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Skv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Agjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/cm0_r04 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Z523z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tfjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/cm0_r11 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ro43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ffjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/cm0_r09 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ay53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Yejvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12701), .q(\CORTEXM0DS_INST/cm0_r08 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J773z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Rejvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/cm0_r03 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J5o2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Dejvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12702), .q(\CORTEXM0DS_INST/cm0_r01 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jl93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Wdjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r00 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rbo2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xhjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(
        \CORTEXM0DS_INST/u_logic/N586 ), .q(\CORTEXM0DS_INST/vis_psp [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I113z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jhjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12737), .q(\CORTEXM0DS_INST/cm0_r14 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jbu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ogjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12725), .q(\CORTEXM0DS_INST/cm0_r06 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/If33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Mfjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12735), .q(\CORTEXM0DS_INST/cm0_r10 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Sg83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Kejvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12728), .q(\CORTEXM0DS_INST/cm0_r02 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nox2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Vihvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/vis_pc [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/C5n2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/C9kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12727), .q(\CORTEXM0DS_INST/vis_msp [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vzz2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/O8kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/cm0_r12 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/N3n2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/H8kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r07 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Y1n2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/T7kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_r05 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Vcv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/M7kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_r04 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cy13z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/F7kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_r11 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ug43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/R6kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_r09 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Dq53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/K6kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_r08 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mz63z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/D6kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_r03 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J0n2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/P5kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_r01 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Md93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/I5kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_r00 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/R6n2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/J9kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/vis_psp [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pw03z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/V8kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_r14 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/M3u2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/A8kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_r06 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/L733z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Y6kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12700), .q(\CORTEXM0DS_INST/cm0_r10 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/V883z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/W5kvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12710), .q(\CORTEXM0DS_INST/cm0_r02 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rix2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xjhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12733), .q(\CORTEXM0DS_INST/vis_pc [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/F4q2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Bdjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12711), .q(\CORTEXM0DS_INST/vis_msp [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/D603z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ncjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12717), .q(\CORTEXM0DS_INST/cm0_r12 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Q2q2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gcjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12724), .q(\CORTEXM0DS_INST/cm0_r07 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/B1q2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Sbjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12729), .q(\CORTEXM0DS_INST/cm0_r05 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hmv2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Lbjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12720), .q(\CORTEXM0DS_INST/cm0_r04 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/O723z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ebjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12716), .q(\CORTEXM0DS_INST/cm0_r11 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gq43z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Qajvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12732), .q(\CORTEXM0DS_INST/cm0_r09 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Pz53z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Jajvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12722), .q(\CORTEXM0DS_INST/cm0_r08 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Y873z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Cajvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12726), .q(\CORTEXM0DS_INST/cm0_r03 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mzp2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/O9jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12708), .q(\CORTEXM0DS_INST/cm0_r01 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/No93z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/H9jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/cm0_r00 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U5q2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Idjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/vis_psp [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/X213z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Ucjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/cm0_r14 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ycu2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zbjvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/cm0_r06 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xg33z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Xajvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/cm0_r10 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Hi83z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/V9jvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/cm0_r02 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J7q2z4_reg  ( .ip(n6099), .ck(HCLK_top), 
        .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/u_logic/Yhdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Y8q2z4_reg  ( .ip(n6106), .ck(HCLK_top), 
        .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/u_logic/Jjdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Rsa3z4_reg  ( .ip(n6130), .ck(HCLK_top), 
        .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Zfh3z4_reg  ( .ip(n6092), .ck(HCLK_top), 
        .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/u_logic/Itdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ym93z4_reg  ( .ip(n6098), .ck(HCLK_top), 
        .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/u_logic/Ukdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xeo2z4_reg  ( .ip(n6128), .ck(HCLK_top), 
        .rb(1'b1), .s(n12699), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xyk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Duhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/vis_pc [23]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U593z4_reg  ( .ip(n6088), .ck(HCLK_top), 
        .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/u_logic/S6dvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kaf3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Zdhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/vis_pc [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/H4p2z4_reg  ( .ip(n6097), .ck(HCLK_top), 
        .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/u_logic/Fmdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ara3z4_reg  ( .ip(n6129), .ck(HCLK_top), 
        .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/W5p2z4_reg  ( .ip(n6096), .ck(HCLK_top), 
        .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/u_logic/Qndvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Foe3z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Gehvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/vis_pc [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/L7p2z4_reg  ( .ip(n6095), .ck(HCLK_top), 
        .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/u_logic/Bpdvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Jpa3z4_reg  ( .ip(n6125), .ck(HCLK_top), 
        .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/u_logic/Irh2z4 [19]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xsx2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Aihvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/vis_pc [26]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Omk2z4_reg  ( .ip(
        \CORTEXM0DS_INST/u_logic/Tvhvx4 ), .ck(HCLK_top), .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/vis_pc [29]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/B6j2z4_reg  ( .ip(n6107), .ck(HCLK_top), 
        .rb(1'b1), .s(n12698), .q(\CORTEXM0DS_INST/u_logic/Tudvx4 ) );
  drsp_1 \CORTEXM0DS_INST/u_logic/B2i3z4_reg  ( .ip(n5967), .ck(HCLK_top), 
        .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [17]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Ieh3z4_reg  ( .ip(n5966), .ck(HCLK_top), 
        .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [21]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Kxe3z4_reg  ( .ip(n5965), .ck(HCLK_top), 
        .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [9]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/I1h3z4_reg  ( .ip(n5964), .ck(HCLK_top), 
        .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [20]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Cma3z4_reg  ( .ip(n5963), .ck(HCLK_top), 
        .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [22]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/C9a3z4_reg  ( .ip(n5962), .ck(HCLK_top), 
        .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [10]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Bge3z4_reg  ( .ip(n5961), .ck(HCLK_top), 
        .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [11]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/T5g3z4_reg  ( .ip(n5960), .ck(HCLK_top), 
        .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [13]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Xyn2z4_reg  ( .ip(n5959), .ck(HCLK_top), 
        .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [18]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/W3f3z4_reg  ( .ip(n5958), .ck(HCLK_top), 
        .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [8]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Aea3z4_reg  ( .ip(n5957), .ck(HCLK_top), 
        .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [0]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Wia3z4_reg  ( .ip(n5956), .ck(HCLK_top), 
        .rb(1'b1), .s(n12697), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [3]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/J7b3z4_reg  ( .ip(n5955), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [6]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Qfa3z4_reg  ( .ip(n5954), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [1]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Mka3z4_reg  ( .ip(n5953), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [5]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Taa3z4_reg  ( .ip(n5952), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [4]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gha3z4_reg  ( .ip(n5951), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [2]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Nfb3z4_reg  ( .ip(n5950), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [7]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/L7a3z4_reg  ( .ip(n5949), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [12]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/U5a3z4_reg  ( .ip(n5948), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [14]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/Gdo2z4_reg  ( .ip(n5947), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [16]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/D4a3z4_reg  ( .ip(n5946), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [15]) );
  drsp_1 \CORTEXM0DS_INST/u_logic/L8m2z4_reg  ( .ip(n5945), .ck(HCLK_top), 
        .rb(1'b1), .s(n12696), .q(\CORTEXM0DS_INST/u_logic/Czh2z4 [19]) );
  mux2_1 U8 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [19]), .ip2(
        PID_hwdata_top[19]), .s(n12695), .op(n5945) );
  mux2_1 U10 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [15]), .ip2(
        PID_hwdata_top[15]), .s(n12695), .op(n5946) );
  mux2_1 U11 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [16]), .ip2(
        PID_hwdata_top[16]), .s(n12695), .op(n5947) );
  mux2_1 U12 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [14]), .ip2(
        PID_hwdata_top[14]), .s(n12695), .op(n5948) );
  mux2_1 U13 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [12]), .ip2(
        PID_hwdata_top[12]), .s(n12695), .op(n5949) );
  mux2_1 U14 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [7]), .ip2(
        PID_hwdata_top[7]), .s(n12695), .op(n5950) );
  mux2_1 U15 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [2]), .ip2(
        PID_hwdata_top[2]), .s(n12695), .op(n5951) );
  mux2_1 U16 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [4]), .ip2(
        PID_hwdata_top[4]), .s(n12695), .op(n5952) );
  mux2_1 U17 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [5]), .ip2(
        PID_hwdata_top[5]), .s(n12695), .op(n5953) );
  mux2_1 U18 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [1]), .ip2(
        PID_hwdata_top[1]), .s(n12695), .op(n5954) );
  mux2_1 U19 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [6]), .ip2(
        PID_hwdata_top[6]), .s(n12695), .op(n5955) );
  mux2_1 U20 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [3]), .ip2(
        PID_hwdata_top[3]), .s(n12695), .op(n5956) );
  mux2_1 U21 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [0]), .ip2(
        PID_hwdata_top[0]), .s(n12689), .op(n5957) );
  mux2_1 U22 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [8]), .ip2(
        PID_hwdata_top[8]), .s(n12689), .op(n5958) );
  mux2_1 U23 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [18]), .ip2(
        PID_hwdata_top[18]), .s(n12689), .op(n5959) );
  mux2_1 U24 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [13]), .ip2(
        PID_hwdata_top[13]), .s(n12695), .op(n5960) );
  mux2_1 U25 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [11]), .ip2(
        PID_hwdata_top[11]), .s(n12695), .op(n5961) );
  mux2_1 U26 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [10]), .ip2(
        PID_hwdata_top[10]), .s(n12695), .op(n5962) );
  mux2_1 U27 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [22]), .ip2(
        PID_hwdata_top[22]), .s(n12695), .op(n5963) );
  mux2_1 U28 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [20]), .ip2(
        PID_hwdata_top[20]), .s(n12695), .op(n5964) );
  mux2_1 U29 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [9]), .ip2(
        PID_hwdata_top[9]), .s(n12695), .op(n5965) );
  mux2_1 U30 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [21]), .ip2(
        PID_hwdata_top[21]), .s(n12695), .op(n5966) );
  mux2_1 U31 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [17]), .ip2(
        PID_hwdata_top[17]), .s(n12689), .op(n5967) );
  mux2_1 U35 ( .ip1(\CORTEXM0DS_INST/u_logic/S0hvx4 ), .ip2(PID_hwdata_top[1]), 
        .s(n1), .op(n5968) );
  inv_1 U36 ( .ip(HRESETn_top), .op(\CORTEXM0DS_INST/u_logic/N586 ) );
  mux2_1 U37 ( .ip1(\CORTEXM0DS_INST/u_logic/F2hvx4 ), .ip2(PID_hwdata_top[0]), 
        .s(n1), .op(n5969) );
  mux2_1 U41 ( .ip1(\CORTEXM0DS_INST/u_logic/Vogvx4 ), .ip2(PID_hwdata_top[4]), 
        .s(n2), .op(n5970) );
  mux2_1 U42 ( .ip1(\CORTEXM0DS_INST/u_logic/Nngvx4 ), .ip2(PID_hwdata_top[2]), 
        .s(n2), .op(n5971) );
  mux2_1 U43 ( .ip1(\CORTEXM0DS_INST/u_logic/Eg8vx4 ), .ip2(PID_hwdata_top[1]), 
        .s(n2), .op(n5972) );
  mux2_1 U47 ( .ip1(PID_hwdata_top[22]), .ip2(
        \CORTEXM0DS_INST/u_logic/Psh2z4 [0]), .s(n488), .op(n5973) );
  mux2_1 U52 ( .ip1(\CORTEXM0DS_INST/u_logic/Uth2z4 [0]), .ip2(
        PID_hwdata_top[30]), .s(n489), .op(n5974) );
  mux2_1 U53 ( .ip1(PID_hwdata_top[30]), .ip2(
        \CORTEXM0DS_INST/u_logic/Txh2z4 [0]), .s(n488), .op(n5975) );
  nand2_1 U647 ( .ip1(\RAM_hresp_top[0] ), .ip2(n5920), .op(n450) );
  nand2_1 U652 ( .ip1(HREADY_top), .ip2(\CORTEXM0DS_INST/u_logic/Xyfvx4 ), 
        .op(n1186) );
  inv_1 U654 ( .ip(HREADY_top), .op(n5938) );
  mux2_1 U655 ( .ip1(PID_hwrite_top), .ip2(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), 
        .s(n5938), .op(n6006) );
  nand2_1 U802 ( .ip1(\CORTEXM0DS_INST/u_logic/Mf8vx4 ), .ip2(
        PID_hwdata_top[23]), .op(n3226) );
  nand2_1 U806 ( .ip1(\CORTEXM0DS_INST/u_logic/Mf8vx4 ), .ip2(
        PID_hwdata_top[31]), .op(n3227) );
  nand2_1 U998 ( .ip1(HREADY_top), .ip2(PID_hprot_top[0]), .op(n4585) );
  ab_or_c_or_d U1590 ( .ip1(n1062), .ip2(n12686), .ip3(HREADY_top), .ip4(n1061), .op(n1063) );
  nand2_1 U1599 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(HREADY_top), 
        .op(n1709) );
  nand2_1 U1603 ( .ip1(RAM_hrdata_top[14]), .ip2(n1148), .op(n1076) );
  inv_1 U1606 ( .ip(RAM_hrdata_top[30]), .op(n1157) );
  nand2_1 U1616 ( .ip1(RAM_hrdata_top[12]), .ip2(n1148), .op(n1081) );
  nand2_1 U1620 ( .ip1(RAM_hrdata_top[28]), .ip2(n1144), .op(n1079) );
  nand2_1 U1622 ( .ip1(RAM_hrdata_top[27]), .ip2(n1144), .op(n1086) );
  nand2_1 U1627 ( .ip1(RAM_hrdata_top[11]), .ip2(n1148), .op(n1084) );
  nand2_1 U1629 ( .ip1(RAM_hrdata_top[26]), .ip2(n1144), .op(n1091) );
  nand2_1 U1634 ( .ip1(RAM_hrdata_top[10]), .ip2(n1148), .op(n1089) );
  nand2_1 U1636 ( .ip1(RAM_hrdata_top[9]), .ip2(n1148), .op(n1096) );
  nand2_1 U1642 ( .ip1(RAM_hrdata_top[25]), .ip2(n1144), .op(n1094) );
  nand2_1 U1644 ( .ip1(RAM_hrdata_top[8]), .ip2(n1148), .op(n1101) );
  inv_1 U1645 ( .ip(RAM_hrdata_top[24]), .op(n1169) );
  nand2_1 U1652 ( .ip1(RAM_hrdata_top[23]), .ip2(n1144), .op(n1106) );
  nand2_1 U1656 ( .ip1(RAM_hrdata_top[7]), .ip2(n1148), .op(n1104) );
  nand2_1 U1658 ( .ip1(RAM_hrdata_top[22]), .ip2(n1144), .op(n1111) );
  nand2_1 U1663 ( .ip1(RAM_hrdata_top[6]), .ip2(n1148), .op(n1109) );
  nand2_1 U1665 ( .ip1(RAM_hrdata_top[21]), .ip2(n1144), .op(n1116) );
  nand2_1 U1671 ( .ip1(RAM_hrdata_top[5]), .ip2(n1148), .op(n1114) );
  nand2_1 U1673 ( .ip1(RAM_hrdata_top[20]), .ip2(n1144), .op(n1121) );
  nand2_1 U1679 ( .ip1(RAM_hrdata_top[4]), .ip2(n1148), .op(n1119) );
  nand2_1 U1681 ( .ip1(RAM_hrdata_top[19]), .ip2(n1144), .op(n1126) );
  nand2_1 U1687 ( .ip1(RAM_hrdata_top[3]), .ip2(n1148), .op(n1124) );
  nand2_1 U1689 ( .ip1(RAM_hrdata_top[18]), .ip2(n1144), .op(n1131) );
  nand2_1 U1695 ( .ip1(RAM_hrdata_top[2]), .ip2(n1148), .op(n1129) );
  nand2_1 U1697 ( .ip1(RAM_hrdata_top[17]), .ip2(n1144), .op(n1136) );
  nand2_1 U1703 ( .ip1(RAM_hrdata_top[1]), .ip2(n1148), .op(n1134) );
  nand2_1 U1705 ( .ip1(RAM_hrdata_top[16]), .ip2(n1144), .op(n1141) );
  nand2_1 U1711 ( .ip1(RAM_hrdata_top[0]), .ip2(n1148), .op(n1139) );
  nand2_1 U1713 ( .ip1(RAM_hrdata_top[13]), .ip2(n1148), .op(n1147) );
  nand2_1 U1718 ( .ip1(RAM_hrdata_top[29]), .ip2(n1144), .op(n1145) );
  nand2_1 U1720 ( .ip1(RAM_hrdata_top[15]), .ip2(n1148), .op(n1154) );
  inv_1 U1721 ( .ip(RAM_hrdata_top[31]), .op(n1155) );
  nand2_1 U1732 ( .ip1(RAM_hrdata_top[29]), .ip2(n12693), .op(n1160) );
  nand2_1 U1735 ( .ip1(RAM_hrdata_top[28]), .ip2(n12693), .op(n1162) );
  nand2_1 U1738 ( .ip1(RAM_hrdata_top[27]), .ip2(n12693), .op(n1164) );
  nand2_1 U1741 ( .ip1(RAM_hrdata_top[26]), .ip2(n12693), .op(n1166) );
  nand2_1 U1744 ( .ip1(RAM_hrdata_top[25]), .ip2(n12693), .op(n1168) );
  nand2_1 U1749 ( .ip1(RAM_hrdata_top[23]), .ip2(n12693), .op(n1172) );
  nand2_1 U1752 ( .ip1(RAM_hrdata_top[22]), .ip2(n12693), .op(n1174) );
  nand2_1 U1755 ( .ip1(RAM_hrdata_top[21]), .ip2(n12693), .op(n1176) );
  nand2_1 U1758 ( .ip1(RAM_hrdata_top[20]), .ip2(n12693), .op(n1178) );
  nand2_1 U1761 ( .ip1(RAM_hrdata_top[19]), .ip2(n12693), .op(n1180) );
  nand2_1 U1764 ( .ip1(RAM_hrdata_top[18]), .ip2(n12693), .op(n1182) );
  nand2_1 U1767 ( .ip1(RAM_hrdata_top[17]), .ip2(n12693), .op(n1184) );
  nand2_1 U1770 ( .ip1(RAM_hrdata_top[16]), .ip2(n12693), .op(n1188) );
  nand2_1 U2034 ( .ip1(n12692), .ip2(RAM_hrdata_top[14]), .op(n1403) );
  nand2_1 U2036 ( .ip1(RAM_hrdata_top[13]), .ip2(n12692), .op(n1473) );
  nand2_1 U2086 ( .ip1(RAM_hrdata_top[12]), .ip2(n12692), .op(n1476) );
  nand2_1 U2090 ( .ip1(RAM_hrdata_top[11]), .ip2(n12692), .op(n1479) );
  nand2_1 U2094 ( .ip1(RAM_hrdata_top[10]), .ip2(n12692), .op(n1482) );
  nand2_1 U2098 ( .ip1(RAM_hrdata_top[9]), .ip2(n12692), .op(n1485) );
  nand2_1 U2102 ( .ip1(RAM_hrdata_top[8]), .ip2(n12692), .op(n1488) );
  nand2_1 U2106 ( .ip1(RAM_hrdata_top[7]), .ip2(n12692), .op(n1491) );
  nand2_1 U2110 ( .ip1(RAM_hrdata_top[6]), .ip2(n12692), .op(n1495) );
  nand2_1 U2117 ( .ip1(n12692), .ip2(RAM_hrdata_top[5]), .op(n1497) );
  nand2_1 U2119 ( .ip1(RAM_hrdata_top[4]), .ip2(n12692), .op(n1501) );
  nand2_1 U2123 ( .ip1(RAM_hrdata_top[3]), .ip2(n12692), .op(n1505) );
  nand2_1 U2129 ( .ip1(RAM_hrdata_top[2]), .ip2(n12692), .op(n1506) );
  nand2_1 U2132 ( .ip1(RAM_hrdata_top[1]), .ip2(n12692), .op(n1510) );
  nand2_1 U2137 ( .ip1(RAM_hrdata_top[0]), .ip2(n12692), .op(n1515) );
  nor2_1 U2143 ( .ip1(PID_hprot_top[0]), .ip2(n1521), .op(n2212) );
  nand3_1 U2269 ( .ip1(PID_haddr_top[29]), .ip2(PID_haddr_top[30]), .ip3(
        PID_haddr_top[31]), .op(n2208) );
  nor3_1 U2274 ( .ip1(PID_haddr_top[5]), .ip2(PID_haddr_top[9]), .ip3(
        PID_haddr_top[7]), .op(n1672) );
  inv_1 U2275 ( .ip(PID_haddr_top[8]), .op(n1630) );
  nor3_1 U2277 ( .ip1(PID_haddr_top[3]), .ip2(PID_haddr_top[4]), .ip3(n2069), 
        .op(n1629) );
  not_ab_or_c_or_d U2278 ( .ip1(PID_haddr_top[11]), .ip2(n1630), .ip3(n1629), 
        .ip4(PID_haddr_top[6]), .op(n1664) );
  nand3_1 U2314 ( .ip1(n2065), .ip2(PID_haddr_top[10]), .ip3(n1851), .op(n1662) );
  nand2_1 U2315 ( .ip1(PID_haddr_top[8]), .ip2(n1662), .op(n1663) );
  nor2_1 U2317 ( .ip1(PID_haddr_top[8]), .ip2(PID_haddr_top[9]), .op(n1665) );
  not_ab_or_c_or_d U2318 ( .ip1(PID_haddr_top[8]), .ip2(PID_haddr_top[9]), 
        .ip3(PID_haddr_top[6]), .ip4(n1665), .op(n1675) );
  nor2_1 U2319 ( .ip1(PID_haddr_top[9]), .ip2(PID_haddr_top[7]), .op(n1666) );
  nand3_1 U2320 ( .ip1(n1666), .ip2(PID_haddr_top[11]), .ip3(PID_haddr_top[10]), .op(n1670) );
  inv_1 U2322 ( .ip(PID_haddr_top[2]), .op(n1667) );
  nor2_1 U2326 ( .ip1(PID_haddr_top[2]), .ip2(n1944), .op(n1671) );
  nor3_1 U2329 ( .ip1(PID_haddr_top[23]), .ip2(PID_haddr_top[27]), .ip3(
        PID_haddr_top[26]), .op(n2213) );
  nor3_1 U2330 ( .ip1(PID_haddr_top[24]), .ip2(PID_haddr_top[22]), .ip3(
        PID_haddr_top[17]), .op(n1676) );
  nor2_1 U2340 ( .ip1(PID_haddr_top[7]), .ip2(PID_haddr_top[2]), .op(n1685) );
  nor2_1 U2343 ( .ip1(PID_haddr_top[3]), .ip2(PID_haddr_top[5]), .op(n1687) );
  inv_1 U2346 ( .ip(PID_haddr_top[10]), .op(n1691) );
  nand2_1 U2366 ( .ip1(HREADY_top), .ip2(n3217), .op(n4831) );
  nand2_1 U2478 ( .ip1(HREADY_top), .ip2(n1744), .op(n1770) );
  nand2_1 U2534 ( .ip1(HREADY_top), .ip2(n1789), .op(n2120) );
  nand2_1 U2567 ( .ip1(PID_haddr_top[29]), .ip2(n12691), .op(n1813) );
  nand2_1 U2640 ( .ip1(PID_haddr_top[30]), .ip2(n12691), .op(n1870) );
  nand2_1 U2861 ( .ip1(PID_haddr_top[14]), .ip2(n12691), .op(n2057) );
  nand2_1 U2865 ( .ip1(PID_haddr_top[13]), .ip2(n12691), .op(n2060) );
  nand2_1 U2907 ( .ip1(PID_haddr_top[15]), .ip2(n12691), .op(n2095) );
  nand2_1 U2932 ( .ip1(PID_haddr_top[31]), .ip2(n12691), .op(n2122) );
  nand2_1 U2948 ( .ip1(HREADY_top), .ip2(n2135), .op(n2136) );
  nand2_1 U2953 ( .ip1(n2140), .ip2(HREADY_top), .op(n5822) );
  nand2_1 U2987 ( .ip1(HREADY_top), .ip2(n2168), .op(n5780) );
  inv_1 U3029 ( .ip(PID_hprot_top[3]), .op(n2197) );
  nand2_1 U3031 ( .ip1(HREADY_top), .ip2(n2212), .op(n2198) );
  nand2_1 U3044 ( .ip1(n12687), .ip2(HREADY_top), .op(n2205) );
  or4_1 U3100 ( .ip1(PID_hwdata_top[30]), .ip2(PID_hwdata_top[29]), .ip3(
        PID_hwdata_top[27]), .ip4(PID_hwdata_top[25]), .op(n3231) );
  nand3_1 U3101 ( .ip1(PID_hwdata_top[26]), .ip2(n4711), .ip3(
        PID_hwdata_top[22]), .op(n2271) );
  inv_1 U3106 ( .ip(PID_hwdata_top[18]), .op(n2266) );
  and4_1 U3107 ( .ip1(PID_hwdata_top[19]), .ip2(PID_hwdata_top[24]), .ip3(
        PID_hwdata_top[17]), .ip4(n2266), .op(n2267) );
  nand2_1 U3191 ( .ip1(n3224), .ip2(PID_hwdata_top[25]), .op(n2328) );
  nand2_1 U3357 ( .ip1(n12690), .ip2(PID_hwdata_top[15]), .op(n2460) );
  not_ab_or_c_or_d U3365 ( .ip1(n12688), .ip2(PID_hwdata_top[15]), .ip3(n2464), 
        .ip4(n2463), .op(\CORTEXM0DS_INST/u_logic/Syhvx4 ) );
  nand2_1 U3393 ( .ip1(n3224), .ip2(PID_hwdata_top[27]), .op(n2490) );
  nand2_1 U3395 ( .ip1(n3224), .ip2(PID_hwdata_top[28]), .op(n2492) );
  nand2_1 U3408 ( .ip1(n12690), .ip2(PID_hwdata_top[13]), .op(n2500) );
  and2_1 U3410 ( .ip1(n12688), .ip2(PID_hwdata_top[13]), .op(n2502) );
  not_ab_or_c_or_d U3421 ( .ip1(n12688), .ip2(PID_hwdata_top[8]), .ip3(n2512), 
        .ip4(n2511), .op(\CORTEXM0DS_INST/u_logic/P0ivx4 ) );
  nand2_1 U3422 ( .ip1(n12690), .ip2(PID_hwdata_top[8]), .op(n2513) );
  nand2_1 U3424 ( .ip1(n12690), .ip2(PID_hwdata_top[9]), .op(n2514) );
  and2_1 U3441 ( .ip1(n12688), .ip2(PID_hwdata_top[9]), .op(n2528) );
  and2_1 U3444 ( .ip1(n12688), .ip2(PID_hwdata_top[11]), .op(n2531) );
  nand2_1 U3447 ( .ip1(n12690), .ip2(PID_hwdata_top[11]), .op(n2533) );
  nand2_1 U3456 ( .ip1(n12690), .ip2(PID_hwdata_top[10]), .op(n2541) );
  not_ab_or_c_or_d U3460 ( .ip1(n12688), .ip2(PID_hwdata_top[10]), .ip3(n2544), 
        .ip4(n2543), .op(\CORTEXM0DS_INST/u_logic/B0ivx4 ) );
  nand2_1 U3500 ( .ip1(n12690), .ip2(PID_hwdata_top[7]), .op(n2577) );
  nand2_1 U3548 ( .ip1(n12688), .ip2(PID_hwdata_top[2]), .op(n2620) );
  nand2_1 U3552 ( .ip1(n12690), .ip2(PID_hwdata_top[2]), .op(n2623) );
  nand2_1 U3554 ( .ip1(n12690), .ip2(PID_hwdata_top[3]), .op(n2624) );
  not_ab_or_c_or_d U3558 ( .ip1(n12688), .ip2(PID_hwdata_top[3]), .ip3(n2627), 
        .ip4(n2626), .op(\CORTEXM0DS_INST/u_logic/Y1ivx4 ) );
  nand2_1 U3572 ( .ip1(n12688), .ip2(PID_hwdata_top[4]), .op(n2641) );
  nand2_1 U3576 ( .ip1(n12690), .ip2(PID_hwdata_top[4]), .op(n2644) );
  nand2_1 U3578 ( .ip1(n12690), .ip2(PID_hwdata_top[12]), .op(n2645) );
  not_ab_or_c_or_d U3582 ( .ip1(n12688), .ip2(PID_hwdata_top[12]), .ip3(n2648), 
        .ip4(n2647), .op(\CORTEXM0DS_INST/u_logic/Nzhvx4 ) );
  nand2_1 U3617 ( .ip1(n12688), .ip2(PID_hwdata_top[5]), .op(n2683) );
  nand2_1 U3621 ( .ip1(n12690), .ip2(PID_hwdata_top[5]), .op(n2686) );
  nand2_1 U3645 ( .ip1(n12690), .ip2(PID_hwdata_top[6]), .op(n2711) );
  not_ab_or_c_or_d U3649 ( .ip1(n12688), .ip2(PID_hwdata_top[6]), .ip3(n2714), 
        .ip4(n2713), .op(\CORTEXM0DS_INST/u_logic/D1ivx4 ) );
  nand2_1 U3674 ( .ip1(PID_hwdata_top[14]), .ip2(n12688), .op(n2754) );
  nand2_1 U3678 ( .ip1(n12690), .ip2(PID_hwdata_top[14]), .op(n2757) );
  nand2_1 U3698 ( .ip1(n12690), .ip2(PID_hwdata_top[1]), .op(n2774) );
  nand2_1 U3701 ( .ip1(n12688), .ip2(PID_hwdata_top[1]), .op(n2776) );
  nand2_1 U3709 ( .ip1(n12690), .ip2(PID_hwdata_top[0]), .op(n2786) );
  not_ab_or_c_or_d U3713 ( .ip1(n12688), .ip2(PID_hwdata_top[0]), .ip3(n2791), 
        .ip4(n2790), .op(\CORTEXM0DS_INST/u_logic/T2ivx4 ) );
  nand2_1 U3967 ( .ip1(n12694), .ip2(RAM_hrdata_top[13]), .op(n2976) );
  not_ab_or_c_or_d U3979 ( .ip1(RAM_hrdata_top[15]), .ip2(n12694), .ip3(n2984), 
        .ip4(n4241), .op(n3002) );
  not_ab_or_c_or_d U4016 ( .ip1(n12694), .ip2(RAM_hrdata_top[31]), .ip3(n3016), 
        .ip4(n3015), .op(n4130) );
  not_ab_or_c_or_d U4028 ( .ip1(n12694), .ip2(RAM_hrdata_top[23]), .ip3(n3025), 
        .ip4(n3024), .op(n3027) );
  not_ab_or_c_or_d U4053 ( .ip1(RAM_hrdata_top[7]), .ip2(n12694), .ip3(n3049), 
        .ip4(n3048), .op(n4150) );
  nand2_1 U4080 ( .ip1(n12694), .ip2(RAM_hrdata_top[29]), .op(n3067) );
  not_ab_or_c_or_d U4102 ( .ip1(RAM_hrdata_top[5]), .ip2(n12694), .ip3(n3082), 
        .ip4(n3081), .op(n3084) );
  nand2_1 U4123 ( .ip1(n12694), .ip2(RAM_hrdata_top[21]), .op(n3101) );
  mux2_1 U4149 ( .ip1(n3128), .ip2(PID_hwrite_top), .s(n3127), .op(
        \CORTEXM0DS_INST/u_logic/F4nvx4 ) );
  nand2_1 U4187 ( .ip1(n12694), .ip2(RAM_hrdata_top[25]), .op(n3164) );
  nand2_1 U4212 ( .ip1(n12694), .ip2(RAM_hrdata_top[1]), .op(n3178) );
  nand2_1 U4234 ( .ip1(n12694), .ip2(RAM_hrdata_top[9]), .op(n3197) );
  nand2_1 U4242 ( .ip1(n12694), .ip2(RAM_hrdata_top[17]), .op(n3204) );
  nand2_1 U4356 ( .ip1(HREADY_top), .ip2(n3317), .op(n3348) );
  nand2_1 U4418 ( .ip1(HREADY_top), .ip2(n3368), .op(n3392) );
  nand2_1 U4468 ( .ip1(n12694), .ip2(RAM_hrdata_top[14]), .op(n3419) );
  nand2_1 U4502 ( .ip1(n12694), .ip2(RAM_hrdata_top[30]), .op(n3485) );
  nand2_1 U4537 ( .ip1(n12694), .ip2(RAM_hrdata_top[6]), .op(n3514) );
  nand2_1 U4552 ( .ip1(n12694), .ip2(RAM_hrdata_top[22]), .op(n3554) );
  nand2_1 U4939 ( .ip1(n12694), .ip2(RAM_hrdata_top[16]), .op(n3958) );
  nand2_1 U4946 ( .ip1(n12694), .ip2(RAM_hrdata_top[0]), .op(n3962) );
  not_ab_or_c_or_d U4958 ( .ip1(n12694), .ip2(RAM_hrdata_top[8]), .ip3(n3978), 
        .ip4(n3977), .op(n4408) );
  and2_1 U4960 ( .ip1(n12694), .ip2(RAM_hrdata_top[24]), .op(n3979) );
  nand2_1 U5057 ( .ip1(n12694), .ip2(RAM_hrdata_top[12]), .op(n4087) );
  nand2_1 U5061 ( .ip1(n12694), .ip2(RAM_hrdata_top[28]), .op(n4092) );
  nand2_1 U5070 ( .ip1(n12694), .ip2(RAM_hrdata_top[4]), .op(n4097) );
  not_ab_or_c_or_d U5079 ( .ip1(n12694), .ip2(RAM_hrdata_top[20]), .ip3(n4110), 
        .ip4(n4109), .op(n4348) );
  nand2_1 U5138 ( .ip1(n12694), .ip2(RAM_hrdata_top[27]), .op(n4175) );
  not_ab_or_c_or_d U5141 ( .ip1(n12694), .ip2(RAM_hrdata_top[19]), .ip3(n4180), 
        .ip4(n4241), .op(n4185) );
  nand2_1 U5151 ( .ip1(n12694), .ip2(RAM_hrdata_top[11]), .op(n4190) );
  nand2_1 U5161 ( .ip1(n12694), .ip2(RAM_hrdata_top[3]), .op(n4203) );
  nand2_1 U5175 ( .ip1(n12694), .ip2(RAM_hrdata_top[26]), .op(n4227) );
  nand2_1 U5185 ( .ip1(n12694), .ip2(RAM_hrdata_top[10]), .op(n4237) );
  nand2_1 U5191 ( .ip1(n12694), .ip2(RAM_hrdata_top[18]), .op(n4243) );
  nand2_1 U5202 ( .ip1(n12694), .ip2(RAM_hrdata_top[2]), .op(n4263) );
  nand2_1 U5945 ( .ip1(HREADY_top), .ip2(n4626), .op(n4627) );
  mux2_1 U6001 ( .ip1(PID_hwdata_top[6]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [0]), .s(n4704), .op(
        \CORTEXM0DS_INST/u_logic/Ggmvx4 ) );
  mux2_1 U6002 ( .ip1(PID_hwdata_top[7]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [1]), .s(n4704), .op(
        \CORTEXM0DS_INST/u_logic/Zfmvx4 ) );
  mux2_1 U6003 ( .ip1(PID_hwdata_top[14]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [2]), .s(n4704), .op(
        \CORTEXM0DS_INST/u_logic/Sfmvx4 ) );
  mux2_1 U6004 ( .ip1(PID_hwdata_top[15]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [3]), .s(n4704), .op(
        \CORTEXM0DS_INST/u_logic/Lfmvx4 ) );
  mux2_1 U6005 ( .ip1(PID_hwdata_top[22]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [4]), .s(n4704), .op(
        \CORTEXM0DS_INST/u_logic/Efmvx4 ) );
  mux2_1 U6007 ( .ip1(PID_hwdata_top[30]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [6]), .s(n4704), .op(
        \CORTEXM0DS_INST/u_logic/Qemvx4 ) );
  mux2_1 U6010 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [8]), .ip2(
        PID_hwdata_top[6]), .s(n4706), .op(\CORTEXM0DS_INST/u_logic/Kimvx4 )
         );
  mux2_1 U6011 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [9]), .ip2(
        PID_hwdata_top[7]), .s(n4706), .op(\CORTEXM0DS_INST/u_logic/Dimvx4 )
         );
  mux2_1 U6012 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [10]), .ip2(
        PID_hwdata_top[14]), .s(n4706), .op(\CORTEXM0DS_INST/u_logic/Whmvx4 )
         );
  mux2_1 U6013 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [11]), .ip2(
        PID_hwdata_top[15]), .s(n4706), .op(\CORTEXM0DS_INST/u_logic/Phmvx4 )
         );
  mux2_1 U6014 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [12]), .ip2(
        PID_hwdata_top[22]), .s(n4706), .op(\CORTEXM0DS_INST/u_logic/Ihmvx4 )
         );
  mux2_1 U6016 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [14]), .ip2(
        PID_hwdata_top[30]), .s(n4706), .op(\CORTEXM0DS_INST/u_logic/Ugmvx4 )
         );
  mux2_1 U6019 ( .ip1(PID_hwdata_top[6]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [16]), .s(n4708), .op(
        \CORTEXM0DS_INST/u_logic/Okmvx4 ) );
  mux2_1 U6020 ( .ip1(PID_hwdata_top[7]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [17]), .s(n4708), .op(
        \CORTEXM0DS_INST/u_logic/Hkmvx4 ) );
  mux2_1 U6021 ( .ip1(PID_hwdata_top[14]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [18]), .s(n4708), .op(
        \CORTEXM0DS_INST/u_logic/Akmvx4 ) );
  mux2_1 U6022 ( .ip1(PID_hwdata_top[15]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [19]), .s(n4708), .op(
        \CORTEXM0DS_INST/u_logic/Tjmvx4 ) );
  mux2_1 U6023 ( .ip1(PID_hwdata_top[22]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [20]), .s(n4708), .op(
        \CORTEXM0DS_INST/u_logic/Mjmvx4 ) );
  mux2_1 U6025 ( .ip1(PID_hwdata_top[30]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [22]), .s(n4708), .op(
        \CORTEXM0DS_INST/u_logic/Yimvx4 ) );
  mux2_1 U6028 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [24]), .ip2(
        PID_hwdata_top[6]), .s(n4712), .op(\CORTEXM0DS_INST/u_logic/Smmvx4 )
         );
  mux2_1 U6029 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [25]), .ip2(
        PID_hwdata_top[7]), .s(n4712), .op(\CORTEXM0DS_INST/u_logic/Lmmvx4 )
         );
  mux2_1 U6030 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [26]), .ip2(
        PID_hwdata_top[14]), .s(n4712), .op(\CORTEXM0DS_INST/u_logic/Emmvx4 )
         );
  mux2_1 U6031 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [27]), .ip2(
        PID_hwdata_top[15]), .s(n4712), .op(\CORTEXM0DS_INST/u_logic/Xlmvx4 )
         );
  mux2_1 U6032 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [28]), .ip2(
        PID_hwdata_top[22]), .s(n4712), .op(\CORTEXM0DS_INST/u_logic/Qlmvx4 )
         );
  mux2_1 U6034 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [30]), .ip2(
        PID_hwdata_top[30]), .s(n4712), .op(\CORTEXM0DS_INST/u_logic/Clmvx4 )
         );
  nand3_1 U6127 ( .ip1(n4815), .ip2(RAM_hrdata_top[15]), .ip3(n4814), .op(
        n4816) );
  mux2_1 U6710 ( .ip1(\CORTEXM0DS_INST/u_logic/Ki8vx4 ), .ip2(n5664), .s(
        HREADY_top), .op(\CORTEXM0DS_INST/u_logic/Lrhvx4 ) );
  not_ab_or_c_or_d U6887 ( .ip1(PID_haddr_top[29]), .ip2(n5889), .ip3(
        \CORTEXM0DS_INST/u_logic/Q462z4 ), .ip4(n5888), .op(n5893) );
  and2_1 U6892 ( .ip1(PID_hprot_top[2]), .ip2(n5894), .op(
        \CORTEXM0DS_INST/u_logic/N4422 ) );
  inv_1 U6907 ( .ip(PID_haddr_top[14]), .op(n5914) );
  nand2_1 U6908 ( .ip1(PID_haddr_top[17]), .ip2(n5914), .op(n5915) );
  inv_1 U6910 ( .ip(\PID_htrans_top[1] ), .op(n5916) );
  or4_1 U6911 ( .ip1(n5932), .ip2(RAM_hsel_top), .ip3(n5938), .ip4(n5916), 
        .op(n5928) );
  nand2_1 U6916 ( .ip1(n5920), .ip2(RAM_hready_resp_top), .op(
        \interconnect_ip_inst/n5991 ) );
  nand2_1 U6917 ( .ip1(HREADY_top), .ip2(n5932), .op(n5921) );
  nor2_1 U6918 ( .ip1(PID_haddr_top[13]), .ip2(n5921), .op(n5937) );
  nand2_1 U6919 ( .ip1(n5937), .ip2(\PID_htrans_top[1] ), .op(n5940) );
  nor2_1 U6920 ( .ip1(PID_hwrite_top), .ip2(n5940), .op(n5939) );
  inv_1 U6924 ( .ip(PID_hwrite_top), .op(n5924) );
  nor2_1 U6927 ( .ip1(RAM_hsel_top), .ip2(n5938), .op(n5926) );
  inv_1 U6929 ( .ip(i_ssi_ssi_rst_n_top), .op(\interconnect_ip_inst/n11572 )
         );
  nand3_1 U6934 ( .ip1(HREADY_top), .ip2(PID_haddr_top[13]), .ip3(n5932), .op(
        n5933) );
  or2_1 U6935 ( .ip1(PID_haddr_top[12]), .ip2(n5933), .op(n5935) );
  and2_1 U6940 ( .ip1(PID_hmastlock_top), .ip2(n5938), .op(
        \interconnect_ip_inst/n4860 ) );
  inv_1 U6945 ( .ip(\CORTEXM0DS_INST/u_logic/N4816 ), .op(PID_haddr_top[0]) );
  inv_1 U6946 ( .ip(\CORTEXM0DS_INST/u_logic/Jxovx4 ), .op(PID_haddr_top[10])
         );
  inv_1 U6947 ( .ip(\CORTEXM0DS_INST/u_logic/Cqovx4 ), .op(PID_haddr_top[12])
         );
  inv_1 U6948 ( .ip(\CORTEXM0DS_INST/u_logic/N4767 ), .op(PID_haddr_top[13])
         );
  inv_1 U6949 ( .ip(\CORTEXM0DS_INST/u_logic/N4751 ), .op(PID_haddr_top[14])
         );
  inv_1 U6950 ( .ip(\CORTEXM0DS_INST/u_logic/Vpovx4 ), .op(PID_haddr_top[16])
         );
  inv_1 U6951 ( .ip(\CORTEXM0DS_INST/u_logic/Bv0wx4 ), .op(PID_haddr_top[17])
         );
  inv_1 U6952 ( .ip(\CORTEXM0DS_INST/u_logic/Fq0wx4 ), .op(PID_haddr_top[18])
         );
  inv_1 U6953 ( .ip(\CORTEXM0DS_INST/u_logic/Ql0wx4 ), .op(PID_haddr_top[19])
         );
  inv_1 U6954 ( .ip(\CORTEXM0DS_INST/u_logic/N4674 ), .op(PID_haddr_top[1]) );
  inv_1 U6955 ( .ip(\CORTEXM0DS_INST/u_logic/Ug0wx4 ), .op(PID_haddr_top[20])
         );
  inv_1 U6956 ( .ip(\CORTEXM0DS_INST/u_logic/Fc0wx4 ), .op(PID_haddr_top[21])
         );
  inv_1 U6957 ( .ip(\CORTEXM0DS_INST/u_logic/C70wx4 ), .op(PID_haddr_top[22])
         );
  inv_1 U6958 ( .ip(\CORTEXM0DS_INST/u_logic/Y92wx4 ), .op(PID_haddr_top[23])
         );
  inv_1 U6959 ( .ip(\CORTEXM0DS_INST/u_logic/Y1pvx4 ), .op(PID_haddr_top[24])
         );
  inv_1 U6960 ( .ip(\CORTEXM0DS_INST/u_logic/Rnovx4 ), .op(PID_haddr_top[25])
         );
  inv_1 U6961 ( .ip(\CORTEXM0DS_INST/u_logic/Nhzvx4 ), .op(PID_haddr_top[26])
         );
  inv_1 U6962 ( .ip(\CORTEXM0DS_INST/u_logic/Vezvx4 ), .op(PID_haddr_top[27])
         );
  inv_1 U6963 ( .ip(\CORTEXM0DS_INST/u_logic/V2qvx4 ), .op(PID_haddr_top[28])
         );
  inv_1 U6964 ( .ip(\CORTEXM0DS_INST/u_logic/N4518 ), .op(PID_haddr_top[31])
         );
  inv_1 U6965 ( .ip(\CORTEXM0DS_INST/u_logic/Yuovx4 ), .op(PID_haddr_top[4])
         );
  inv_1 U6966 ( .ip(\CORTEXM0DS_INST/u_logic/Rxzvx4 ), .op(PID_haddr_top[5])
         );
  inv_1 U6967 ( .ip(\CORTEXM0DS_INST/u_logic/Hszvx4 ), .op(PID_haddr_top[6])
         );
  inv_1 U6968 ( .ip(\CORTEXM0DS_INST/u_logic/S4qvx4 ), .op(PID_haddr_top[7])
         );
  inv_1 U6969 ( .ip(\CORTEXM0DS_INST/u_logic/N4439 ), .op(PID_haddr_top[30])
         );
  or2_1 U6970 ( .ip1(\CORTEXM0DS_INST/u_logic/E562z4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Q462z4 ), .op(PID_haddr_top[29]) );
  or2_1 U6971 ( .ip1(PID_haddr_top[30]), .ip2(PID_haddr_top[29]), .op(
        PID_hprot_top[2]) );
  inv_1 U6972 ( .ip(\CORTEXM0DS_INST/u_logic/N4422 ), .op(PID_hprot_top[3]) );
  and2_1 U6973 ( .ip1(\CORTEXM0DS_INST/u_logic/A362z4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Oq42z4 ), .op(PID_hsize_top[0]) );
  inv_1 U6974 ( .ip(\CORTEXM0DS_INST/u_logic/N4421 ), .op(PID_hsize_top[1]) );
  inv_1 U6975 ( .ip(\CORTEXM0DS_INST/u_logic/N4396 ), .op(PID_hprot_top[0]) );
  and2_1 U6976 ( .ip1(n6116), .ip2(\CORTEXM0DS_INST/u_logic/Xmywx4 ), .op(
        \PID_htrans_top[1] ) );
  inv_1 U6977 ( .ip(\CORTEXM0DS_INST/u_logic/N4359 ), .op(PID_hwdata_top[0])
         );
  inv_1 U6978 ( .ip(\CORTEXM0DS_INST/u_logic/N4282 ), .op(PID_hwdata_top[24])
         );
  inv_1 U6979 ( .ip(\CORTEXM0DS_INST/u_logic/N4227 ), .op(PID_hwdata_top[25])
         );
  inv_1 U6980 ( .ip(\CORTEXM0DS_INST/u_logic/N4170 ), .op(PID_hwdata_top[26])
         );
  inv_1 U6981 ( .ip(\CORTEXM0DS_INST/u_logic/N4116 ), .op(PID_hwdata_top[27])
         );
  inv_1 U6982 ( .ip(\CORTEXM0DS_INST/u_logic/Sx3wx4 ), .op(PID_hwdata_top[28])
         );
  inv_1 U6983 ( .ip(\CORTEXM0DS_INST/u_logic/N4005 ), .op(PID_hwdata_top[29])
         );
  inv_1 U6984 ( .ip(\CORTEXM0DS_INST/u_logic/N3967 ), .op(PID_hwdata_top[31])
         );
  inv_1 U6985 ( .ip(\CORTEXM0DS_INST/u_logic/N3966 ), .op(PID_hwdata_top[3])
         );
  inv_1 U6986 ( .ip(n6176), .op(PID_hwdata_top[4]) );
  inv_1 U6987 ( .ip(n6181), .op(PID_hwdata_top[5]) );
  inv_1 U6988 ( .ip(\CORTEXM0DS_INST/u_logic/N3946 ), .op(PID_hwdata_top[6])
         );
  inv_1 U6989 ( .ip(n6167), .op(PID_hwdata_top[7]) );
  inv_1 U6990 ( .ip(n6172), .op(PID_hwdata_top[2]) );
  inv_1 U6991 ( .ip(\CORTEXM0DS_INST/u_logic/N3783 ), .op(PID_hwdata_top[30])
         );
  inv_1 U6992 ( .ip(\CORTEXM0DS_INST/u_logic/N2678 ), .op(PID_hwrite_top) );
  inv_1 U6993 ( .ip(\CORTEXM0DS_INST/u_logic/Bq5wx4 ), .op(PID_hwdata_top[14])
         );
  inv_1 U6994 ( .ip(n6190), .op(PID_hwdata_top[1]) );
  inv_1 U6995 ( .ip(\CORTEXM0DS_INST/u_logic/O24wx4 ), .op(PID_hwdata_top[16])
         );
  inv_1 U6996 ( .ip(\CORTEXM0DS_INST/u_logic/N1447 ), .op(PID_haddr_top[15])
         );
  inv_1 U6997 ( .ip(\CORTEXM0DS_INST/u_logic/Xxovx4 ), .op(PID_haddr_top[9])
         );
  inv_1 U6998 ( .ip(\CORTEXM0DS_INST/u_logic/Ekovx4 ), .op(PID_haddr_top[3])
         );
  inv_1 U6999 ( .ip(\CORTEXM0DS_INST/u_logic/Owovx4 ), .op(PID_haddr_top[11])
         );
  inv_1 U7000 ( .ip(\CORTEXM0DS_INST/u_logic/Z6ovx4 ), .op(PID_haddr_top[8])
         );
  inv_1 U7001 ( .ip(\CORTEXM0DS_INST/u_logic/Fvovx4 ), .op(PID_haddr_top[2])
         );
  nand2_1 U7002 ( .ip1(n5978), .ip2(n5977), .op(PID_hwdata_top[23]) );
  nand2_1 U7003 ( .ip1(n5980), .ip2(n5979), .op(PID_hwdata_top[22]) );
  nand2_1 U7004 ( .ip1(n5982), .ip2(n5981), .op(PID_hwdata_top[21]) );
  nand2_1 U7005 ( .ip1(n5984), .ip2(n5983), .op(PID_hwdata_top[19]) );
  nand2_1 U7006 ( .ip1(n5986), .ip2(n5985), .op(PID_hwdata_top[20]) );
  nand2_1 U7007 ( .ip1(n5988), .ip2(n5987), .op(PID_hwdata_top[17]) );
  nand2_1 U7008 ( .ip1(n5990), .ip2(n5989), .op(PID_hwdata_top[18]) );
  nand2_1 U7009 ( .ip1(n5992), .ip2(n5991), .op(PID_hwdata_top[15]) );
  nand2_1 U7010 ( .ip1(n5994), .ip2(n5993), .op(PID_hwdata_top[13]) );
  nand2_1 U7011 ( .ip1(n5996), .ip2(n5995), .op(PID_hwdata_top[12]) );
  nand2_1 U7012 ( .ip1(n5998), .ip2(n5997), .op(PID_hwdata_top[11]) );
  nand2_1 U7013 ( .ip1(n6000), .ip2(n5999), .op(PID_hwdata_top[10]) );
  nand2_1 U7014 ( .ip1(n6002), .ip2(n6001), .op(PID_hwdata_top[9]) );
  nand2_1 U7015 ( .ip1(n6004), .ip2(n6003), .op(PID_hwdata_top[8]) );
  nand4_1 U7016 ( .ip1(n6656), .ip2(n6655), .ip3(n6654), .ip4(n6653), .op(
        n6657) );
  nand4_1 U7017 ( .ip1(n6771), .ip2(n6770), .ip3(n6769), .ip4(n6768), .op(
        n6772) );
  nand4_1 U7018 ( .ip1(n6601), .ip2(n6600), .ip3(n6599), .ip4(n6598), .op(
        n6602) );
  nand4_1 U7019 ( .ip1(n6552), .ip2(n6551), .ip3(n6550), .ip4(n6549), .op(
        n6553) );
  nand4_1 U7020 ( .ip1(n6675), .ip2(n6674), .ip3(n6673), .ip4(n6672), .op(
        n6676) );
  nand4_1 U7021 ( .ip1(n6666), .ip2(n6665), .ip3(n6664), .ip4(n6663), .op(
        n6667) );
  nand4_1 U7022 ( .ip1(n6717), .ip2(n6716), .ip3(n6715), .ip4(n6714), .op(
        n6718) );
  nand4_1 U7023 ( .ip1(n6472), .ip2(n6471), .ip3(n6470), .ip4(n6469), .op(
        n6473) );
  nand4_1 U7024 ( .ip1(n6543), .ip2(n6542), .ip3(n6541), .ip4(n6540), .op(
        n6544) );
  nand4_1 U7025 ( .ip1(n6561), .ip2(n6560), .ip3(n6559), .ip4(n6558), .op(
        n6562) );
  nand4_1 U7026 ( .ip1(n6616), .ip2(n6615), .ip3(n6614), .ip4(n6613), .op(
        n6617) );
  nor4_1 U7027 ( .ip1(n11755), .ip2(n6871), .ip3(n6870), .ip4(n6869), .op(
        n7536) );
  nand4_1 U7028 ( .ip1(n6520), .ip2(n6519), .ip3(n6518), .ip4(n6517), .op(
        n6521) );
  nand4_1 U7029 ( .ip1(n6634), .ip2(n6633), .ip3(n6632), .ip4(n6631), .op(
        n6635) );
  nand4_1 U7030 ( .ip1(n6643), .ip2(n6642), .ip3(n6641), .ip4(n6640), .op(
        n6644) );
  nand4_1 U7031 ( .ip1(n6738), .ip2(n6737), .ip3(n6736), .ip4(n6735), .op(
        n6739) );
  nand4_1 U7032 ( .ip1(n6534), .ip2(n6533), .ip3(n6532), .ip4(n6531), .op(
        n6535) );
  nand4_1 U7033 ( .ip1(n6625), .ip2(n6624), .ip3(n6623), .ip4(n6622), .op(
        n6626) );
  nand4_1 U7034 ( .ip1(n6423), .ip2(n6422), .ip3(n6421), .ip4(n6420), .op(
        n6424) );
  nand4_1 U7035 ( .ip1(n6816), .ip2(n6815), .ip3(n6814), .ip4(n6813), .op(
        n6817) );
  nand4_1 U7036 ( .ip1(n6684), .ip2(n6683), .ip3(n6682), .ip4(n6681), .op(
        n6685) );
  nand4_1 U7037 ( .ip1(n6574), .ip2(n6573), .ip3(n6572), .ip4(n6571), .op(
        n6575) );
  nand4_1 U7038 ( .ip1(n6493), .ip2(n6492), .ip3(n6491), .ip4(n6490), .op(
        n6494) );
  nand4_1 U7039 ( .ip1(n6693), .ip2(n6692), .ip3(n6691), .ip4(n6690), .op(
        n6694) );
  nand4_1 U7040 ( .ip1(n6652), .ip2(n6651), .ip3(n6650), .ip4(n6649), .op(
        n6695) );
  nand4_1 U7041 ( .ip1(n6570), .ip2(n6569), .ip3(n6568), .ip4(n6567), .op(
        n6612) );
  nor4_1 U7042 ( .ip1(n6873), .ip2(n6872), .ip3(n10938), .ip4(n11195), .op(
        n6874) );
  nand4_1 U7043 ( .ip1(n6880), .ip2(n6879), .ip3(n6878), .ip4(n6877), .op(
        n6881) );
  nor4_1 U7044 ( .ip1(n7575), .ip2(n6452), .ip3(n6451), .ip4(n6450), .op(n6453) );
  nand4_1 U7045 ( .ip1(n6255), .ip2(n6254), .ip3(n12650), .ip4(n6253), .op(
        n6256) );
  nand4_1 U7046 ( .ip1(n6417), .ip2(n6416), .ip3(n11722), .ip4(n6415), .op(
        n7827) );
  nand4_1 U7047 ( .ip1(n6921), .ip2(n6920), .ip3(n6919), .ip4(n6918), .op(
        n6922) );
  nand4_1 U7048 ( .ip1(n6853), .ip2(n6852), .ip3(n6851), .ip4(n6850), .op(
        n6854) );
  nand4_1 U7049 ( .ip1(n7007), .ip2(n7006), .ip3(n7005), .ip4(n7004), .op(
        n7008) );
  nand4_1 U7050 ( .ip1(n7028), .ip2(n7027), .ip3(n7026), .ip4(n7025), .op(
        n7029) );
  nand4_1 U7051 ( .ip1(n7046), .ip2(n7045), .ip3(n7044), .ip4(n7043), .op(
        n7047) );
  nand4_1 U7052 ( .ip1(n7037), .ip2(n7036), .ip3(n7035), .ip4(n7034), .op(
        n7038) );
  nor4_1 U7053 ( .ip1(n10970), .ip2(n11752), .ip3(n10472), .ip4(n6209), .op(
        n6220) );
  nand4_1 U7054 ( .ip1(n8230), .ip2(n8229), .ip3(n8228), .ip4(n8227), .op(
        n8231) );
  nand4_1 U7055 ( .ip1(n8194), .ip2(n8193), .ip3(n8192), .ip4(n8191), .op(
        n8195) );
  nand4_1 U7056 ( .ip1(n8121), .ip2(n8120), .ip3(n8119), .ip4(n8118), .op(
        n8122) );
  nand4_1 U7057 ( .ip1(n8052), .ip2(n8051), .ip3(n8050), .ip4(n8049), .op(
        n8053) );
  nand4_1 U7058 ( .ip1(n7942), .ip2(n7941), .ip3(n7940), .ip4(n7939), .op(
        n7943) );
  nand4_1 U7059 ( .ip1(n8348), .ip2(n8347), .ip3(n8346), .ip4(n8345), .op(
        n8349) );
  nand4_1 U7060 ( .ip1(n7655), .ip2(n7654), .ip3(n7653), .ip4(n7652), .op(
        n7656) );
  nand4_1 U7061 ( .ip1(n7626), .ip2(n7625), .ip3(n7624), .ip4(n7623), .op(
        n7627) );
  nand4_1 U7062 ( .ip1(n7686), .ip2(n7685), .ip3(n7684), .ip4(n7683), .op(
        n7687) );
  nand4_1 U7063 ( .ip1(n7599), .ip2(n7598), .ip3(n7597), .ip4(n7596), .op(
        n7600) );
  nand4_1 U7064 ( .ip1(n7561), .ip2(n7560), .ip3(n7559), .ip4(n7558), .op(
        n7562) );
  nand4_1 U7065 ( .ip1(n6938), .ip2(n6937), .ip3(n6936), .ip4(n6935), .op(
        n6939) );
  nand4_1 U7066 ( .ip1(n6291), .ip2(n6290), .ip3(n6289), .ip4(n6288), .op(
        n8577) );
  nand4_1 U7067 ( .ip1(n6304), .ip2(n6303), .ip3(n6302), .ip4(n6301), .op(
        n8576) );
  nand4_1 U7068 ( .ip1(n7364), .ip2(n7363), .ip3(n7362), .ip4(n7361), .op(
        n7365) );
  nand4_1 U7069 ( .ip1(n6904), .ip2(n6903), .ip3(n6902), .ip4(n6901), .op(
        n6905) );
  nand4_1 U7070 ( .ip1(n6334), .ip2(n6333), .ip3(n6332), .ip4(n6331), .op(
        n8585) );
  nand4_1 U7071 ( .ip1(n11698), .ip2(n11697), .ip3(n6210), .ip4(n11700), .op(
        n6340) );
  nor4_1 U7072 ( .ip1(n6374), .ip2(n9520), .ip3(n6373), .ip4(n9582), .op(n6380) );
  nand4_1 U7073 ( .ip1(n8213), .ip2(n8212), .ip3(n8211), .ip4(n8210), .op(
        n8214) );
  nand4_1 U7074 ( .ip1(n8209), .ip2(n8208), .ip3(n8207), .ip4(n8206), .op(
        n8215) );
  nand4_1 U7075 ( .ip1(n8180), .ip2(n8179), .ip3(n8178), .ip4(n8177), .op(
        n8181) );
  nand4_1 U7076 ( .ip1(n8176), .ip2(n8175), .ip3(n8174), .ip4(n8173), .op(
        n8182) );
  nand4_1 U7077 ( .ip1(n8106), .ip2(n8105), .ip3(n8104), .ip4(n8103), .op(
        n8107) );
  nand4_1 U7078 ( .ip1(n8102), .ip2(n8101), .ip3(n8100), .ip4(n8099), .op(
        n8108) );
  nand4_1 U7079 ( .ip1(n8067), .ip2(n8066), .ip3(n8065), .ip4(n8064), .op(
        n8073) );
  nand4_1 U7080 ( .ip1(n8071), .ip2(n8070), .ip3(n8069), .ip4(n8068), .op(
        n8072) );
  nand4_1 U7081 ( .ip1(n8037), .ip2(n8036), .ip3(n8035), .ip4(n8034), .op(
        n8038) );
  nand4_1 U7082 ( .ip1(n8033), .ip2(n8032), .ip3(n8031), .ip4(n8030), .op(
        n8039) );
  nand4_1 U7083 ( .ip1(n7862), .ip2(n7861), .ip3(n7860), .ip4(n7859), .op(
        n7863) );
  nand4_1 U7084 ( .ip1(n7841), .ip2(n7840), .ip3(n7839), .ip4(n7838), .op(
        n7842) );
  nand4_1 U7085 ( .ip1(n7837), .ip2(n7836), .ip3(n7835), .ip4(n7834), .op(
        n7843) );
  nand4_1 U7086 ( .ip1(n7442), .ip2(n7441), .ip3(n7440), .ip4(n7439), .op(
        n7443) );
  nand4_1 U7087 ( .ip1(n7438), .ip2(n7437), .ip3(n7436), .ip4(n7435), .op(
        n7444) );
  nand4_1 U7088 ( .ip1(n8246), .ip2(n8245), .ip3(n8244), .ip4(n8243), .op(
        n8251) );
  nand4_1 U7089 ( .ip1(n6220), .ip2(n6219), .ip3(n6218), .ip4(n6345), .op(
        n6221) );
  nand4_1 U7090 ( .ip1(n6888), .ip2(n6887), .ip3(n6886), .ip4(n6885), .op(
        n6889) );
  nand4_1 U7091 ( .ip1(n7371), .ip2(n7370), .ip3(n7369), .ip4(n7368), .op(
        n7372) );
  nand4_1 U7092 ( .ip1(n7693), .ip2(n7692), .ip3(n7691), .ip4(n7690), .op(
        n7694) );
  nand4_1 U7093 ( .ip1(n7661), .ip2(n7660), .ip3(n7659), .ip4(n7658), .op(
        n7662) );
  nand4_1 U7094 ( .ip1(n7634), .ip2(n7633), .ip3(n7632), .ip4(n7631), .op(
        n7635) );
  nand4_1 U7095 ( .ip1(n7604), .ip2(n7603), .ip3(n7602), .ip4(n7601), .op(
        n7605) );
  nand4_1 U7096 ( .ip1(n7566), .ip2(n7565), .ip3(n7564), .ip4(n7563), .op(
        n7567) );
  nand4_1 U7097 ( .ip1(n7527), .ip2(n7526), .ip3(n7525), .ip4(n7524), .op(
        n7528) );
  nand4_1 U7098 ( .ip1(n7490), .ip2(n7489), .ip3(n7488), .ip4(n7487), .op(
        n7491) );
  nand4_1 U7099 ( .ip1(n7456), .ip2(n7455), .ip3(n7454), .ip4(n7453), .op(
        n7457) );
  nand4_1 U7100 ( .ip1(n8304), .ip2(n8303), .ip3(n8302), .ip4(n8301), .op(
        n8305) );
  nand4_1 U7101 ( .ip1(n8158), .ip2(n8157), .ip3(n8156), .ip4(n8155), .op(
        n8159) );
  nand4_1 U7102 ( .ip1(n8089), .ip2(n8088), .ip3(n8087), .ip4(n8086), .op(
        n8090) );
  nand4_1 U7103 ( .ip1(n8020), .ip2(n8019), .ip3(n8018), .ip4(n8017), .op(
        n8021) );
  nand4_1 U7104 ( .ip1(n7910), .ip2(n7909), .ip3(n7908), .ip4(n7907), .op(
        n7911) );
  nand4_1 U7105 ( .ip1(n7874), .ip2(n7873), .ip3(n7872), .ip4(n7871), .op(
        n7875) );
  nand4_1 U7106 ( .ip1(n7816), .ip2(n7815), .ip3(n7814), .ip4(n7813), .op(
        n7817) );
  nand4_1 U7107 ( .ip1(n8354), .ip2(n8353), .ip3(n8352), .ip4(n8351), .op(
        n9160) );
  nand4_1 U7108 ( .ip1(n8953), .ip2(n8952), .ip3(n8951), .ip4(n8950), .op(
        n8954) );
  nand4_1 U7109 ( .ip1(n8894), .ip2(n8893), .ip3(n8892), .ip4(n8891), .op(
        n8895) );
  nand4_1 U7110 ( .ip1(n8838), .ip2(n8837), .ip3(n8836), .ip4(n8835), .op(
        n8839) );
  nor4_1 U7111 ( .ip1(n6336), .ip2(n11851), .ip3(n12011), .ip4(n11859), .op(
        n8588) );
  nand4_1 U7112 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10539), .ip3(
        n10734), .ip4(n11038), .op(n8813) );
  nand4_1 U7113 ( .ip1(n8873), .ip2(n8872), .ip3(n8871), .ip4(n8870), .op(
        n8878) );
  nand4_1 U7114 ( .ip1(n6269), .ip2(n6268), .ip3(n6267), .ip4(n6266), .op(
        n2140) );
  nand4_1 U7115 ( .ip1(n8332), .ip2(n8331), .ip3(n8330), .ip4(n8329), .op(
        n8333) );
  nand4_1 U7116 ( .ip1(n8328), .ip2(n8327), .ip3(n8326), .ip4(n8325), .op(
        n8334) );
  nor4_1 U7117 ( .ip1(n10679), .ip2(n6279), .ip3(n10678), .ip4(n11652), .op(
        n6342) );
  nand4_1 U7118 ( .ip1(n8929), .ip2(n8928), .ip3(n8927), .ip4(n8926), .op(
        n8930) );
  nand4_1 U7119 ( .ip1(n8921), .ip2(n8920), .ip3(n8919), .ip4(n8918), .op(
        n8931) );
  nor4_1 U7120 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip4(n10771), .op(n12627) );
  nand4_1 U7121 ( .ip1(n7589), .ip2(n7588), .ip3(n7587), .ip4(n7586), .op(
        n7590) );
  nand4_1 U7122 ( .ip1(n7585), .ip2(n7584), .ip3(n7583), .ip4(n7582), .op(
        n7591) );
  nand4_1 U7123 ( .ip1(n7544), .ip2(n7543), .ip3(n7542), .ip4(n7541), .op(
        n7545) );
  nand4_1 U7124 ( .ip1(n7540), .ip2(n7539), .ip3(n7538), .ip4(n7537), .op(
        n7546) );
  nand4_1 U7125 ( .ip1(n6436), .ip2(n6435), .ip3(n6434), .ip4(n6433), .op(
        n6437) );
  nand4_1 U7126 ( .ip1(n6826), .ip2(n6825), .ip3(n6824), .ip4(n6823), .op(
        n6827) );
  nand4_1 U7127 ( .ip1(n8186), .ip2(n8185), .ip3(n8184), .ip4(n8183), .op(
        n8187) );
  nand4_1 U7128 ( .ip1(n8140), .ip2(n8139), .ip3(n8138), .ip4(n8137), .op(
        n8141) );
  nand4_1 U7129 ( .ip1(n8136), .ip2(n8135), .ip3(n8134), .ip4(n8133), .op(
        n8142) );
  nand4_1 U7130 ( .ip1(n8001), .ip2(n8000), .ip3(n7999), .ip4(n7998), .op(
        n8002) );
  nand4_1 U7131 ( .ip1(n7997), .ip2(n7996), .ip3(n7995), .ip4(n7994), .op(
        n8003) );
  nand4_1 U7132 ( .ip1(n7964), .ip2(n7963), .ip3(n7962), .ip4(n7961), .op(
        n7965) );
  nand4_1 U7133 ( .ip1(n7960), .ip2(n7959), .ip3(n7958), .ip4(n7957), .op(
        n7966) );
  nand4_1 U7134 ( .ip1(n7926), .ip2(n7925), .ip3(n7924), .ip4(n7923), .op(
        n7932) );
  nand4_1 U7135 ( .ip1(n7930), .ip2(n7929), .ip3(n7928), .ip4(n7927), .op(
        n7931) );
  nand4_1 U7136 ( .ip1(n7896), .ip2(n7895), .ip3(n7894), .ip4(n7893), .op(
        n7897) );
  nand4_1 U7137 ( .ip1(n7892), .ip2(n7891), .ip3(n7890), .ip4(n7889), .op(
        n7898) );
  nand4_1 U7138 ( .ip1(n7868), .ip2(n7867), .ip3(n7866), .ip4(n7865), .op(
        n7869) );
  nand4_1 U7139 ( .ip1(n7512), .ip2(n7511), .ip3(n7510), .ip4(n7509), .op(
        n7513) );
  nand4_1 U7140 ( .ip1(n7508), .ip2(n7507), .ip3(n7506), .ip4(n7505), .op(
        n7514) );
  nand4_1 U7141 ( .ip1(n7847), .ip2(n7846), .ip3(n7845), .ip4(n7844), .op(
        n7848) );
  nand4_1 U7142 ( .ip1(n7475), .ip2(n7474), .ip3(n7473), .ip4(n7472), .op(
        n7476) );
  nand4_1 U7143 ( .ip1(n7471), .ip2(n7470), .ip3(n7469), .ip4(n7468), .op(
        n7477) );
  nand4_1 U7144 ( .ip1(n7448), .ip2(n7447), .ip3(n7446), .ip4(n7445), .op(
        n7449) );
  nand4_1 U7145 ( .ip1(n7405), .ip2(n7404), .ip3(n7403), .ip4(n7402), .op(
        n7406) );
  nand4_1 U7146 ( .ip1(n7401), .ip2(n7400), .ip3(n7399), .ip4(n7398), .op(
        n7407) );
  nand4_1 U7147 ( .ip1(n8282), .ip2(n8281), .ip3(n8280), .ip4(n8279), .op(
        n8283) );
  nand4_1 U7148 ( .ip1(n8278), .ip2(n8277), .ip3(n8276), .ip4(n8275), .op(
        n8284) );
  nand4_1 U7149 ( .ip1(n8857), .ip2(n8856), .ip3(n8855), .ip4(n8854), .op(
        n8858) );
  nand4_1 U7150 ( .ip1(n8255), .ip2(n8254), .ip3(n8253), .ip4(n8252), .op(
        n8256) );
  nand4_1 U7151 ( .ip1(n6845), .ip2(n11191), .ip3(n12305), .ip4(n12600), .op(
        n2209) );
  nand4_1 U7152 ( .ip1(n6409), .ip2(n6408), .ip3(n6407), .ip4(n6406), .op(
        n6410) );
  nand4_1 U7153 ( .ip1(n6810), .ip2(n6809), .ip3(n6808), .ip4(n6807), .op(
        n6811) );
  nand4_1 U7154 ( .ip1(n7699), .ip2(n7698), .ip3(n7697), .ip4(n7696), .op(
        n12233) );
  nand4_1 U7155 ( .ip1(n7420), .ip2(n7419), .ip3(n7418), .ip4(n7417), .op(
        n7421) );
  nand4_1 U7156 ( .ip1(n8263), .ip2(n8262), .ip3(n8261), .ip4(n8260), .op(
        n8264) );
  nand4_1 U7157 ( .ip1(n8095), .ip2(n8094), .ip3(n8093), .ip4(n8092), .op(
        n12201) );
  nand4_1 U7158 ( .ip1(n8026), .ip2(n8025), .ip3(n8024), .ip4(n8023), .op(
        n12222) );
  nand4_1 U7159 ( .ip1(n7916), .ip2(n7915), .ip3(n7914), .ip4(n7913), .op(
        n12253) );
  nand4_1 U7160 ( .ip1(n7822), .ip2(n7821), .ip3(n7820), .ip4(n7819), .op(
        n12274) );
  nand4_1 U7161 ( .ip1(n8963), .ip2(n8962), .ip3(n8961), .ip4(n8960), .op(
        n8964) );
  nand4_1 U7162 ( .ip1(n8900), .ip2(n8899), .ip3(n8898), .ip4(n8897), .op(
        n9122) );
  nand4_1 U7163 ( .ip1(n8844), .ip2(n8843), .ip3(n8842), .ip4(n8841), .op(
        n9776) );
  nand4_1 U7164 ( .ip1(n9002), .ip2(n9653), .ip3(n6797), .ip4(n8457), .op(
        n6798) );
  nand4_1 U7165 ( .ip1(n8869), .ip2(n8868), .ip3(n8867), .ip4(n8866), .op(
        n8886) );
  nand4_1 U7166 ( .ip1(n8338), .ip2(n8337), .ip3(n8336), .ip4(n8335), .op(
        n8339) );
  nand4_1 U7167 ( .ip1(n6206), .ip2(n12042), .ip3(n6205), .ip4(n6204), .op(
        n10908) );
  nor4_1 U7168 ( .ip1(n12068), .ip2(n12390), .ip3(n12373), .ip4(n12362), .op(
        n6206) );
  nand4_1 U7169 ( .ip1(n8938), .ip2(n8937), .ip3(n8936), .ip4(n8935), .op(
        n8939) );
  nand4_1 U7170 ( .ip1(n7595), .ip2(n7594), .ip3(n7593), .ip4(n7592), .op(
        n12658) );
  nand4_1 U7171 ( .ip1(n7553), .ip2(n7552), .ip3(n7551), .ip4(n7550), .op(
        n7554) );
  nand4_1 U7172 ( .ip1(n6934), .ip2(n6933), .ip3(n6932), .ip4(n6931), .op(
        n12667) );
  nand4_1 U7173 ( .ip1(n6867), .ip2(n6866), .ip3(n6865), .ip4(n6864), .op(
        n12673) );
  nand4_1 U7174 ( .ip1(n7360), .ip2(n7359), .ip3(n7358), .ip4(n7357), .op(
        n12671) );
  nand4_1 U7175 ( .ip1(n7681), .ip2(n7680), .ip3(n7679), .ip4(n7678), .op(
        n12675) );
  nand4_1 U7176 ( .ip1(n8007), .ip2(n8006), .ip3(n8005), .ip4(n8004), .op(
        n12676) );
  nand4_1 U7177 ( .ip1(n7650), .ip2(n7649), .ip3(n7648), .ip4(n7647), .op(
        n12677) );
  nand4_1 U7178 ( .ip1(n7970), .ip2(n7969), .ip3(n7968), .ip4(n7967), .op(
        n12678) );
  nand4_1 U7179 ( .ip1(n7622), .ip2(n7621), .ip3(n7620), .ip4(n7619), .op(
        n12681) );
  nand4_1 U7180 ( .ip1(n7936), .ip2(n7935), .ip3(n7934), .ip4(n7933), .op(
        n7937) );
  nand4_1 U7181 ( .ip1(n7902), .ip2(n7901), .ip3(n7900), .ip4(n7899), .op(
        n7903) );
  nand4_1 U7182 ( .ip1(n7518), .ip2(n7517), .ip3(n7516), .ip4(n7515), .op(
        n7519) );
  nand4_1 U7183 ( .ip1(n8863), .ip2(n8862), .ip3(n8861), .ip4(n8860), .op(
        n8864) );
  nand4_1 U7184 ( .ip1(n9841), .ip2(n6238), .ip3(n6237), .ip4(n6236), .op(
        n12305) );
  nor4_1 U7185 ( .ip1(n8558), .ip2(n8557), .ip3(n9836), .ip4(n8556), .op(
        \CORTEXM0DS_INST/u_logic/N2678 ) );
  nand4_1 U7186 ( .ip1(n9841), .ip2(n9840), .ip3(n9839), .ip4(n10731), .op(
        n9842) );
  inv_1 U7187 ( .ip(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .op(n10865) );
  inv_1 U7188 ( .ip(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .op(n11754) );
  nand2_1 U7189 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(n11754), .op(
        n12613) );
  inv_1 U7190 ( .ip(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .op(n12095) );
  inv_1 U7191 ( .ip(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .op(n10547) );
  nor2_1 U7192 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10547), .op(
        n9597) );
  inv_1 U7193 ( .ip(n9597), .op(n7094) );
  inv_1 U7194 ( .ip(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .op(n11730) );
  inv_1 U7195 ( .ip(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .op(n12625) );
  nor2_1 U7196 ( .ip1(n11730), .ip2(n12625), .op(n11654) );
  inv_1 U7197 ( .ip(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(n6210) );
  nand2_1 U7198 ( .ip1(n11654), .ip2(n6210), .op(n8831) );
  nor4_1 U7199 ( .ip1(n10865), .ip2(n12613), .ip3(n7094), .ip4(n8831), .op(
        TXEV_top_out) );
  inv_1 U7200 ( .ip(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .op(n12686) );
  inv_1 U7201 ( .ip(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .op(n11038) );
  nor2_1 U7202 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Cn8vx4 ), .op(n9639) );
  nor2_1 U7203 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n10547), .op(
        n10937) );
  nor2_1 U7204 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n10547), .op(
        n11651) );
  inv_1 U7205 ( .ip(n11651), .op(n8823) );
  inv_1 U7206 ( .ip(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .op(n12096) );
  nand2_1 U7207 ( .ip1(n12096), .ip2(n11038), .op(n10770) );
  nor2_1 U7208 ( .ip1(n11754), .ip2(n10770), .op(n11744) );
  inv_1 U7209 ( .ip(n11744), .op(n11231) );
  or2_1 U7210 ( .ip1(n8823), .ip2(n11231), .op(n6198) );
  nor2_1 U7211 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [4]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [5]), .op(n6300) );
  inv_1 U7212 ( .ip(\CORTEXM0DS_INST/vis_ipsr [3]), .op(n6322) );
  nand2_1 U7213 ( .ip1(n6300), .ip2(n6322), .op(n9781) );
  nor4_1 U7214 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [1]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [2]), .ip3(\CORTEXM0DS_INST/vis_ipsr [0]), 
        .ip4(n9781), .op(n11769) );
  nand2_1 U7215 ( .ip1(\CORTEXM0DS_INST/vis_pc [28]), .ip2(
        \CORTEXM0DS_INST/vis_pc [29]), .op(n10417) );
  nor2_1 U7216 ( .ip1(n11769), .ip2(n10417), .op(n6196) );
  nand4_1 U7217 ( .ip1(\CORTEXM0DS_INST/vis_pc [27]), .ip2(
        \CORTEXM0DS_INST/u_logic/Hx8vx4 ), .ip3(\CORTEXM0DS_INST/vis_pc [30]), 
        .ip4(n6196), .op(n11771) );
  nand2_1 U7218 ( .ip1(n12625), .ip2(n11771), .op(n10489) );
  or2_1 U7219 ( .ip1(n10489), .ip2(n11231), .op(n6197) );
  nand2_1 U7220 ( .ip1(n6198), .ip2(n6197), .op(n6201) );
  nor2_1 U7221 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n12095), .op(
        n11206) );
  nor2_1 U7222 ( .ip1(n11206), .ip2(n10865), .op(n10648) );
  nor2_1 U7223 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n10770), .op(
        n11697) );
  inv_1 U7224 ( .ip(n11697), .op(n6199) );
  nor2_1 U7225 ( .ip1(n10648), .ip2(n6199), .op(n6200) );
  not_ab_or_c_or_d U7226 ( .ip1(n9639), .ip2(n10937), .ip3(n6201), .ip4(n6200), 
        .op(n6208) );
  nor4_1 U7227 ( .ip1(\CORTEXM0DS_INST/u_logic/Bx9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Wv9vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Su9vx4 ), .ip4(
        \CORTEXM0DS_INST/u_logic/Ot9vx4 ), .op(n8698) );
  inv_1 U7228 ( .ip(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .op(n12065) );
  nor2_1 U7229 ( .ip1(n8698), .ip2(n12065), .op(n12068) );
  nor3_1 U7230 ( .ip1(\CORTEXM0DS_INST/u_logic/Wv9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Su9vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Ot9vx4 ), .op(n6202) );
  inv_1 U7231 ( .ip(\CORTEXM0DS_INST/u_logic/Bx9vx4 ), .op(n12376) );
  nor2_1 U7232 ( .ip1(n6202), .ip2(n12376), .op(n12390) );
  inv_1 U7233 ( .ip(\CORTEXM0DS_INST/u_logic/Su9vx4 ), .op(n12365) );
  inv_1 U7234 ( .ip(\CORTEXM0DS_INST/u_logic/Ot9vx4 ), .op(n11159) );
  nor2_1 U7235 ( .ip1(n12365), .ip2(n11159), .op(n12373) );
  nor2_1 U7236 ( .ip1(\CORTEXM0DS_INST/u_logic/Su9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Ot9vx4 ), .op(n8656) );
  inv_1 U7237 ( .ip(\CORTEXM0DS_INST/u_logic/Wv9vx4 ), .op(n12356) );
  nor2_1 U7238 ( .ip1(n8656), .ip2(n12356), .op(n12362) );
  nand2_1 U7239 ( .ip1(n8698), .ip2(n12065), .op(n8675) );
  nand2_1 U7240 ( .ip1(\CORTEXM0DS_INST/u_logic/Cq9vx4 ), .ip2(n8675), .op(
        n12042) );
  nor2_1 U7241 ( .ip1(n8675), .ip2(\CORTEXM0DS_INST/u_logic/Cq9vx4 ), .op(
        n6203) );
  inv_1 U7242 ( .ip(n6203), .op(n10040) );
  nand2_1 U7243 ( .ip1(\CORTEXM0DS_INST/u_logic/Gr9vx4 ), .ip2(n10040), .op(
        n6205) );
  inv_1 U7244 ( .ip(\CORTEXM0DS_INST/u_logic/Gr9vx4 ), .op(n10038) );
  nand2_1 U7245 ( .ip1(n6203), .ip2(n10038), .op(n10030) );
  nand2_1 U7246 ( .ip1(\CORTEXM0DS_INST/u_logic/Ks9vx4 ), .ip2(n10030), .op(
        n6204) );
  nand2_1 U7247 ( .ip1(n11754), .ip2(n10908), .op(n9722) );
  inv_1 U7248 ( .ip(n9722), .op(n10936) );
  nand2_1 U7249 ( .ip1(n10547), .ip2(n11730), .op(n12603) );
  nor3_1 U7250 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n12096), .ip3(
        n12603), .op(n10661) );
  nand2_1 U7251 ( .ip1(n10936), .ip2(n10661), .op(n6207) );
  nor2_1 U7252 ( .ip1(n12096), .ip2(n6210), .op(n11184) );
  nand2_1 U7253 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n11184), .op(
        n10816) );
  nor2_1 U7254 ( .ip1(n10865), .ip2(n10816), .op(n10586) );
  nand2_1 U7255 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10586), .op(
        n10498) );
  nand3_1 U7256 ( .ip1(n6208), .ip2(n6207), .ip3(n10498), .op(n6223) );
  inv_1 U7257 ( .ip(\CORTEXM0DS_INST/u_logic/Ki8vx4 ), .op(n10894) );
  nand3_1 U7258 ( .ip1(n10894), .ip2(\CORTEXM0DS_INST/vis_pc [2]), .ip3(
        \CORTEXM0DS_INST/u_logic/Eg8vx4 ), .op(n11089) );
  inv_1 U7259 ( .ip(n11089), .op(n9723) );
  and3_1 U7260 ( .ip1(n10936), .ip2(n9723), .ip3(n10661), .op(n6222) );
  inv_1 U7261 ( .ip(\CORTEXM0DS_INST/u_logic/Q5gvx4 ), .op(n9700) );
  nor2_1 U7262 ( .ip1(n12095), .ip2(n11730), .op(n12078) );
  nand2_1 U7263 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n12078), .op(
        n11035) );
  nor3_1 U7264 ( .ip1(n6210), .ip2(n9700), .ip3(n11035), .op(n10970) );
  nand2_1 U7265 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(n12095), .op(
        n8986) );
  nand2_1 U7266 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Z6gvx4 ), .op(n10943) );
  or2_1 U7267 ( .ip1(n11730), .ip2(n10943), .op(n10800) );
  nor2_1 U7268 ( .ip1(n8986), .ip2(n10800), .op(n11752) );
  nor3_1 U7269 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip3(n10800), .op(n10472) );
  nand2_1 U7270 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n10865), .op(
        n9620) );
  nor2_1 U7271 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n6210), .op(
        n8495) );
  inv_1 U7272 ( .ip(n8495), .op(n10665) );
  nor2_1 U7273 ( .ip1(n9620), .ip2(n10665), .op(n6209) );
  inv_1 U7274 ( .ip(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .op(n12338) );
  nor2_1 U7275 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n12338), .op(
        n11736) );
  nand2_1 U7276 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n11730), .op(
        n12614) );
  nor2_1 U7277 ( .ip1(n11754), .ip2(n12614), .op(n9757) );
  nor2_1 U7278 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n6210), .op(
        n10539) );
  inv_1 U7279 ( .ip(n12613), .op(n10734) );
  nor2_1 U7280 ( .ip1(n11730), .ip2(n8813), .op(n10495) );
  nand3_1 U7281 ( .ip1(n11730), .ip2(n10865), .ip3(n11038), .op(n8678) );
  inv_1 U7282 ( .ip(n8678), .op(n10727) );
  nor2_1 U7283 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n11730), .op(
        n8819) );
  nor2_1 U7284 ( .ip1(n12095), .ip2(n12625), .op(n10822) );
  nand2_1 U7285 ( .ip1(n8819), .ip2(n10822), .op(n6254) );
  nor2_1 U7286 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n6254), .op(
        n6799) );
  or2_1 U7287 ( .ip1(n10727), .ip2(n6799), .op(n6212) );
  or2_1 U7288 ( .ip1(n11736), .ip2(n6799), .op(n6211) );
  nand2_1 U7289 ( .ip1(n6212), .ip2(n6211), .op(n6213) );
  nor2_1 U7290 ( .ip1(n6213), .ip2(n12613), .op(n6214) );
  not_ab_or_c_or_d U7291 ( .ip1(n11736), .ip2(n9757), .ip3(n10495), .ip4(n6214), .op(n6219) );
  nor2_1 U7292 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .op(n10880) );
  nor2_1 U7293 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n12096), .op(
        n10874) );
  inv_1 U7294 ( .ip(n10874), .op(n11729) );
  nor2_1 U7295 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n11729), .op(
        n11745) );
  nand2_1 U7296 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n12095), .op(
        n11751) );
  nor2_1 U7297 ( .ip1(n12096), .ip2(n11751), .op(n11198) );
  inv_1 U7298 ( .ip(n11198), .op(n11132) );
  or2_1 U7299 ( .ip1(n11132), .ip2(n6210), .op(n6216) );
  nand2_1 U7300 ( .ip1(n12095), .ip2(n11730), .op(n11212) );
  inv_1 U7301 ( .ip(n11212), .op(n11746) );
  nor2_1 U7302 ( .ip1(n9620), .ip2(n9700), .op(n12079) );
  nand2_1 U7303 ( .ip1(n11746), .ip2(n12079), .op(n10475) );
  or2_1 U7304 ( .ip1(n10475), .ip2(n6210), .op(n6215) );
  nand2_1 U7305 ( .ip1(n6216), .ip2(n6215), .op(n6217) );
  inv_1 U7306 ( .ip(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .op(n10949) );
  nor4_1 U7307 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10865), .ip3(
        n12686), .ip4(n10949), .op(n6355) );
  not_ab_or_c_or_d U7308 ( .ip1(n10880), .ip2(n11745), .ip3(n6217), .ip4(n6355), .op(n6218) );
  nand2_1 U7309 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n10865), .op(
        n11168) );
  nand2_1 U7310 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n11754), .op(
        n10903) );
  nor3_1 U7311 ( .ip1(n6210), .ip2(n11168), .ip3(n10903), .op(n6374) );
  nand3_1 U7312 ( .ip1(n10734), .ip2(n6374), .ip3(n12095), .op(n6345) );
  not_ab_or_c_or_d U7313 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n6223), 
        .ip3(n6222), .ip4(n6221), .op(n6845) );
  nor2_1 U7314 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n12686), .op(
        n10779) );
  inv_1 U7315 ( .ip(n10779), .op(n11191) );
  nor2_1 U7316 ( .ip1(n12614), .ip2(n9620), .op(n6230) );
  nor2_1 U7317 ( .ip1(n10547), .ip2(n12096), .op(n10027) );
  or2_1 U7318 ( .ip1(n6230), .ip2(n10027), .op(n6225) );
  or2_1 U7319 ( .ip1(n9722), .ip2(n10027), .op(n6224) );
  nand2_1 U7320 ( .ip1(n6225), .ip2(n6224), .op(n9841) );
  nor2_1 U7321 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n11754), .op(
        n9570) );
  inv_1 U7322 ( .ip(n9570), .op(n6226) );
  or2_1 U7323 ( .ip1(n6226), .ip2(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(n6228) );
  nor2_1 U7324 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n10547), .op(
        n10713) );
  nand2_1 U7325 ( .ip1(n10713), .ip2(n11038), .op(n10900) );
  inv_1 U7326 ( .ip(n10900), .op(n10726) );
  nand2_1 U7327 ( .ip1(n10726), .ip2(n12095), .op(n11130) );
  or2_1 U7328 ( .ip1(n11130), .ip2(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(
        n6227) );
  nand2_1 U7329 ( .ip1(n6228), .ip2(n6227), .op(n9831) );
  nor2_1 U7330 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n10865), .op(
        n10830) );
  nand2_1 U7331 ( .ip1(n10830), .ip2(n11754), .op(n10677) );
  nor2_1 U7332 ( .ip1(n10547), .ip2(n10677), .op(n6229) );
  not_ab_or_c_or_d U7333 ( .ip1(n6230), .ip2(n12338), .ip3(n9831), .ip4(n6229), 
        .op(n6238) );
  nand2_1 U7334 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Vdgvx4 ), .op(n11750) );
  inv_1 U7335 ( .ip(n11750), .op(n12032) );
  nand2_1 U7336 ( .ip1(n12032), .ip2(n6210), .op(n11084) );
  nor2_1 U7337 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n12625), .op(
        n9634) );
  nand2_1 U7338 ( .ip1(n12096), .ip2(n12338), .op(n8738) );
  nor2_1 U7339 ( .ip1(n11754), .ip2(n8738), .op(n11177) );
  nand2_1 U7340 ( .ip1(n9634), .ip2(n11177), .op(n6231) );
  nand2_1 U7341 ( .ip1(n11084), .ip2(n6231), .op(n6232) );
  nor2_1 U7342 ( .ip1(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Mj8vx4 ), .op(n10728) );
  inv_1 U7343 ( .ip(n10728), .op(n12608) );
  nor2_1 U7344 ( .ip1(n10770), .ip2(n12608), .op(n10959) );
  nor2_1 U7345 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .op(n11169) );
  nand2_1 U7346 ( .ip1(n10959), .ip2(n11169), .op(n10934) );
  inv_1 U7347 ( .ip(n10934), .op(n9652) );
  not_ab_or_c_or_d U7348 ( .ip1(n12686), .ip2(n6232), .ip3(n9652), .ip4(n10495), .op(n6237) );
  nand2_1 U7349 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n10865), .op(
        n10771) );
  inv_1 U7350 ( .ip(n10771), .op(n12607) );
  nand2_1 U7351 ( .ip1(n10547), .ip2(n6210), .op(n8993) );
  nor2_1 U7352 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Efgvx4 ), .op(n12628) );
  nand2_1 U7353 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n11038), .op(
        n12649) );
  inv_1 U7354 ( .ip(n12649), .op(n11650) );
  nand2_1 U7355 ( .ip1(n12628), .ip2(n11650), .op(n9009) );
  nor3_1 U7356 ( .ip1(n12625), .ip2(n8993), .ip3(n9009), .op(n6235) );
  inv_1 U7357 ( .ip(n6254), .op(n11743) );
  nor3_1 U7358 ( .ip1(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip2(n8738), .ip3(
        n8678), .op(n10906) );
  nor3_1 U7359 ( .ip1(\CORTEXM0DS_INST/u_logic/Q5gvx4 ), .ip2(n10771), .ip3(
        n10943), .op(n9702) );
  not_ab_or_c_or_d U7360 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n11743), .ip3(n10906), .ip4(n9702), .op(n6233) );
  nor2_1 U7361 ( .ip1(n6233), .ip2(n10949), .op(n6234) );
  not_ab_or_c_or_d U7362 ( .ip1(n11752), .ip2(n12607), .ip3(n6235), .ip4(n6234), .op(n6236) );
  inv_1 U7363 ( .ip(n11751), .op(n10776) );
  or2_1 U7364 ( .ip1(n10776), .ip2(n11206), .op(n6240) );
  or2_1 U7365 ( .ip1(n10665), .ip2(n11206), .op(n6239) );
  nand2_1 U7366 ( .ip1(n6240), .ip2(n6239), .op(n8564) );
  nand2_1 U7367 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(n8553) );
  inv_1 U7368 ( .ip(n8553), .op(n9869) );
  nor2_1 U7369 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .op(n9598) );
  nand2_1 U7370 ( .ip1(n11730), .ip2(n11038), .op(n10781) );
  nor2_1 U7371 ( .ip1(n10949), .ip2(n6210), .op(n11200) );
  nand2_1 U7372 ( .ip1(n11200), .ip2(n10880), .op(n6241) );
  nand2_1 U7373 ( .ip1(n10781), .ip2(n6241), .op(n6242) );
  not_ab_or_c_or_d U7374 ( .ip1(n9869), .ip2(n10822), .ip3(n9598), .ip4(n6242), 
        .op(n9813) );
  inv_1 U7375 ( .ip(n9813), .op(n8563) );
  nor2_1 U7376 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n12095), .op(
        n8456) );
  nand2_1 U7377 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n10949), .op(
        n8826) );
  inv_1 U7378 ( .ip(n8826), .op(n11170) );
  nand2_1 U7379 ( .ip1(n10949), .ip2(n6210), .op(n8996) );
  inv_1 U7380 ( .ip(n8996), .op(n11182) );
  nand2_1 U7381 ( .ip1(n11182), .ip2(n10822), .op(n9530) );
  inv_1 U7382 ( .ip(n9530), .op(n6246) );
  nand2_1 U7383 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(n10892) );
  inv_1 U7384 ( .ip(n10892), .op(n6999) );
  nor2_1 U7385 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Whgvx4 ), .op(n11715) );
  nand2_1 U7386 ( .ip1(n6999), .ip2(n11715), .op(n6244) );
  nand2_1 U7387 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n6210), .op(
        n10588) );
  inv_1 U7388 ( .ip(n10588), .op(n10708) );
  nand3_1 U7389 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n11654), .ip3(
        n10708), .op(n6243) );
  not_ab_or_c_or_d U7390 ( .ip1(n6244), .ip2(n6243), .ip3(
        \CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip4(n12338), .op(n6245) );
  not_ab_or_c_or_d U7391 ( .ip1(n8456), .ip2(n11170), .ip3(n6246), .ip4(n6245), 
        .op(n6269) );
  nand2_1 U7392 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n12686), .op(
        n12615) );
  inv_1 U7393 ( .ip(n12615), .op(n11229) );
  or4_1 U7394 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(n11651), .ip3(
        n10539), .ip4(n10776), .op(n6263) );
  nor2_1 U7395 ( .ip1(n12096), .ip2(n12686), .op(n12405) );
  inv_1 U7396 ( .ip(n10713), .op(n11211) );
  nor2_1 U7397 ( .ip1(n12625), .ip2(n11211), .op(n6257) );
  inv_1 U7398 ( .ip(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .op(n12075) );
  inv_1 U7399 ( .ip(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .op(n12329) );
  nor2_1 U7400 ( .ip1(n12329), .ip2(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .op(
        n11033) );
  and2_1 U7401 ( .ip1(n12075), .ip2(n11033), .op(n10679) );
  inv_1 U7402 ( .ip(\CORTEXM0DS_INST/u_logic/Ho8vx4 ), .op(n10811) );
  nand2_1 U7403 ( .ip1(n12329), .ip2(n10811), .op(n10782) );
  inv_1 U7404 ( .ip(n10782), .op(n9657) );
  nor3_1 U7405 ( .ip1(n9657), .ip2(n11033), .ip3(n12075), .op(n6279) );
  nor3_1 U7406 ( .ip1(n10679), .ip2(n6279), .ip3(n8738), .op(n6247) );
  nand2_1 U7407 ( .ip1(n6247), .ip2(n11754), .op(n6250) );
  inv_1 U7408 ( .ip(\CORTEXM0DS_INST/u_logic/K79vx4 ), .op(n12564) );
  not_ab_or_c_or_d U7409 ( .ip1(\CORTEXM0DS_INST/u_logic/W49vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/D69vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/R89vx4 ), .ip4(n12564), .op(n9571) );
  nand2_1 U7410 ( .ip1(n12075), .ip2(n12338), .op(n10652) );
  nor3_1 U7411 ( .ip1(n9571), .ip2(n11730), .ip3(n10652), .op(n6344) );
  nand2_1 U7412 ( .ip1(n6344), .ip2(n11754), .op(n6249) );
  inv_1 U7413 ( .ip(n8738), .op(n11725) );
  nand3_1 U7414 ( .ip1(n11654), .ip2(n11725), .ip3(n12075), .op(n6248) );
  nand3_1 U7415 ( .ip1(n6250), .ip2(n6249), .ip3(n6248), .op(n6252) );
  inv_1 U7416 ( .ip(n11184), .op(n12616) );
  nor2_1 U7417 ( .ip1(n12616), .ip2(n11212), .op(n6251) );
  nor2_1 U7418 ( .ip1(n6210), .ip2(n11729), .op(n10790) );
  not_ab_or_c_or_d U7419 ( .ip1(\CORTEXM0DS_INST/u_logic/Rkgvx4 ), .ip2(n6252), 
        .ip3(n6251), .ip4(n10790), .op(n6255) );
  nand2_1 U7420 ( .ip1(n11206), .ip2(n10728), .op(n12650) );
  nand3_1 U7421 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n10734), .ip3(
        n12686), .op(n6253) );
  not_ab_or_c_or_d U7422 ( .ip1(n12405), .ip2(n11754), .ip3(n6257), .ip4(n6256), .op(n6258) );
  nor2_1 U7423 ( .ip1(n6258), .ip2(n10865), .op(n6262) );
  nand2_1 U7424 ( .ip1(n11177), .ip2(n10547), .op(n10646) );
  or2_1 U7425 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10646), .op(
        n6260) );
  or2_1 U7426 ( .ip1(n11168), .ip2(n10646), .op(n6259) );
  nand2_1 U7427 ( .ip1(n6260), .ip2(n6259), .op(n6261) );
  not_ab_or_c_or_d U7428 ( .ip1(n11229), .ip2(n6263), .ip3(n6262), .ip4(n6261), 
        .op(n6268) );
  or2_1 U7429 ( .ip1(n8993), .ip2(n9009), .op(n6267) );
  nand4_1 U7430 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n11654), .ip3(
        n10734), .ip4(n12095), .op(n6264) );
  nand2_1 U7431 ( .ip1(n12096), .ip2(n10949), .op(n11214) );
  inv_1 U7432 ( .ip(n11214), .op(n7001) );
  nand2_1 U7433 ( .ip1(n7001), .ip2(n11754), .op(n8987) );
  nand2_1 U7434 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n12625), .op(
        n8623) );
  nand3_1 U7435 ( .ip1(n10779), .ip2(n8987), .ip3(n8623), .op(n6356) );
  nand2_1 U7436 ( .ip1(n6264), .ip2(n6356), .op(n6265) );
  nand2_1 U7437 ( .ip1(\CORTEXM0DS_INST/u_logic/Rkgvx4 ), .ip2(n6265), .op(
        n6266) );
  nand3_1 U7438 ( .ip1(n9634), .ip2(n8823), .ip3(n2140), .op(n6276) );
  and2_1 U7439 ( .ip1(n6276), .ip2(\CORTEXM0DS_INST/u_logic/I4gvx4 ), .op(
        n6946) );
  nor2_1 U7440 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n12095), .op(
        n11202) );
  nor2_1 U7441 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n10865), .op(
        n11207) );
  inv_1 U7442 ( .ip(n11207), .op(n12651) );
  nor2_1 U7443 ( .ip1(n12096), .ip2(n12651), .op(n10819) );
  or2_1 U7444 ( .ip1(n11202), .ip2(n10819), .op(n6271) );
  or2_1 U7445 ( .ip1(n10830), .ip2(n10819), .op(n6270) );
  nand2_1 U7446 ( .ip1(n6271), .ip2(n6270), .op(n11016) );
  inv_1 U7447 ( .ip(n11016), .op(n6272) );
  nand2_1 U7448 ( .ip1(n2140), .ip2(n6272), .op(n12089) );
  inv_1 U7449 ( .ip(n12089), .op(n12641) );
  nor2_1 U7450 ( .ip1(n6946), .ip2(n12641), .op(n6273) );
  or2_1 U7451 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n6273), .op(n6275) );
  inv_1 U7452 ( .ip(\CORTEXM0DS_INST/u_logic/Xyfvx4 ), .op(n8538) );
  or2_1 U7453 ( .ip1(n8538), .ip2(n6273), .op(n6274) );
  nand2_1 U7454 ( .ip1(n6275), .ip2(n6274), .op(n6278) );
  nand2_1 U7455 ( .ip1(\CORTEXM0DS_INST/u_logic/A3gvx4 ), .ip2(n6276), .op(
        n12639) );
  nand2_1 U7456 ( .ip1(n12639), .ip2(n12089), .op(n6277) );
  inv_1 U7457 ( .ip(\CORTEXM0DS_INST/vis_pc [0]), .op(n8537) );
  mux2_1 U7458 ( .ip1(n6278), .ip2(n6277), .s(n8537), .op(n6357) );
  nor3_1 U7459 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n10665), .ip3(
        n12651), .op(n6343) );
  nor2_1 U7460 ( .ip1(n12075), .ip2(n10811), .op(n10678) );
  nor2_1 U7461 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Efgvx4 ), .op(n11698) );
  nand4_1 U7462 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n11698), .ip3(
        n11200), .ip4(n11725), .op(n11652) );
  inv_1 U7463 ( .ip(n9781), .op(n6957) );
  inv_1 U7464 ( .ip(\CORTEXM0DS_INST/vis_ipsr [2]), .op(n10980) );
  nand3_1 U7465 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [1]), .ip2(n6957), .ip3(
        n10980), .op(n12646) );
  inv_1 U7466 ( .ip(\CORTEXM0DS_INST/vis_ipsr [0]), .op(n12403) );
  inv_1 U7467 ( .ip(\CORTEXM0DS_INST/vis_ipsr [4]), .op(n6280) );
  nor2_1 U7468 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [5]), .ip2(n6280), .op(n6336)
         );
  nand2_1 U7469 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [3]), .ip2(n6336), .op(n11863) );
  nor4_1 U7470 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [1]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [2]), .ip3(n12403), .ip4(n11863), .op(n8546)
         );
  inv_1 U7471 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [10]), .op(n6281) );
  nor3_1 U7472 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [5]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [3]), .ip3(n6280), .op(n6293) );
  inv_1 U7473 ( .ip(\CORTEXM0DS_INST/vis_ipsr [1]), .op(n10991) );
  nand4_1 U7474 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [2]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [0]), .ip3(n6293), .ip4(n10991), .op(n9787)
         );
  nor2_1 U7475 ( .ip1(n6281), .ip2(n9787), .op(n6283) );
  inv_1 U7476 ( .ip(n6293), .op(n11847) );
  nor3_1 U7477 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [2]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [0]), .ip3(n10991), .op(n6956) );
  inv_1 U7478 ( .ip(n6956), .op(n9782) );
  nor2_1 U7479 ( .ip1(n11847), .ip2(n9782), .op(n8774) );
  and2_1 U7480 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [4]), .ip2(n8774), .op(
        n6282) );
  not_ab_or_c_or_d U7481 ( .ip1(n8546), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [18]), .ip3(n6283), .ip4(n6282), .op(
        n6291) );
  nand3_1 U7482 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [1]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [2]), .ip3(\CORTEXM0DS_INST/vis_ipsr [0]), 
        .op(n11864) );
  nor2_1 U7483 ( .ip1(n11847), .ip2(n11864), .op(n8768) );
  inv_1 U7484 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [24]), .op(n10186) );
  nor4_1 U7485 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [1]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [0]), .ip3(n10980), .ip4(n11863), .op(n6325)
         );
  inv_1 U7486 ( .ip(n6325), .op(n11845) );
  nor2_1 U7487 ( .ip1(n10186), .ip2(n11845), .op(n6285) );
  inv_1 U7488 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [28]), .op(n10202) );
  inv_1 U7489 ( .ip(n11863), .op(n6297) );
  nor3_1 U7490 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [0]), .ip2(n10980), .ip3(
        n10991), .op(n6292) );
  nand2_1 U7491 ( .ip1(n6297), .ip2(n6292), .op(n6313) );
  nor2_1 U7492 ( .ip1(n10202), .ip2(n6313), .op(n6284) );
  not_ab_or_c_or_d U7493 ( .ip1(n8768), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [14]), .ip3(n6285), .ip4(n6284), .op(
        n6290) );
  nand3_1 U7494 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [3]), .ip2(n6300), .ip3(n6292), .op(n6310) );
  inv_1 U7495 ( .ip(n6310), .op(n11859) );
  nor4_1 U7496 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [1]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [2]), .ip3(n12403), .ip4(n11847), .op(n8793)
         );
  and2_1 U7497 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [2]), .ip2(n8793), .op(
        n6287) );
  inv_1 U7498 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [0]), .op(n7223) );
  nor3_1 U7499 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [1]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [2]), .ip3(\CORTEXM0DS_INST/vis_ipsr [0]), 
        .op(n6296) );
  nand2_1 U7500 ( .ip1(n6296), .ip2(n6293), .op(n11843) );
  nor2_1 U7501 ( .ip1(n7223), .ip2(n11843), .op(n6286) );
  not_ab_or_c_or_d U7502 ( .ip1(n11859), .ip2(
        \CORTEXM0DS_INST/u_logic/Psh2z4 [0]), .ip3(n6287), .ip4(n6286), .op(
        n6289) );
  nand3_1 U7503 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [1]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [0]), .ip3(n10980), .op(n11846) );
  nor2_1 U7504 ( .ip1(n11847), .ip2(n11846), .op(n6326) );
  nand2_1 U7505 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [6]), .ip2(n6326), .op(
        n6288) );
  nor4_1 U7506 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [1]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [0]), .ip3(n10980), .ip4(n11847), .op(n8780)
         );
  inv_1 U7507 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [12]), .op(n7201) );
  nand2_1 U7508 ( .ip1(n6293), .ip2(n6292), .op(n11844) );
  nor2_1 U7509 ( .ip1(n7201), .ip2(n11844), .op(n6295) );
  inv_1 U7510 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [20]), .op(n10204) );
  nand2_1 U7511 ( .ip1(n6297), .ip2(n6956), .op(n11857) );
  nor2_1 U7512 ( .ip1(n10204), .ip2(n11857), .op(n6294) );
  not_ab_or_c_or_d U7513 ( .ip1(n8780), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [8]), .ip3(n6295), .ip4(n6294), .op(
        n6304) );
  nor2_1 U7514 ( .ip1(n11863), .ip2(n11846), .op(n6309) );
  inv_1 U7515 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [16]), .op(n7144) );
  nand2_1 U7516 ( .ip1(n6296), .ip2(n6297), .op(n11858) );
  nor2_1 U7517 ( .ip1(n7144), .ip2(n11858), .op(n6299) );
  inv_1 U7518 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [26]), .op(n7169) );
  nand4_1 U7519 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [2]), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [0]), .ip3(n6297), .ip4(n10991), .op(n8543)
         );
  nor2_1 U7520 ( .ip1(n7169), .ip2(n8543), .op(n6298) );
  not_ab_or_c_or_d U7521 ( .ip1(n6309), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [22]), .ip3(n6299), .ip4(n6298), .op(
        n6303) );
  nor2_1 U7522 ( .ip1(n11864), .ip2(n11863), .op(n6308) );
  nand2_1 U7523 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [30]), .ip2(n6308), 
        .op(n6302) );
  inv_1 U7524 ( .ip(n6300), .op(n6321) );
  nor3_1 U7525 ( .ip1(n6322), .ip2(n6321), .ip3(n11864), .op(n12011) );
  nand2_1 U7526 ( .ip1(\CORTEXM0DS_INST/u_logic/Txh2z4 [0]), .ip2(n12011), 
        .op(n6301) );
  nor2_1 U7527 ( .ip1(n8577), .ip2(n8576), .op(n6305) );
  nor2_1 U7528 ( .ip1(\CORTEXM0DS_INST/u_logic/Uth2z4 [0]), .ip2(n6305), .op(
        n6338) );
  inv_1 U7529 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [27]), .op(n7306) );
  nor2_1 U7530 ( .ip1(n7306), .ip2(n8543), .op(n6307) );
  inv_1 U7531 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [13]), .op(n7202) );
  nor2_1 U7532 ( .ip1(n7202), .ip2(n11844), .op(n6306) );
  not_ab_or_c_or_d U7533 ( .ip1(n6308), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [31]), .ip3(n6307), .ip4(n6306), .op(
        n6334) );
  inv_1 U7534 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [21]), .op(n7139) );
  nor2_1 U7535 ( .ip1(n7139), .ip2(n11857), .op(n6318) );
  nand2_1 U7536 ( .ip1(n6309), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [23]), 
        .op(n6316) );
  and2_1 U7537 ( .ip1(\CORTEXM0DS_INST/u_logic/Txh2z4 [1]), .ip2(n12011), .op(
        n6312) );
  inv_1 U7538 ( .ip(\CORTEXM0DS_INST/u_logic/Psh2z4 [1]), .op(n7290) );
  nor2_1 U7539 ( .ip1(n7290), .ip2(n6310), .op(n6311) );
  not_ab_or_c_or_d U7540 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [3]), .ip2(
        n8793), .ip3(n6312), .ip4(n6311), .op(n6315) );
  inv_1 U7541 ( .ip(n6313), .op(n8786) );
  nand2_1 U7542 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [29]), .ip2(n8786), 
        .op(n6314) );
  nand3_1 U7543 ( .ip1(n6316), .ip2(n6315), .ip3(n6314), .op(n6317) );
  not_ab_or_c_or_d U7544 ( .ip1(n8768), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [15]), .ip3(n6318), .ip4(n6317), .op(
        n6333) );
  inv_1 U7545 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [1]), .op(n11796) );
  nor2_1 U7546 ( .ip1(n11796), .ip2(n11843), .op(n6320) );
  inv_1 U7547 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [17]), .op(n11794) );
  nor2_1 U7548 ( .ip1(n11794), .ip2(n11858), .op(n6319) );
  not_ab_or_c_or_d U7549 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [19]), .ip2(
        n8546), .ip3(n6320), .ip4(n6319), .op(n6330) );
  inv_1 U7550 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [11]), .op(n7213) );
  nor2_1 U7551 ( .ip1(n7213), .ip2(n9787), .op(n6324) );
  nor3_1 U7552 ( .ip1(n6322), .ip2(n6321), .ip3(n11846), .op(n11851) );
  and2_1 U7553 ( .ip1(\CORTEXM0DS_INST/u_logic/Uth2z4 [1]), .ip2(n11851), .op(
        n6323) );
  not_ab_or_c_or_d U7554 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [25]), .ip2(
        n6325), .ip3(n6324), .ip4(n6323), .op(n6329) );
  nand2_1 U7555 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [5]), .ip2(n8774), .op(
        n6328) );
  nand2_1 U7556 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [7]), .ip2(n6326), .op(
        n6327) );
  and4_1 U7557 ( .ip1(n6330), .ip2(n6329), .ip3(n6328), .ip4(n6327), .op(n6332) );
  nand2_1 U7558 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [9]), .ip2(n8780), .op(
        n6331) );
  nor2_1 U7559 ( .ip1(n8585), .ip2(n6338), .op(n6335) );
  nor2_1 U7560 ( .ip1(\CORTEXM0DS_INST/u_logic/Uth2z4 [1]), .ip2(n6335), .op(
        n6337) );
  ab_or_c_or_d U7561 ( .ip1(n6338), .ip2(n8585), .ip3(n6337), .ip4(n8588), 
        .op(n6339) );
  inv_1 U7562 ( .ip(\CORTEXM0DS_INST/cm0_primask[0] ), .op(n11477) );
  nand3_1 U7563 ( .ip1(n12646), .ip2(n6339), .ip3(n11477), .op(n11700) );
  nand2_1 U7564 ( .ip1(n6356), .ip2(n6340), .op(n6341) );
  not_ab_or_c_or_d U7565 ( .ip1(n6344), .ip2(n6343), .ip3(n6342), .ip4(n6341), 
        .op(n11658) );
  inv_1 U7566 ( .ip(\CORTEXM0DS_INST/u_logic/Rkgvx4 ), .op(n12647) );
  or2_1 U7567 ( .ip1(n11658), .ip2(n12647), .op(n6347) );
  or2_1 U7568 ( .ip1(n6345), .ip2(n12647), .op(n6346) );
  nand2_1 U7569 ( .ip1(n6347), .ip2(n6346), .op(n6354) );
  nand2_1 U7570 ( .ip1(n10547), .ip2(n10865), .op(n11164) );
  or2_1 U7571 ( .ip1(n11164), .ip2(n9009), .op(n6348) );
  or2_1 U7572 ( .ip1(n6348), .ip2(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .op(n6352) );
  nor3_1 U7573 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip3(n10892), .op(n6439) );
  nor2_1 U7574 ( .ip1(n11730), .ip2(n10652), .op(n6349) );
  nand4_1 U7575 ( .ip1(n6439), .ip2(\CORTEXM0DS_INST/u_logic/Rkgvx4 ), .ip3(
        n6349), .ip4(n11038), .op(n6350) );
  or2_1 U7576 ( .ip1(n6350), .ip2(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .op(n6351) );
  nand2_1 U7577 ( .ip1(n6352), .ip2(n6351), .op(n6353) );
  not_ab_or_c_or_d U7578 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n6355), 
        .ip3(n6354), .ip4(n6353), .op(n6958) );
  nand3_1 U7579 ( .ip1(n6958), .ip2(n6845), .ip3(n6356), .op(n8501) );
  nor2_1 U7580 ( .ip1(n6357), .ip2(n8501), .op(n9826) );
  or2_1 U7581 ( .ip1(n8563), .ip2(n9826), .op(n8796) );
  nor2_1 U7582 ( .ip1(n8564), .ip2(n8796), .op(n9801) );
  nand2_1 U7583 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .op(n10587) );
  nand2_1 U7584 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10949), .op(
        n9664) );
  nor2_1 U7585 ( .ip1(n10587), .ip2(n9664), .op(n11217) );
  nor3_1 U7586 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip3(n11038), .op(n9550) );
  not_ab_or_c_or_d U7587 ( .ip1(n11207), .ip2(n11184), .ip3(n11217), .ip4(
        n9550), .op(n6417) );
  inv_1 U7588 ( .ip(\CORTEXM0DS_INST/u_logic/O8gvx4 ), .op(n9582) );
  or2_1 U7589 ( .ip1(n6417), .ip2(n9582), .op(n6370) );
  inv_1 U7590 ( .ip(n9620), .op(n8419) );
  nor2_1 U7591 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n12625), .op(
        n10899) );
  nor3_1 U7592 ( .ip1(n10587), .ip2(n10771), .ip3(n8986), .op(n6358) );
  or2_1 U7593 ( .ip1(n10899), .ip2(n6358), .op(n6359) );
  nand2_1 U7594 ( .ip1(n6359), .ip2(n11651), .op(n6360) );
  nor2_1 U7595 ( .ip1(n6360), .ip2(n11754), .op(n6367) );
  inv_1 U7596 ( .ip(n11200), .op(n6442) );
  nor2_1 U7597 ( .ip1(n6442), .ip2(n10903), .op(n10531) );
  or2_1 U7598 ( .ip1(\CORTEXM0DS_INST/vis_apsr [1]), .ip2(n10531), .op(n6364)
         );
  nor3_1 U7599 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(n8553), .ip3(
        n11730), .op(n6361) );
  or2_1 U7600 ( .ip1(n6361), .ip2(n9570), .op(n6362) );
  or2_1 U7601 ( .ip1(n6362), .ip2(n10531), .op(n6363) );
  nand2_1 U7602 ( .ip1(n6364), .ip2(n6363), .op(n6365) );
  nor2_1 U7603 ( .ip1(n6365), .ip2(n11038), .op(n6366) );
  not_ab_or_c_or_d U7604 ( .ip1(n10776), .ip2(n8419), .ip3(n6367), .ip4(n6366), 
        .op(n6368) );
  or2_1 U7605 ( .ip1(n6368), .ip2(n9582), .op(n6369) );
  nand2_1 U7606 ( .ip1(n6370), .ip2(n6369), .op(n6838) );
  nor2_1 U7607 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n8553), .op(
        n9520) );
  or2_1 U7608 ( .ip1(n9620), .ip2(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(n6372) );
  or2_1 U7609 ( .ip1(n8623), .ip2(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(n6371) );
  nand2_1 U7610 ( .ip1(n6372), .ip2(n6371), .op(n6373) );
  inv_1 U7611 ( .ip(n12614), .op(n12606) );
  nor2_1 U7612 ( .ip1(n12614), .ip2(n10949), .op(n8554) );
  nor3_1 U7613 ( .ip1(n8456), .ip2(n8554), .ip3(n11164), .op(n6375) );
  or2_1 U7614 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n6375), .op(n6377) );
  nor2_1 U7615 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n6210), .op(
        n10729) );
  nand2_1 U7616 ( .ip1(n10729), .ip2(n11650), .op(n9594) );
  or2_1 U7617 ( .ip1(n9594), .ip2(n6375), .op(n6376) );
  nand2_1 U7618 ( .ip1(n6377), .ip2(n6376), .op(n6378) );
  nor2_1 U7619 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n12613), .op(
        n10864) );
  not_ab_or_c_or_d U7620 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n12606), .ip3(n6378), .ip4(n10864), .op(n6379) );
  nand2_1 U7621 ( .ip1(n6380), .ip2(n6379), .op(n8969) );
  inv_1 U7622 ( .ip(n8969), .op(n8974) );
  nand2_1 U7623 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [1]), .ip2(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [0]), .op(n6395) );
  nand2_1 U7624 ( .ip1(n10495), .ip2(n12338), .op(n12353) );
  nand4_1 U7625 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip3(n11651), .ip4(n12625), .op(
        n6381) );
  nand2_1 U7626 ( .ip1(n12353), .ip2(n6381), .op(n8948) );
  or2_1 U7627 ( .ip1(n11654), .ip2(n10819), .op(n6382) );
  nand2_1 U7628 ( .ip1(n6382), .ip2(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .op(
        n6387) );
  nor2_1 U7629 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n10665), .op(
        n11077) );
  nor2_1 U7630 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n12625), .op(
        n11181) );
  inv_1 U7631 ( .ip(n11181), .op(n11022) );
  nor3_1 U7632 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n12614), .ip3(
        n11022), .op(n6383) );
  not_ab_or_c_or_d U7633 ( .ip1(n11077), .ip2(n12606), .ip3(n12627), .ip4(
        n6383), .op(n6386) );
  nand4_1 U7634 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [1]), .ip2(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [0]), .ip3(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [3]), .ip4(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [2]), .op(n6385) );
  nand3_1 U7635 ( .ip1(n10547), .ip2(n11754), .ip3(n11214), .op(n6384) );
  nand4_1 U7636 ( .ip1(n6387), .ip2(n6386), .ip3(n6385), .ip4(n6384), .op(
        n6389) );
  nor2_1 U7637 ( .ip1(n8948), .ip2(n6389), .op(n8946) );
  inv_1 U7638 ( .ip(\CORTEXM0DS_INST/u_logic/Tjh2z4 [2]), .op(n8756) );
  nand3_1 U7639 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [3]), .ip2(n8946), 
        .ip3(n8756), .op(n6405) );
  nor2_1 U7640 ( .ip1(n6395), .ip2(n6405), .op(n8957) );
  nor3_1 U7641 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [1]), .ip2(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [0]), .ip3(n6405), .op(n8945) );
  and2_1 U7642 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [0]), .op(n6411)
         );
  nand2_1 U7643 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [3]), .ip2(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [2]), .op(n6388) );
  inv_1 U7644 ( .ip(n8946), .op(n8887) );
  or2_1 U7645 ( .ip1(n6388), .ip2(n8887), .op(n6884) );
  inv_1 U7646 ( .ip(\CORTEXM0DS_INST/u_logic/Tjh2z4 [0]), .op(n11158) );
  nand2_1 U7647 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [1]), .ip2(n11158), 
        .op(n6404) );
  nor2_1 U7648 ( .ip1(n6884), .ip2(n6404), .op(n8958) );
  inv_1 U7649 ( .ip(n8948), .op(n12051) );
  nand2_1 U7650 ( .ip1(n6389), .ip2(n12051), .op(n7975) );
  inv_1 U7651 ( .ip(\CORTEXM0DS_INST/u_logic/Kycvx4 ), .op(n12288) );
  nor2_1 U7652 ( .ip1(n7975), .ip2(n12288), .op(n6402) );
  nor3_1 U7653 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [3]), .ip2(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [2]), .ip3(n6404), .op(n6765) );
  nor4_1 U7654 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [1]), .ip2(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [0]), .ip3(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [3]), .ip4(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [2]), .op(n6763) );
  and2_1 U7655 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [0]), .op(n6400)
         );
  inv_1 U7656 ( .ip(\CORTEXM0DS_INST/u_logic/Tjh2z4 [3]), .op(n8720) );
  nand2_1 U7657 ( .ip1(n8720), .ip2(\CORTEXM0DS_INST/u_logic/Tjh2z4 [2]), .op(
        n6390) );
  nor2_1 U7658 ( .ip1(n6395), .ip2(n6390), .op(n6762) );
  nand2_1 U7659 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [0]), .op(n6398)
         );
  nor2_1 U7660 ( .ip1(n6404), .ip2(n6390), .op(n6775) );
  nand2_1 U7661 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [0]), .op(n6394)
         );
  inv_1 U7662 ( .ip(\CORTEXM0DS_INST/u_logic/Tjh2z4 [1]), .op(n8745) );
  nand2_1 U7663 ( .ip1(n8745), .ip2(\CORTEXM0DS_INST/u_logic/Tjh2z4 [0]), .op(
        n6883) );
  nor2_1 U7664 ( .ip1(n6883), .ip2(n6390), .op(n6764) );
  nand2_1 U7665 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [0]), .op(n6393)
         );
  nor3_1 U7666 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [3]), .ip2(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [2]), .ip3(n6883), .op(n6774) );
  nand2_1 U7667 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [0]), .op(n6392)
         );
  nand2_1 U7668 ( .ip1(n8745), .ip2(n11158), .op(n6403) );
  nor2_1 U7669 ( .ip1(n6403), .ip2(n6390), .op(n6766) );
  nand2_1 U7670 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [0]), .op(n6391)
         );
  and4_1 U7671 ( .ip1(n6394), .ip2(n6393), .ip3(n6392), .ip4(n6391), .op(n6397) );
  nor3_1 U7672 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [3]), .ip2(
        \CORTEXM0DS_INST/u_logic/Tjh2z4 [2]), .ip3(n6395), .op(n6767) );
  nand2_1 U7673 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [0]), .op(n6396)
         );
  nand3_1 U7674 ( .ip1(n6398), .ip2(n6397), .ip3(n6396), .op(n6399) );
  not_ab_or_c_or_d U7675 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [0]), 
        .ip3(n6400), .ip4(n6399), .op(n9294) );
  nor2_1 U7676 ( .ip1(n9294), .ip2(n8887), .op(n6401) );
  not_ab_or_c_or_d U7677 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [0]), .ip2(n8958), 
        .ip3(n6402), .ip4(n6401), .op(n6409) );
  nor2_1 U7678 ( .ip1(n6403), .ip2(n6884), .op(n8966) );
  nand2_1 U7679 ( .ip1(n8966), .ip2(\CORTEXM0DS_INST/cm0_r12 [0]), .op(n6408)
         );
  nor2_1 U7680 ( .ip1(n6404), .ip2(n6405), .op(n8944) );
  nand2_1 U7681 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [0]), .op(n6407)
         );
  nor2_1 U7682 ( .ip1(n6405), .ip2(n6883), .op(n8956) );
  nand2_1 U7683 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [0]), .op(n6406)
         );
  not_ab_or_c_or_d U7684 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [0]), .ip2(n8957), 
        .ip3(n6411), .ip4(n6410), .op(n9183) );
  nor2_1 U7685 ( .ip1(n8974), .ip2(n9183), .op(n6833) );
  or2_1 U7686 ( .ip1(n11200), .ip2(n9570), .op(n6413) );
  or2_1 U7687 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n9570), .op(n6412) );
  nand2_1 U7688 ( .ip1(n6413), .ip2(n6412), .op(n6414) );
  or2_1 U7689 ( .ip1(n6414), .ip2(n10587), .op(n6416) );
  nand2_1 U7690 ( .ip1(n11198), .ip2(n6210), .op(n11722) );
  nor2_1 U7691 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(n10865), .op(
        n10705) );
  nand3_1 U7692 ( .ip1(n10705), .ip2(n8553), .ip3(n8993), .op(n6415) );
  nand2_1 U7693 ( .ip1(\CORTEXM0DS_INST/u_logic/O8gvx4 ), .ip2(n7827), .op(
        n8297) );
  inv_1 U7694 ( .ip(n8297), .op(n8013) );
  nand2_1 U7695 ( .ip1(\CORTEXM0DS_INST/u_logic/Vu8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nt8vx4 ), .op(n6846) );
  nor3_1 U7696 ( .ip1(\CORTEXM0DS_INST/u_logic/Fs8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Xq8vx4 ), .ip3(n6846), .op(n8924) );
  nand2_1 U7697 ( .ip1(\CORTEXM0DS_INST/u_logic/Fs8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Xq8vx4 ), .op(n6431) );
  nor2_1 U7698 ( .ip1(n6846), .ip2(n6431), .op(n8853) );
  inv_1 U7699 ( .ip(n8853), .op(n8909) );
  nor2_1 U7700 ( .ip1(n8909), .ip2(n12288), .op(n6438) );
  inv_1 U7701 ( .ip(\CORTEXM0DS_INST/u_logic/Fs8vx4 ), .op(n8666) );
  nand2_1 U7702 ( .ip1(\CORTEXM0DS_INST/u_logic/Xq8vx4 ), .ip2(n8666), .op(
        n6847) );
  inv_1 U7703 ( .ip(\CORTEXM0DS_INST/u_logic/Nt8vx4 ), .op(n8695) );
  nand2_1 U7704 ( .ip1(\CORTEXM0DS_INST/u_logic/Vu8vx4 ), .ip2(n8695), .op(
        n6432) );
  nor2_1 U7705 ( .ip1(n6847), .ip2(n6432), .op(n8933) );
  inv_1 U7706 ( .ip(\CORTEXM0DS_INST/u_logic/Xq8vx4 ), .op(n11160) );
  nand2_1 U7707 ( .ip1(\CORTEXM0DS_INST/u_logic/Fs8vx4 ), .ip2(n11160), .op(
        n6430) );
  nor2_1 U7708 ( .ip1(n6430), .ip2(n6432), .op(n8916) );
  and2_1 U7709 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [0]), .op(n6429)
         );
  nor3_1 U7710 ( .ip1(\CORTEXM0DS_INST/u_logic/Vu8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nt8vx4 ), .ip3(n6430), .op(n8941) );
  nand2_1 U7711 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [0]), .op(n6428)
         );
  nor3_1 U7712 ( .ip1(\CORTEXM0DS_INST/u_logic/Vu8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nt8vx4 ), .ip3(n6847), .op(n8917) );
  nand2_1 U7713 ( .ip1(n8666), .ip2(n11160), .op(n6418) );
  inv_1 U7714 ( .ip(\CORTEXM0DS_INST/u_logic/Vu8vx4 ), .op(n8707) );
  nand2_1 U7715 ( .ip1(n8707), .ip2(\CORTEXM0DS_INST/u_logic/Nt8vx4 ), .op(
        n6419) );
  nor2_1 U7716 ( .ip1(n6418), .ip2(n6419), .op(n8904) );
  and2_1 U7717 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [0]), .op(n6425)
         );
  nor2_1 U7718 ( .ip1(n6431), .ip2(n6419), .op(n8934) );
  nand2_1 U7719 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [0]), .op(n6423)
         );
  nor2_1 U7720 ( .ip1(n6430), .ip2(n6419), .op(n8925) );
  nand2_1 U7721 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [0]), .op(n6422)
         );
  nor2_1 U7722 ( .ip1(n6847), .ip2(n6419), .op(n8903) );
  nand2_1 U7723 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [0]), .op(n6421)
         );
  nor4_1 U7724 ( .ip1(\CORTEXM0DS_INST/u_logic/Vu8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nt8vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Fs8vx4 ), .ip4(
        \CORTEXM0DS_INST/u_logic/Xq8vx4 ), .op(n8932) );
  nand2_1 U7725 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [0]), .op(n6420)
         );
  not_ab_or_c_or_d U7726 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [0]), .ip2(n8917), 
        .ip3(n6425), .ip4(n6424), .op(n6427) );
  nor3_1 U7727 ( .ip1(\CORTEXM0DS_INST/u_logic/Vu8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nt8vx4 ), .ip3(n6431), .op(n8915) );
  nand2_1 U7728 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [0]), .op(n6426)
         );
  nand3_1 U7729 ( .ip1(n6428), .ip2(n6427), .ip3(n6426), .op(n6971) );
  not_ab_or_c_or_d U7730 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [0]), 
        .ip3(n6429), .ip4(n6971), .op(n6436) );
  nor2_1 U7731 ( .ip1(n6430), .ip2(n6846), .op(n8910) );
  nand2_1 U7732 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [0]), .op(n6435)
         );
  nor2_1 U7733 ( .ip1(n6432), .ip2(n6431), .op(n8914) );
  nand2_1 U7734 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [0]), .op(n6434)
         );
  nor3_1 U7735 ( .ip1(\CORTEXM0DS_INST/u_logic/Fs8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Xq8vx4 ), .ip3(n6432), .op(n8902) );
  nand2_1 U7736 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [0]), .op(n6433)
         );
  not_ab_or_c_or_d U7737 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [0]), 
        .ip3(n6438), .ip4(n6437), .op(n8598) );
  nand2_1 U7738 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10865), .op(
        n11183) );
  nor2_1 U7739 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n10865), .op(
        n11186) );
  not_ab_or_c_or_d U7740 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n11183), .ip3(n6439), .ip4(n11186), .op(n6440) );
  nor2_1 U7741 ( .ip1(n6440), .ip2(n11754), .op(n6441) );
  not_ab_or_c_or_d U7742 ( .ip1(n10880), .ip2(n10937), .ip3(n10705), .ip4(
        n6441), .op(n6445) );
  nor2_1 U7743 ( .ip1(n11730), .ip2(n6442), .op(n9748) );
  nand3_1 U7744 ( .ip1(n11202), .ip2(n9748), .ip3(n11754), .op(n6444) );
  nand3_1 U7745 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n9598), .ip3(
        n8495), .op(n6443) );
  nand2_1 U7746 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n11715), .op(
        n8616) );
  nand4_1 U7747 ( .ip1(n6445), .ip2(n6444), .ip3(n6443), .ip4(n8616), .op(
        n6446) );
  nand2_1 U7748 ( .ip1(\CORTEXM0DS_INST/u_logic/O8gvx4 ), .ip2(n6446), .op(
        n8292) );
  nor2_1 U7749 ( .ip1(n8598), .ip2(n8292), .op(n6455) );
  or2_1 U7750 ( .ip1(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip2(n6455), .op(n6457) );
  nand4_1 U7751 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/O8gvx4 ), .ip4(n9639), .op(n7823) );
  inv_1 U7752 ( .ip(n7823), .op(n7575) );
  nor2_1 U7753 ( .ip1(n11754), .ip2(n12095), .op(n12334) );
  or2_1 U7754 ( .ip1(n11181), .ip2(n12334), .op(n6448) );
  or2_1 U7755 ( .ip1(n11730), .ip2(n12334), .op(n6447) );
  nand2_1 U7756 ( .ip1(n6448), .ip2(n6447), .op(n6449) );
  nor2_1 U7757 ( .ip1(n6449), .ip2(n11038), .op(n6452) );
  not_ab_or_c_or_d U7758 ( .ip1(n8996), .ip2(n8623), .ip3(
        \CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip4(n12095), .op(n6451) );
  nand2_1 U7759 ( .ip1(n10949), .ip2(n12625), .op(n8474) );
  nand2_1 U7760 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n6210), .op(
        n10676) );
  not_ab_or_c_or_d U7761 ( .ip1(n8474), .ip2(n10676), .ip3(n12095), .ip4(
        n10547), .op(n6450) );
  nor2_1 U7762 ( .ip1(n6453), .ip2(n9582), .op(n7670) );
  nor4_1 U7763 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip3(n10587), .ip4(n10771), .op(
        n11714) );
  and2_1 U7764 ( .ip1(\CORTEXM0DS_INST/u_logic/O8gvx4 ), .ip2(n11714), .op(
        n6454) );
  nor2_1 U7765 ( .ip1(n7670), .ip2(n6454), .op(n6829) );
  inv_1 U7766 ( .ip(n6829), .op(n6914) );
  or2_1 U7767 ( .ip1(n6914), .ip2(n6455), .op(n6456) );
  nand2_1 U7768 ( .ip1(n6457), .ip2(n6456), .op(n6458) );
  mux2_1 U7769 ( .ip1(n8297), .ip2(n8013), .s(n6458), .op(n9181) );
  xor2_1 U7770 ( .ip1(n6833), .ip2(n9181), .op(n6839) );
  xor2_1 U7771 ( .ip1(n6838), .ip2(n6839), .op(n11476) );
  inv_1 U7772 ( .ip(n11476), .op(n11018) );
  inv_1 U7773 ( .ip(n12305), .op(n12599) );
  nand2_1 U7774 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n11730), .op(
        n10976) );
  nand2_1 U7775 ( .ip1(n10976), .ip2(n8623), .op(n6794) );
  inv_1 U7776 ( .ip(n11164), .op(n11661) );
  nor3_1 U7777 ( .ip1(n11661), .ip2(n11169), .ip3(n11754), .op(n6793) );
  inv_1 U7778 ( .ip(n11168), .op(n6459) );
  inv_1 U7779 ( .ip(n12603), .op(n9584) );
  not_ab_or_c_or_d U7780 ( .ip1(n12628), .ip2(n6459), .ip3(n9584), .ip4(n10949), .op(n6791) );
  inv_1 U7781 ( .ip(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .op(n11145) );
  nor2_1 U7782 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n11145), .op(
        n11120) );
  and2_1 U7783 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [31]), .ip2(n6766), .op(n6468)
         );
  nand2_1 U7784 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [31]), .op(n6466)
         );
  nand2_1 U7785 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [31]), .ip2(n6764), .op(n6463)
         );
  nand2_1 U7786 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [31]), .ip2(n6775), .op(n6462)
         );
  nand2_1 U7787 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [31]), .ip2(n6765), .op(n6461)
         );
  nand2_1 U7788 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [31]), .ip2(n6763), .op(n6460)
         );
  and4_1 U7789 ( .ip1(n6463), .ip2(n6462), .ip3(n6461), .ip4(n6460), .op(n6465) );
  nand2_1 U7790 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [31]), .ip2(n6774), .op(n6464)
         );
  nand3_1 U7791 ( .ip1(n6466), .ip2(n6465), .ip3(n6464), .op(n6467) );
  not_ab_or_c_or_d U7792 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [31]), .ip2(n6767), 
        .ip3(n6468), .ip4(n6467), .op(n8832) );
  inv_1 U7793 ( .ip(n8832), .op(n9329) );
  nand2_1 U7794 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [29]), .ip2(n6764), .op(n6477)
         );
  and2_1 U7795 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [29]), .op(n6474)
         );
  nand2_1 U7796 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [29]), .op(n6472)
         );
  nand2_1 U7797 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [29]), .op(n6471)
         );
  nand2_1 U7798 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [29]), .op(n6470)
         );
  nand2_1 U7799 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [29]), .op(n6469)
         );
  not_ab_or_c_or_d U7800 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [29]), 
        .ip3(n6474), .ip4(n6473), .op(n6476) );
  nand2_1 U7801 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [29]), .op(n6475)
         );
  nand3_1 U7802 ( .ip1(n6477), .ip2(n6476), .ip3(n6475), .op(n9304) );
  inv_1 U7803 ( .ip(n9304), .op(n9320) );
  nand2_1 U7804 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Ik9vx4 ), .op(n11105) );
  nor2_1 U7805 ( .ip1(n9320), .ip2(n11105), .op(n6489) );
  and2_1 U7806 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [30]), .op(n6486)
         );
  nand2_1 U7807 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [30]), .op(n6484)
         );
  nand2_1 U7808 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [30]), .op(n6481)
         );
  nand2_1 U7809 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [30]), .op(n6480)
         );
  nand2_1 U7810 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [30]), .op(n6479)
         );
  nand2_1 U7811 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [30]), .op(n6478)
         );
  and4_1 U7812 ( .ip1(n6481), .ip2(n6480), .ip3(n6479), .ip4(n6478), .op(n6483) );
  nand2_1 U7813 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [30]), .op(n6482)
         );
  nand3_1 U7814 ( .ip1(n6484), .ip2(n6483), .ip3(n6482), .op(n6485) );
  not_ab_or_c_or_d U7815 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [30]), 
        .ip3(n6486), .ip4(n6485), .op(n8888) );
  inv_1 U7816 ( .ip(n9294), .op(n9331) );
  nor2_1 U7817 ( .ip1(n9331), .ip2(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .op(
        n6487) );
  not_ab_or_c_or_d U7818 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n8888), 
        .ip3(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip4(n6487), .op(n6488) );
  not_ab_or_c_or_d U7819 ( .ip1(n11120), .ip2(n9329), .ip3(n6489), .ip4(n6488), 
        .op(n6530) );
  nand2_1 U7820 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [23]), .ip2(n6775), .op(n6498)
         );
  and2_1 U7821 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [23]), .op(n6495)
         );
  nand2_1 U7822 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [23]), .op(n6493)
         );
  nand2_1 U7823 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [23]), .op(n6492)
         );
  nand2_1 U7824 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [23]), .op(n6491)
         );
  nand2_1 U7825 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [23]), .op(n6490)
         );
  not_ab_or_c_or_d U7826 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [23]), .ip2(n6766), 
        .ip3(n6495), .ip4(n6494), .op(n6497) );
  nand2_1 U7827 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [23]), .op(n6496)
         );
  nand3_1 U7828 ( .ip1(n6498), .ip2(n6497), .ip3(n6496), .op(n9403) );
  and2_1 U7829 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [21]), .op(n6507)
         );
  nand2_1 U7830 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [21]), .op(n6505)
         );
  nand2_1 U7831 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [21]), .op(n6502)
         );
  nand2_1 U7832 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [21]), .op(n6501)
         );
  nand2_1 U7833 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [21]), .op(n6500)
         );
  nand2_1 U7834 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [21]), .op(n6499)
         );
  and4_1 U7835 ( .ip1(n6502), .ip2(n6501), .ip3(n6500), .ip4(n6499), .op(n6504) );
  nand2_1 U7836 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [21]), .op(n6503)
         );
  nand3_1 U7837 ( .ip1(n6505), .ip2(n6504), .ip3(n6503), .op(n6506) );
  not_ab_or_c_or_d U7838 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [21]), 
        .ip3(n6507), .ip4(n6506), .op(n7774) );
  nor2_1 U7839 ( .ip1(n7774), .ip2(n11105), .op(n6528) );
  and2_1 U7840 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [22]), .op(n6516)
         );
  nand2_1 U7841 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [22]), .op(n6514)
         );
  nand2_1 U7842 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [22]), .op(n6511)
         );
  nand2_1 U7843 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [22]), .op(n6510)
         );
  nand2_1 U7844 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [22]), .op(n6509)
         );
  nand2_1 U7845 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [22]), .op(n6508)
         );
  and4_1 U7846 ( .ip1(n6511), .ip2(n6510), .ip3(n6509), .ip4(n6508), .op(n6513) );
  nand2_1 U7847 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [22]), .op(n6512)
         );
  nand3_1 U7848 ( .ip1(n6514), .ip2(n6513), .ip3(n6512), .op(n6515) );
  not_ab_or_c_or_d U7849 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [22]), 
        .ip3(n6516), .ip4(n6515), .op(n8014) );
  nand2_1 U7850 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [24]), .ip2(n6774), .op(n6525)
         );
  and2_1 U7851 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [24]), .op(n6522)
         );
  nand2_1 U7852 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [24]), .op(n6520)
         );
  nand2_1 U7853 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [24]), .op(n6519)
         );
  nand2_1 U7854 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [24]), .op(n6518)
         );
  nand2_1 U7855 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [24]), .op(n6517)
         );
  not_ab_or_c_or_d U7856 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [24]), 
        .ip3(n6522), .ip4(n6521), .op(n6524) );
  nand2_1 U7857 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [24]), .op(n6523)
         );
  nand3_1 U7858 ( .ip1(n6525), .ip2(n6524), .ip3(n6523), .op(n9402) );
  nor2_1 U7859 ( .ip1(n9402), .ip2(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .op(
        n6526) );
  not_ab_or_c_or_d U7860 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n8014), 
        .ip3(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip4(n6526), .op(n6527) );
  not_ab_or_c_or_d U7861 ( .ip1(n11120), .ip2(n9403), .ip3(n6528), .ip4(n6527), 
        .op(n6529) );
  mux2_1 U7862 ( .ip1(n6530), .ip2(n6529), .s(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .op(n6789) );
  nor2_1 U7863 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Qm9vx4 ), .op(n11008) );
  nor2_1 U7864 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Ik9vx4 ), .op(n7055) );
  nand2_1 U7865 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [8]), .op(n6539)
         );
  and2_1 U7866 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [8]), .op(n6536)
         );
  nand2_1 U7867 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [8]), .op(n6534)
         );
  nand2_1 U7868 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [8]), .op(n6533)
         );
  nand2_1 U7869 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [8]), .op(n6532)
         );
  nand2_1 U7870 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [8]), .op(n6531)
         );
  not_ab_or_c_or_d U7871 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [8]), .ip2(n6762), 
        .ip3(n6536), .ip4(n6535), .op(n6538) );
  nand2_1 U7872 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [8]), .op(n6537)
         );
  nand3_1 U7873 ( .ip1(n6539), .ip2(n6538), .ip3(n6537), .op(n9283) );
  nand2_1 U7874 ( .ip1(n7055), .ip2(n9283), .op(n6570) );
  nand2_1 U7875 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [7]), .ip2(n6767), .op(n6548)
         );
  and2_1 U7876 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [7]), .op(n6545)
         );
  nand2_1 U7877 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [7]), .op(n6543)
         );
  nand2_1 U7878 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [7]), .op(n6542)
         );
  nand2_1 U7879 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [7]), .op(n6541)
         );
  nand2_1 U7880 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [7]), .op(n6540)
         );
  not_ab_or_c_or_d U7881 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [7]), 
        .ip3(n6545), .ip4(n6544), .op(n6547) );
  nand2_1 U7882 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [7]), .op(n6546)
         );
  nand3_1 U7883 ( .ip1(n6548), .ip2(n6547), .ip3(n6546), .op(n9281) );
  nand2_1 U7884 ( .ip1(n11120), .ip2(n9281), .op(n6569) );
  inv_1 U7885 ( .ip(n11105), .op(n11073) );
  nand2_1 U7886 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [5]), .op(n6557)
         );
  and2_1 U7887 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [5]), .op(n6554)
         );
  nand2_1 U7888 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [5]), .op(n6552)
         );
  nand2_1 U7889 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [5]), .op(n6551)
         );
  nand2_1 U7890 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [5]), .op(n6550)
         );
  nand2_1 U7891 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [5]), .op(n6549)
         );
  not_ab_or_c_or_d U7892 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [5]), .ip2(n6764), 
        .ip3(n6554), .ip4(n6553), .op(n6556) );
  nand2_1 U7893 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [5]), .op(n6555)
         );
  nand3_1 U7894 ( .ip1(n6557), .ip2(n6556), .ip3(n6555), .op(n9263) );
  nand2_1 U7895 ( .ip1(n11073), .ip2(n9263), .op(n6568) );
  inv_1 U7896 ( .ip(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .op(n6965) );
  nor2_1 U7897 ( .ip1(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip2(n6965), .op(
        n6662) );
  nand2_1 U7898 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [6]), .op(n6566)
         );
  and2_1 U7899 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [6]), .op(n6563)
         );
  nand2_1 U7900 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [6]), .op(n6561)
         );
  nand2_1 U7901 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [6]), .op(n6560)
         );
  nand2_1 U7902 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [6]), .op(n6559)
         );
  nand2_1 U7903 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [6]), .op(n6558)
         );
  not_ab_or_c_or_d U7904 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [6]), 
        .ip3(n6563), .ip4(n6562), .op(n6565) );
  nand2_1 U7905 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [6]), .op(n6564)
         );
  nand3_1 U7906 ( .ip1(n6566), .ip2(n6565), .ip3(n6564), .op(n9282) );
  nand2_1 U7907 ( .ip1(n6662), .ip2(n9282), .op(n6567) );
  nand2_1 U7908 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [15]), .ip2(n6766), .op(n6579)
         );
  and2_1 U7909 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [15]), .op(n6576)
         );
  nand2_1 U7910 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [15]), .op(n6574)
         );
  nand2_1 U7911 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [15]), .op(n6573)
         );
  nand2_1 U7912 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [15]), .op(n6572)
         );
  nand2_1 U7913 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [15]), .op(n6571)
         );
  not_ab_or_c_or_d U7914 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [15]), .ip2(n6775), 
        .ip3(n6576), .ip4(n6575), .op(n6578) );
  nand2_1 U7915 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [15]), .op(n6577)
         );
  nand3_1 U7916 ( .ip1(n6579), .ip2(n6578), .ip3(n6577), .op(n9428) );
  and2_1 U7917 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [13]), .op(n6588)
         );
  nand2_1 U7918 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [13]), .op(n6586)
         );
  nand2_1 U7919 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [13]), .op(n6583)
         );
  nand2_1 U7920 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [13]), .op(n6582)
         );
  nand2_1 U7921 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [13]), .op(n6581)
         );
  nand2_1 U7922 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [13]), .op(n6580)
         );
  and4_1 U7923 ( .ip1(n6583), .ip2(n6582), .ip3(n6581), .ip4(n6580), .op(n6585) );
  nand2_1 U7924 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [13]), .op(n6584)
         );
  nand3_1 U7925 ( .ip1(n6586), .ip2(n6585), .ip3(n6584), .op(n6587) );
  not_ab_or_c_or_d U7926 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [13]), 
        .ip3(n6588), .ip4(n6587), .op(n9417) );
  nor2_1 U7927 ( .ip1(n9417), .ip2(n11105), .op(n6609) );
  and2_1 U7928 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [14]), .op(n6597)
         );
  nand2_1 U7929 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [14]), .ip2(n6762), .op(n6595)
         );
  nand2_1 U7930 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [14]), .op(n6592)
         );
  nand2_1 U7931 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [14]), .op(n6591)
         );
  nand2_1 U7932 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [14]), .op(n6590)
         );
  nand2_1 U7933 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [14]), .op(n6589)
         );
  and4_1 U7934 ( .ip1(n6592), .ip2(n6591), .ip3(n6590), .ip4(n6589), .op(n6594) );
  nand2_1 U7935 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [14]), .op(n6593)
         );
  nand3_1 U7936 ( .ip1(n6595), .ip2(n6594), .ip3(n6593), .op(n6596) );
  not_ab_or_c_or_d U7937 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [14]), .ip2(n6765), 
        .ip3(n6597), .ip4(n6596), .op(n9419) );
  nand2_1 U7938 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [16]), .ip2(n6767), .op(n6606)
         );
  and2_1 U7939 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [16]), .op(n6603)
         );
  nand2_1 U7940 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [16]), .op(n6601)
         );
  nand2_1 U7941 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [16]), .op(n6600)
         );
  nand2_1 U7942 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [16]), .op(n6599)
         );
  nand2_1 U7943 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [16]), .op(n6598)
         );
  not_ab_or_c_or_d U7944 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [16]), 
        .ip3(n6603), .ip4(n6602), .op(n6605) );
  nand2_1 U7945 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [16]), .op(n6604)
         );
  nand3_1 U7946 ( .ip1(n6606), .ip2(n6605), .ip3(n6604), .op(n9432) );
  nor2_1 U7947 ( .ip1(n9432), .ip2(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .op(
        n6607) );
  not_ab_or_c_or_d U7948 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n9419), 
        .ip3(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip4(n6607), .op(n6608) );
  not_ab_or_c_or_d U7949 ( .ip1(n11120), .ip2(n9428), .ip3(n6609), .ip4(n6608), 
        .op(n6610) );
  nor2_1 U7950 ( .ip1(n6610), .ip2(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .op(
        n6611) );
  inv_1 U7951 ( .ip(\CORTEXM0DS_INST/u_logic/Qm9vx4 ), .op(n10891) );
  nand2_1 U7952 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(n10891), .op(
        n11479) );
  not_ab_or_c_or_d U7953 ( .ip1(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .ip2(n6612), 
        .ip3(n6611), .ip4(n11479), .op(n6788) );
  nand2_1 U7954 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [12]), .ip2(n6767), .op(n6621)
         );
  and2_1 U7955 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [12]), .op(n6618)
         );
  nand2_1 U7956 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [12]), .op(n6616)
         );
  nand2_1 U7957 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [12]), .op(n6615)
         );
  nand2_1 U7958 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [12]), .op(n6614)
         );
  nand2_1 U7959 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [12]), .op(n6613)
         );
  not_ab_or_c_or_d U7960 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [12]), .ip2(n6774), 
        .ip3(n6618), .ip4(n6617), .op(n6620) );
  nand2_1 U7961 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [12]), .op(n6619)
         );
  nand3_1 U7962 ( .ip1(n6621), .ip2(n6620), .ip3(n6619), .op(n9269) );
  nand2_1 U7963 ( .ip1(n7055), .ip2(n9269), .op(n6652) );
  nand2_1 U7964 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [9]), .ip2(n6766), .op(n6630)
         );
  and2_1 U7965 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [9]), .op(n6627)
         );
  nand2_1 U7966 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [9]), .op(n6625)
         );
  nand2_1 U7967 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [9]), .op(n6624)
         );
  nand2_1 U7968 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [9]), .op(n6623)
         );
  nand2_1 U7969 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [9]), .op(n6622)
         );
  not_ab_or_c_or_d U7970 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [9]), 
        .ip3(n6627), .ip4(n6626), .op(n6629) );
  nand2_1 U7971 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [9]), .op(n6628)
         );
  nand3_1 U7972 ( .ip1(n6630), .ip2(n6629), .ip3(n6628), .op(n9284) );
  nand2_1 U7973 ( .ip1(n11073), .ip2(n9284), .op(n6651) );
  nand2_1 U7974 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [10]), .ip2(n6766), .op(n6639)
         );
  and2_1 U7975 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [10]), .op(n6636)
         );
  nand2_1 U7976 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [10]), .op(n6634)
         );
  nand2_1 U7977 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [10]), .op(n6633)
         );
  nand2_1 U7978 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [10]), .op(n6632)
         );
  nand2_1 U7979 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [10]), .op(n6631)
         );
  not_ab_or_c_or_d U7980 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [10]), 
        .ip3(n6636), .ip4(n6635), .op(n6638) );
  nand2_1 U7981 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [10]), .op(n6637)
         );
  nand3_1 U7982 ( .ip1(n6639), .ip2(n6638), .ip3(n6637), .op(n9275) );
  nand2_1 U7983 ( .ip1(n6662), .ip2(n9275), .op(n6650) );
  nand2_1 U7984 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [11]), .ip2(n6774), .op(n6648)
         );
  and2_1 U7985 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [11]), .op(n6645)
         );
  nand2_1 U7986 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [11]), .op(n6643)
         );
  nand2_1 U7987 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [11]), .op(n6642)
         );
  nand2_1 U7988 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [11]), .op(n6641)
         );
  nand2_1 U7989 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [11]), .op(n6640)
         );
  not_ab_or_c_or_d U7990 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [11]), .ip2(n6767), 
        .ip3(n6645), .ip4(n6644), .op(n6647) );
  nand2_1 U7991 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [11]), .op(n6646)
         );
  nand3_1 U7992 ( .ip1(n6648), .ip2(n6647), .ip3(n6646), .op(n9276) );
  nand2_1 U7993 ( .ip1(n11120), .ip2(n9276), .op(n6649) );
  nand2_1 U7994 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [2]), .ip2(n6762), .op(n6661)
         );
  and2_1 U7995 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [2]), .op(n6658)
         );
  nand2_1 U7996 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [2]), .op(n6656)
         );
  nand2_1 U7997 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [2]), .op(n6655)
         );
  nand2_1 U7998 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [2]), .op(n6654)
         );
  nand2_1 U7999 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [2]), .op(n6653)
         );
  not_ab_or_c_or_d U8000 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [2]), 
        .ip3(n6658), .ip4(n6657), .op(n6660) );
  nand2_1 U8001 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [2]), .op(n6659)
         );
  nand3_1 U8002 ( .ip1(n6661), .ip2(n6660), .ip3(n6659), .op(n7100) );
  nand2_1 U8003 ( .ip1(n6662), .ip2(n7100), .op(n6693) );
  nand2_1 U8004 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [4]), .op(n6671)
         );
  and2_1 U8005 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [4]), .op(n6668)
         );
  nand2_1 U8006 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [4]), .op(n6666)
         );
  nand2_1 U8007 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [4]), .op(n6665)
         );
  nand2_1 U8008 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [4]), .op(n6664)
         );
  nand2_1 U8009 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [4]), .op(n6663)
         );
  not_ab_or_c_or_d U8010 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [4]), .ip2(n6765), 
        .ip3(n6668), .ip4(n6667), .op(n6670) );
  nand2_1 U8011 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [4]), .op(n6669)
         );
  nand3_1 U8012 ( .ip1(n6671), .ip2(n6670), .ip3(n6669), .op(n9264) );
  nand2_1 U8013 ( .ip1(n7055), .ip2(n9264), .op(n6692) );
  nand2_1 U8014 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [3]), .op(n6680)
         );
  and2_1 U8015 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [3]), .op(n6677)
         );
  nand2_1 U8016 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [3]), .op(n6675)
         );
  nand2_1 U8017 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [3]), .op(n6674)
         );
  nand2_1 U8018 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [3]), .op(n6673)
         );
  nand2_1 U8019 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [3]), .op(n6672)
         );
  not_ab_or_c_or_d U8020 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [3]), .ip2(n6767), 
        .ip3(n6677), .ip4(n6676), .op(n6679) );
  nand2_1 U8021 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [3]), .op(n6678)
         );
  nand3_1 U8022 ( .ip1(n6680), .ip2(n6679), .ip3(n6678), .op(n6976) );
  nand2_1 U8023 ( .ip1(n11120), .ip2(n6976), .op(n6691) );
  nand2_1 U8024 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [1]), .ip2(n6774), .op(n6689)
         );
  and2_1 U8025 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [1]), .op(n6686)
         );
  nand2_1 U8026 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [1]), .op(n6684)
         );
  nand2_1 U8027 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [1]), .op(n6683)
         );
  nand2_1 U8028 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [1]), .op(n6682)
         );
  nand2_1 U8029 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [1]), .op(n6681)
         );
  not_ab_or_c_or_d U8030 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [1]), 
        .ip3(n6686), .ip4(n6685), .op(n6688) );
  nand2_1 U8031 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [1]), .op(n6687)
         );
  nand3_1 U8032 ( .ip1(n6689), .ip2(n6688), .ip3(n6687), .op(n9332) );
  nand2_1 U8033 ( .ip1(n11073), .ip2(n9332), .op(n6690) );
  mux2_1 U8034 ( .ip1(n6695), .ip2(n6694), .s(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .op(n6786) );
  and2_1 U8035 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [27]), .op(n6704)
         );
  nand2_1 U8036 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [27]), .ip2(n6762), .op(n6702)
         );
  nand2_1 U8037 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [27]), .op(n6699)
         );
  nand2_1 U8038 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [27]), .op(n6698)
         );
  nand2_1 U8039 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [27]), .op(n6697)
         );
  nand2_1 U8040 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [27]), .op(n6696)
         );
  and4_1 U8041 ( .ip1(n6699), .ip2(n6698), .ip3(n6697), .ip4(n6696), .op(n6701) );
  nand2_1 U8042 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [27]), .op(n6700)
         );
  nand3_1 U8043 ( .ip1(n6702), .ip2(n6701), .ip3(n6700), .op(n6703) );
  not_ab_or_c_or_d U8044 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [27]), .ip2(n6774), 
        .ip3(n6704), .ip4(n6703), .op(n9319) );
  inv_1 U8045 ( .ip(n9319), .op(n9351) );
  and2_1 U8046 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [25]), .op(n6713)
         );
  nand2_1 U8047 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [25]), .op(n6711)
         );
  nand2_1 U8048 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [25]), .op(n6708)
         );
  nand2_1 U8049 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [25]), .op(n6707)
         );
  nand2_1 U8050 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [25]), .op(n6706)
         );
  nand2_1 U8051 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [25]), .op(n6705)
         );
  and4_1 U8052 ( .ip1(n6708), .ip2(n6707), .ip3(n6706), .ip4(n6705), .op(n6710) );
  nand2_1 U8053 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [25]), .op(n6709)
         );
  nand3_1 U8054 ( .ip1(n6711), .ip2(n6710), .ip3(n6709), .op(n6712) );
  not_ab_or_c_or_d U8055 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [25]), 
        .ip3(n6713), .ip4(n6712), .op(n9350) );
  nor2_1 U8056 ( .ip1(n9350), .ip2(n11105), .op(n6734) );
  nand2_1 U8057 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [26]), .op(n6722)
         );
  and2_1 U8058 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [26]), .op(n6719)
         );
  nand2_1 U8059 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [26]), .op(n6717)
         );
  nand2_1 U8060 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [26]), .op(n6716)
         );
  nand2_1 U8061 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [26]), .op(n6715)
         );
  nand2_1 U8062 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [26]), .op(n6714)
         );
  not_ab_or_c_or_d U8063 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [26]), 
        .ip3(n6719), .ip4(n6718), .op(n6721) );
  nand2_1 U8064 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [26]), .op(n6720)
         );
  nand3_1 U8065 ( .ip1(n6722), .ip2(n6721), .ip3(n6720), .op(n9377) );
  inv_1 U8066 ( .ip(n9377), .op(n9318) );
  and2_1 U8067 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [28]), .op(n6731)
         );
  nand2_1 U8068 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [28]), .op(n6729)
         );
  nand2_1 U8069 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [28]), .op(n6726)
         );
  nand2_1 U8070 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [28]), .op(n6725)
         );
  nand2_1 U8071 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [28]), .op(n6724)
         );
  nand2_1 U8072 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [28]), .op(n6723)
         );
  and4_1 U8073 ( .ip1(n6726), .ip2(n6725), .ip3(n6724), .ip4(n6723), .op(n6728) );
  nand2_1 U8074 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [28]), .op(n6727)
         );
  nand3_1 U8075 ( .ip1(n6729), .ip2(n6728), .ip3(n6727), .op(n6730) );
  not_ab_or_c_or_d U8076 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [28]), 
        .ip3(n6731), .ip4(n6730), .op(n9317) );
  inv_1 U8077 ( .ip(n9317), .op(n9303) );
  nor2_1 U8078 ( .ip1(n9303), .ip2(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .op(
        n6732) );
  not_ab_or_c_or_d U8079 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n9318), 
        .ip3(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip4(n6732), .op(n6733) );
  not_ab_or_c_or_d U8080 ( .ip1(n11120), .ip2(n9351), .ip3(n6734), .ip4(n6733), 
        .op(n6783) );
  nand2_1 U8081 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [19]), .op(n6743)
         );
  and2_1 U8082 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [19]), .op(n6740)
         );
  nand2_1 U8083 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [19]), .op(n6738)
         );
  nand2_1 U8084 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [19]), .op(n6737)
         );
  nand2_1 U8085 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [19]), .op(n6736)
         );
  nand2_1 U8086 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [19]), .op(n6735)
         );
  not_ab_or_c_or_d U8087 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [19]), .ip2(n6764), 
        .ip3(n6740), .ip4(n6739), .op(n6742) );
  nand2_1 U8088 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [19]), .op(n6741)
         );
  nand3_1 U8089 ( .ip1(n6743), .ip2(n6742), .ip3(n6741), .op(n9369) );
  and2_1 U8090 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [17]), .op(n6752)
         );
  nand2_1 U8091 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [17]), .ip2(n6762), .op(n6750)
         );
  nand2_1 U8092 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [17]), .op(n6747)
         );
  nand2_1 U8093 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [17]), .op(n6746)
         );
  nand2_1 U8094 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [17]), .op(n6745)
         );
  nand2_1 U8095 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [17]), .op(n6744)
         );
  and4_1 U8096 ( .ip1(n6747), .ip2(n6746), .ip3(n6745), .ip4(n6744), .op(n6749) );
  nand2_1 U8097 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [17]), .op(n6748)
         );
  nand3_1 U8098 ( .ip1(n6750), .ip2(n6749), .ip3(n6748), .op(n6751) );
  not_ab_or_c_or_d U8099 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [17]), 
        .ip3(n6752), .ip4(n6751), .op(n9389) );
  nor2_1 U8100 ( .ip1(n9389), .ip2(n11105), .op(n6781) );
  and2_1 U8101 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [18]), .op(n6761)
         );
  nand2_1 U8102 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [18]), .op(n6759)
         );
  nand2_1 U8103 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [18]), .op(n6756)
         );
  nand2_1 U8104 ( .ip1(n6762), .ip2(\CORTEXM0DS_INST/cm0_r07 [18]), .op(n6755)
         );
  nand2_1 U8105 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [18]), .op(n6754)
         );
  nand2_1 U8106 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [18]), .op(n6753)
         );
  and4_1 U8107 ( .ip1(n6756), .ip2(n6755), .ip3(n6754), .ip4(n6753), .op(n6758) );
  nand2_1 U8108 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [18]), .op(n6757)
         );
  nand3_1 U8109 ( .ip1(n6759), .ip2(n6758), .ip3(n6757), .op(n6760) );
  not_ab_or_c_or_d U8110 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [18]), .ip2(n6766), 
        .ip3(n6761), .ip4(n6760), .op(n9391) );
  nand2_1 U8111 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [20]), .ip2(n6762), .op(n6778)
         );
  and2_1 U8112 ( .ip1(n6763), .ip2(\CORTEXM0DS_INST/cm0_r00 [20]), .op(n6773)
         );
  nand2_1 U8113 ( .ip1(n6764), .ip2(\CORTEXM0DS_INST/cm0_r05 [20]), .op(n6771)
         );
  nand2_1 U8114 ( .ip1(n6765), .ip2(\CORTEXM0DS_INST/cm0_r02 [20]), .op(n6770)
         );
  nand2_1 U8115 ( .ip1(n6766), .ip2(\CORTEXM0DS_INST/cm0_r04 [20]), .op(n6769)
         );
  nand2_1 U8116 ( .ip1(n6767), .ip2(\CORTEXM0DS_INST/cm0_r03 [20]), .op(n6768)
         );
  not_ab_or_c_or_d U8117 ( .ip1(n6774), .ip2(\CORTEXM0DS_INST/cm0_r01 [20]), 
        .ip3(n6773), .ip4(n6772), .op(n6777) );
  nand2_1 U8118 ( .ip1(n6775), .ip2(\CORTEXM0DS_INST/cm0_r06 [20]), .op(n6776)
         );
  nand3_1 U8119 ( .ip1(n6778), .ip2(n6777), .ip3(n6776), .op(n9367) );
  nor2_1 U8120 ( .ip1(n9367), .ip2(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .op(
        n6779) );
  not_ab_or_c_or_d U8121 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n9391), 
        .ip3(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip4(n6779), .op(n6780) );
  not_ab_or_c_or_d U8122 ( .ip1(n11120), .ip2(n9369), .ip3(n6781), .ip4(n6780), 
        .op(n6782) );
  mux2_1 U8123 ( .ip1(n6783), .ip2(n6782), .s(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .op(n6784) );
  nor2_1 U8124 ( .ip1(n6784), .ip2(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .op(
        n6785) );
  not_ab_or_c_or_d U8125 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(n6786), 
        .ip3(n6785), .ip4(n10891), .op(n6787) );
  not_ab_or_c_or_d U8126 ( .ip1(n6789), .ip2(n11008), .ip3(n6788), .ip4(n6787), 
        .op(n6796) );
  nand2_1 U8127 ( .ip1(n6796), .ip2(n8948), .op(n8992) );
  nand2_1 U8128 ( .ip1(n12625), .ip2(n6210), .op(n12072) );
  nand2_1 U8129 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n11654), .op(
        n6790) );
  nand4_1 U8130 ( .ip1(n6791), .ip2(n8992), .ip3(n12072), .ip4(n6790), .op(
        n6792) );
  not_ab_or_c_or_d U8131 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n6794), 
        .ip3(n6793), .ip4(n6792), .op(n6795) );
  nor2_1 U8132 ( .ip1(n12599), .ip2(n6795), .op(n12300) );
  inv_1 U8133 ( .ip(n12300), .op(n12309) );
  nor2_1 U8134 ( .ip1(n11018), .ip2(n12309), .op(n6802) );
  nor2_1 U8135 ( .ip1(n12096), .ip2(n11730), .op(n12034) );
  or2_1 U8136 ( .ip1(n12051), .ip2(n6796), .op(n9002) );
  nand2_1 U8137 ( .ip1(n10937), .ip2(n10899), .op(n9653) );
  inv_1 U8138 ( .ip(n10903), .op(n9753) );
  inv_1 U8139 ( .ip(n8819), .op(n7765) );
  nand2_1 U8140 ( .ip1(n7765), .ip2(n11212), .op(n10490) );
  nand3_1 U8141 ( .ip1(n9753), .ip2(n12603), .ip3(n10490), .op(n6797) );
  inv_1 U8142 ( .ip(n8623), .op(n10972) );
  nand3_1 U8143 ( .ip1(n10972), .ip2(n12096), .ip3(n11730), .op(n8457) );
  not_ab_or_c_or_d U8144 ( .ip1(n12034), .ip2(n12095), .ip3(n6799), .ip4(n6798), .op(n6800) );
  nor2_1 U8145 ( .ip1(n12599), .ip2(n6800), .op(n12314) );
  inv_1 U8146 ( .ip(n12314), .op(n12295) );
  nor2_1 U8147 ( .ip1(n9183), .ip2(n12295), .op(n6801) );
  or2_1 U8148 ( .ip1(n6802), .ip2(n6801), .op(n12286) );
  or2_1 U8149 ( .ip1(n8796), .ip2(n12286), .op(n6843) );
  and2_1 U8150 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [1]), .op(n6812)
         );
  nand2_1 U8151 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [1]), .op(n6806)
         );
  nand2_1 U8152 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [1]), .op(n6805)
         );
  nand2_1 U8153 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [1]), .op(n6804)
         );
  nand2_1 U8154 ( .ip1(n8966), .ip2(\CORTEXM0DS_INST/cm0_r12 [1]), .op(n6803)
         );
  and4_1 U8155 ( .ip1(n6806), .ip2(n6805), .ip3(n6804), .ip4(n6803), .op(n6810) );
  nand2_1 U8156 ( .ip1(n8946), .ip2(n9332), .op(n6809) );
  nand2_1 U8157 ( .ip1(\CORTEXM0DS_INST/u_logic/Kycvx4 ), .ip2(n8948), .op(
        n6808) );
  inv_1 U8158 ( .ip(n7975), .op(n8947) );
  nand2_1 U8159 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/Uzcvx4 ), .op(
        n6807) );
  ab_or_c_or_d U8160 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [1]), .ip2(n8957), .ip3(
        n6812), .ip4(n6811), .op(n9074) );
  nor2_1 U8161 ( .ip1(n12639), .ip2(n8537), .op(n6945) );
  not_ab_or_c_or_d U8162 ( .ip1(n12639), .ip2(n8537), .ip3(n6945), .ip4(n12305), .op(n6841) );
  nand4_1 U8163 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/O8gvx4 ), .ip4(n11206), .op(n8008) );
  inv_1 U8164 ( .ip(n8008), .op(n8295) );
  and2_1 U8165 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [1]), .op(n6828)
         );
  and2_1 U8166 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [1]), .op(n6822)
         );
  nand2_1 U8167 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [1]), .op(n6821)
         );
  and2_1 U8168 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [1]), .op(n6818)
         );
  nand2_1 U8169 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [1]), .op(n6816)
         );
  nand2_1 U8170 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [1]), .op(n6815)
         );
  nand2_1 U8171 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [1]), .op(n6814)
         );
  nand2_1 U8172 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [1]), .op(n6813)
         );
  not_ab_or_c_or_d U8173 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [1]), .ip2(n8903), 
        .ip3(n6818), .ip4(n6817), .op(n6820) );
  nand2_1 U8174 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [1]), .op(n6819)
         );
  nand3_1 U8175 ( .ip1(n6821), .ip2(n6820), .ip3(n6819), .op(n6967) );
  not_ab_or_c_or_d U8176 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [1]), .ip2(n8910), 
        .ip3(n6822), .ip4(n6967), .op(n6826) );
  nand2_1 U8177 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [1]), .op(n6825)
         );
  nand2_1 U8178 ( .ip1(n8853), .ip2(\CORTEXM0DS_INST/u_logic/Uzcvx4 ), .op(
        n6824) );
  nand2_1 U8179 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [1]), .op(n6823)
         );
  not_ab_or_c_or_d U8180 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [1]), .ip2(n8914), 
        .ip3(n6828), .ip4(n6827), .op(n8789) );
  nor2_1 U8181 ( .ip1(n8789), .ip2(n8292), .op(n6831) );
  nor2_1 U8182 ( .ip1(n6829), .ip2(n6965), .op(n6830) );
  not_ab_or_c_or_d U8183 ( .ip1(n8295), .ip2(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), 
        .ip3(n6831), .ip4(n6830), .op(n6832) );
  mux2_1 U8184 ( .ip1(n8013), .ip2(n8297), .s(n6832), .op(n9077) );
  and2_1 U8185 ( .ip1(n6833), .ip2(n9181), .op(n6834) );
  nand2_1 U8186 ( .ip1(n9074), .ip2(n6834), .op(n6899) );
  inv_1 U8187 ( .ip(n6899), .op(n6836) );
  or2_1 U8188 ( .ip1(n9074), .ip2(n6834), .op(n6835) );
  nand2_1 U8189 ( .ip1(n8969), .ip2(n6835), .op(n6898) );
  nor2_1 U8190 ( .ip1(n6836), .ip2(n6898), .op(n6837) );
  xor2_1 U8191 ( .ip1(n9077), .ip2(n6837), .op(n6942) );
  nand2_1 U8192 ( .ip1(n6839), .ip2(n6838), .op(n6941) );
  xnor2_1 U8193 ( .ip1(n6942), .ip2(n6941), .op(n10856) );
  nor2_1 U8194 ( .ip1(n10856), .ip2(n12309), .op(n6840) );
  ab_or_c_or_d U8195 ( .ip1(n12314), .ip2(n9074), .ip3(n6841), .ip4(n6840), 
        .op(n11153) );
  or2_1 U8196 ( .ip1(n11153), .ip2(n12286), .op(n6842) );
  nand2_1 U8197 ( .ip1(n6843), .ip2(n6842), .op(n6844) );
  or2_1 U8198 ( .ip1(n9801), .ip2(n6844), .op(n12600) );
  inv_1 U8199 ( .ip(n8292), .op(n8011) );
  inv_1 U8200 ( .ip(\CORTEXM0DS_INST/u_logic/O7evx4 ), .op(n11526) );
  nor2_1 U8201 ( .ip1(n6847), .ip2(n6846), .op(n6863) );
  and2_1 U8202 ( .ip1(n11526), .ip2(n6863), .op(n8922) );
  and2_1 U8203 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [3]), .op(n6849)
         );
  inv_1 U8204 ( .ip(n8910), .op(n8143) );
  inv_1 U8205 ( .ip(\CORTEXM0DS_INST/cm0_r14 [3]), .op(n6882) );
  nor2_1 U8206 ( .ip1(n8143), .ip2(n6882), .op(n6848) );
  not_ab_or_c_or_d U8207 ( .ip1(\CORTEXM0DS_INST/vis_msp [1]), .ip2(n8922), 
        .ip3(n6849), .ip4(n6848), .op(n6867) );
  nand2_1 U8208 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [3]), .op(n6858)
         );
  and2_1 U8209 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [3]), .op(n6855)
         );
  nand2_1 U8210 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [3]), .op(n6853)
         );
  nand2_1 U8211 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [3]), .op(n6852)
         );
  nand2_1 U8212 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [3]), .op(n6851)
         );
  nand2_1 U8213 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [3]), .op(n6850)
         );
  not_ab_or_c_or_d U8214 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [3]), .ip2(n8934), 
        .ip3(n6855), .ip4(n6854), .op(n6857) );
  nand2_1 U8215 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [3]), .op(n6856)
         );
  nand3_1 U8216 ( .ip1(n6858), .ip2(n6857), .ip3(n6856), .op(n7017) );
  nand2_1 U8217 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [3]), .op(n6861)
         );
  nand2_1 U8218 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [3]), .op(n6860)
         );
  nand2_1 U8219 ( .ip1(n8853), .ip2(\CORTEXM0DS_INST/u_logic/O2dvx4 ), .op(
        n6859) );
  nand3_1 U8220 ( .ip1(n6861), .ip2(n6860), .ip3(n6859), .op(n6862) );
  not_ab_or_c_or_d U8221 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [3]), 
        .ip3(n7017), .ip4(n6862), .op(n6866) );
  and2_1 U8222 ( .ip1(n6863), .ip2(\CORTEXM0DS_INST/u_logic/O7evx4 ), .op(
        n8923) );
  nand2_1 U8223 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [1]), .op(n6865)
         );
  nand2_1 U8224 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [3]), .op(n6864)
         );
  nand2_1 U8225 ( .ip1(n8011), .ip2(n12673), .op(n6880) );
  nand2_1 U8226 ( .ip1(\CORTEXM0DS_INST/u_logic/I29vx4 ), .ip2(n8295), .op(
        n6879) );
  nand2_1 U8227 ( .ip1(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .ip2(n7670), .op(
        n6878) );
  nor4_1 U8228 ( .ip1(n12625), .ip2(n8553), .ip3(n11183), .ip4(n12649), .op(
        n11755) );
  and3_1 U8229 ( .ip1(n9748), .ip2(n10880), .ip3(n11754), .op(n6871) );
  nor4_1 U8230 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip3(n10865), .ip4(n12613), .op(
        n6870) );
  nor2_1 U8231 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n12614), .op(
        n6868) );
  nor3_1 U8232 ( .ip1(n6868), .ip2(n10899), .ip3(n12616), .op(n6869) );
  or2_1 U8233 ( .ip1(n7536), .ip2(n9582), .op(n6876) );
  nand2_1 U8234 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10547), .op(
        n12618) );
  not_ab_or_c_or_d U8235 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n12618), .ip3(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip4(n12625), .op(n6873) );
  nor2_1 U8236 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n10547), .op(
        n10538) );
  nor2_1 U8237 ( .ip1(n9598), .ip2(n10538), .op(n11162) );
  nor4_1 U8238 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n10937), .ip3(
        n11162), .ip4(n10949), .op(n6872) );
  nor2_1 U8239 ( .ip1(n12096), .ip2(n12072), .op(n10938) );
  nor2_1 U8240 ( .ip1(n12613), .ip2(n12603), .op(n11195) );
  or2_1 U8241 ( .ip1(n6874), .ip2(n9582), .op(n6875) );
  nand2_1 U8242 ( .ip1(n6876), .ip2(n6875), .op(n7682) );
  nand2_1 U8243 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n7682), .op(
        n6877) );
  mux2_1 U8244 ( .ip1(n8297), .ip2(n8013), .s(n6881), .op(n9071) );
  inv_1 U8245 ( .ip(n9071), .op(n9066) );
  inv_1 U8246 ( .ip(n8958), .op(n8154) );
  nor2_1 U8247 ( .ip1(n8154), .ip2(n6882), .op(n6897) );
  and2_1 U8248 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [3]), .op(n6890)
         );
  nand2_1 U8249 ( .ip1(n8946), .ip2(n6976), .op(n6888) );
  nand2_1 U8250 ( .ip1(\CORTEXM0DS_INST/u_logic/E1dvx4 ), .ip2(n8948), .op(
        n6887) );
  nand2_1 U8251 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/O2dvx4 ), .op(
        n6886) );
  or2_1 U8252 ( .ip1(n6884), .ip2(n6883), .op(n6891) );
  nor2_1 U8253 ( .ip1(\CORTEXM0DS_INST/u_logic/O7evx4 ), .ip2(n6891), .op(
        n8949) );
  nand2_1 U8254 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [1]), .op(n6885)
         );
  not_ab_or_c_or_d U8255 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [3]), .ip2(n8966), 
        .ip3(n6890), .ip4(n6889), .op(n6895) );
  nand2_1 U8256 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [3]), .op(n6894)
         );
  nand2_1 U8257 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [3]), .op(n6893)
         );
  nor2_1 U8258 ( .ip1(n11526), .ip2(n6891), .op(n8959) );
  nand2_1 U8259 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [1]), .op(n6892)
         );
  nand4_1 U8260 ( .ip1(n6895), .ip2(n6894), .ip3(n6893), .ip4(n6892), .op(
        n6896) );
  not_ab_or_c_or_d U8261 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [3]), 
        .ip3(n6897), .ip4(n6896), .op(n9070) );
  nor2_1 U8262 ( .ip1(n8974), .ip2(n9070), .op(n7381) );
  or2_1 U8263 ( .ip1(n9077), .ip2(n6898), .op(n6900) );
  nand2_1 U8264 ( .ip1(n6900), .ip2(n6899), .op(n6944) );
  nor3_1 U8265 ( .ip1(n12096), .ip2(n12625), .ip3(n9582), .op(n6913) );
  inv_1 U8266 ( .ip(n8944), .op(n7367) );
  inv_1 U8267 ( .ip(\CORTEXM0DS_INST/cm0_r10 [2]), .op(n6915) );
  nor2_1 U8268 ( .ip1(n7367), .ip2(n6915), .op(n6912) );
  and2_1 U8269 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [2]), .op(n6906)
         );
  nand2_1 U8270 ( .ip1(n8946), .ip2(n7100), .op(n6904) );
  nand2_1 U8271 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/E1dvx4 ), .op(
        n6903) );
  nand2_1 U8272 ( .ip1(\CORTEXM0DS_INST/u_logic/Uzcvx4 ), .ip2(n8948), .op(
        n6902) );
  nand2_1 U8273 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [0]), .op(n6901)
         );
  not_ab_or_c_or_d U8274 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [2]), .ip2(n8958), 
        .ip3(n6906), .ip4(n6905), .op(n6910) );
  nand2_1 U8275 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [2]), .op(n6909)
         );
  nand2_1 U8276 ( .ip1(n8966), .ip2(\CORTEXM0DS_INST/cm0_r12 [2]), .op(n6908)
         );
  nand2_1 U8277 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [0]), .op(n6907)
         );
  nand4_1 U8278 ( .ip1(n6910), .ip2(n6909), .ip3(n6908), .ip4(n6907), .op(
        n6911) );
  not_ab_or_c_or_d U8279 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [2]), .ip2(n8956), 
        .ip3(n6912), .ip4(n6911), .op(n9180) );
  not_ab_or_c_or_d U8280 ( .ip1(n6913), .ip2(n11746), .ip3(n8974), .ip4(n9180), 
        .op(n6943) );
  nand2_1 U8281 ( .ip1(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip2(n7682), .op(
        n6938) );
  nand2_1 U8282 ( .ip1(\CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip2(n6914), .op(
        n6937) );
  nand2_1 U8283 ( .ip1(n8295), .ip2(\CORTEXM0DS_INST/u_logic/B19vx4 ), .op(
        n6936) );
  inv_1 U8284 ( .ip(n8916), .op(n7349) );
  nor2_1 U8285 ( .ip1(n7349), .ip2(n6915), .op(n6917) );
  and2_1 U8286 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [0]), .op(n6916)
         );
  not_ab_or_c_or_d U8287 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [2]), .ip2(n8914), 
        .ip3(n6917), .ip4(n6916), .op(n6934) );
  nand2_1 U8288 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [2]), .op(n6926)
         );
  and2_1 U8289 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [2]), .op(n6923)
         );
  nand2_1 U8290 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [2]), .op(n6921)
         );
  nand2_1 U8291 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [2]), .op(n6920)
         );
  nand2_1 U8292 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [2]), .op(n6919)
         );
  nand2_1 U8293 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [2]), .op(n6918)
         );
  not_ab_or_c_or_d U8294 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [2]), .ip2(n8925), 
        .ip3(n6923), .ip4(n6922), .op(n6925) );
  nand2_1 U8295 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [2]), .op(n6924)
         );
  nand3_1 U8296 ( .ip1(n6926), .ip2(n6925), .ip3(n6924), .op(n6962) );
  nand2_1 U8297 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [2]), .ip2(n8910), .op(n6929)
         );
  nand2_1 U8298 ( .ip1(n8853), .ip2(\CORTEXM0DS_INST/u_logic/E1dvx4 ), .op(
        n6928) );
  nand2_1 U8299 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [2]), .op(n6927)
         );
  nand3_1 U8300 ( .ip1(n6929), .ip2(n6928), .ip3(n6927), .op(n6930) );
  not_ab_or_c_or_d U8301 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [2]), 
        .ip3(n6962), .ip4(n6930), .op(n6933) );
  nand2_1 U8302 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [0]), .op(n6932)
         );
  nand2_1 U8303 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [2]), .op(n6931)
         );
  nand2_1 U8304 ( .ip1(n8011), .ip2(n12667), .op(n6935) );
  mux2_1 U8305 ( .ip1(n8013), .ip2(n8297), .s(n6939), .op(n9175) );
  inv_1 U8306 ( .ip(n6940), .op(n7383) );
  nor2_1 U8307 ( .ip1(n6942), .ip2(n6941), .op(n7338) );
  fulladder U8308 ( .a(n6944), .b(n6943), .ci(n9175), .co(n7380), .s(n7337) );
  nand2_1 U8309 ( .ip1(n7338), .ip2(n7337), .op(n7382) );
  xor2_1 U8310 ( .ip1(n7383), .ip2(n7382), .op(n11390) );
  nand2_1 U8311 ( .ip1(\CORTEXM0DS_INST/u_logic/I4gvx4 ), .ip2(n6945), .op(
        n6947) );
  inv_1 U8312 ( .ip(\CORTEXM0DS_INST/u_logic/I4gvx4 ), .op(n8500) );
  mux2_1 U8313 ( .ip1(n6946), .ip2(n8500), .s(n6945), .op(n7339) );
  nand2_1 U8314 ( .ip1(n7339), .ip2(\CORTEXM0DS_INST/vis_pc [1]), .op(n7340)
         );
  and2_1 U8315 ( .ip1(n6947), .ip2(n7340), .op(n6948) );
  inv_1 U8316 ( .ip(\CORTEXM0DS_INST/vis_pc [2]), .op(n7392) );
  nor2_1 U8317 ( .ip1(n7392), .ip2(n6948), .op(n7384) );
  not_ab_or_c_or_d U8318 ( .ip1(n6948), .ip2(n7392), .ip3(n7384), .ip4(n12305), 
        .op(n6950) );
  nor2_1 U8319 ( .ip1(n9070), .ip2(n12295), .op(n6949) );
  not_ab_or_c_or_d U8320 ( .ip1(n12300), .ip2(n11390), .ip3(n6950), .ip4(n6949), .op(\CORTEXM0DS_INST/u_logic/Ekovx4 ) );
  nand2_1 U8321 ( .ip1(\CORTEXM0DS_INST/u_logic/Uzcvx4 ), .ip2(n2120), .op(
        n6955) );
  nor2_1 U8322 ( .ip1(n2120), .ip2(n11729), .op(n12321) );
  nand2_1 U8323 ( .ip1(\CORTEXM0DS_INST/vis_pc [0]), .ip2(n12321), .op(n6954)
         );
  nand2_1 U8324 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n11184), .op(
        n11222) );
  nor2_1 U8325 ( .ip1(n2120), .ip2(n11222), .op(n12320) );
  nand2_1 U8326 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [1]), .ip2(n12320), .op(n6953) );
  nand2_1 U8327 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n10547), .op(
        n8451) );
  inv_1 U8328 ( .ip(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .op(n12588) );
  nor2_1 U8329 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Ud9vx4 ), .op(n9463) );
  nor2_1 U8330 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n11038), .op(
        n6989) );
  and3_1 U8331 ( .ip1(n9463), .ip2(n6989), .ip3(n12329), .op(n6951) );
  not_ab_or_c_or_d U8332 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n8451), 
        .ip3(n2120), .ip4(n6951), .op(n12691) );
  nand2_1 U8333 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n12075), .op(
        n10701) );
  inv_1 U8334 ( .ip(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .op(n12592) );
  nand2_1 U8335 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n12592), .op(
        n10506) );
  inv_1 U8336 ( .ip(n10506), .op(n10454) );
  nand2_1 U8337 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n10454), .op(
        n11053) );
  nand4_1 U8338 ( .ip1(n12691), .ip2(n10701), .ip3(n11153), .ip4(n11053), .op(
        n6952) );
  nand4_1 U8339 ( .ip1(n6955), .ip2(n6954), .ip3(n6953), .ip4(n6952), .op(
        n6083) );
  nor2_1 U8340 ( .ip1(n9781), .ip2(n11846), .op(n12395) );
  and3_1 U8341 ( .ip1(n6957), .ip2(n6956), .ip3(
        \CORTEXM0DS_INST/u_logic/Ul8vx4 ), .op(n6959) );
  inv_1 U8342 ( .ip(n6958), .op(LOCKUP_top_out) );
  not_ab_or_c_or_d U8343 ( .ip1(\CORTEXM0DS_INST/u_logic/Mk8vx4 ), .ip2(n12395), .ip3(n6959), .ip4(LOCKUP_top_out), .op(n6960) );
  nor2_1 U8344 ( .ip1(n5822), .ip2(n6960), .op(n10858) );
  inv_1 U8345 ( .ip(n10858), .op(n10573) );
  nand2_1 U8346 ( .ip1(n9634), .ip2(n8823), .op(n11017) );
  nor2_1 U8347 ( .ip1(n5822), .ip2(n11017), .op(n10572) );
  nand2_1 U8348 ( .ip1(n11390), .ip2(n10572), .op(n7336) );
  nor2_1 U8349 ( .ip1(n11016), .ip2(n5822), .op(n10859) );
  nor2_1 U8350 ( .ip1(n10859), .ip2(n10572), .op(n12091) );
  inv_1 U8351 ( .ip(\CORTEXM0DS_INST/vis_pc [1]), .op(n12394) );
  nor3_1 U8352 ( .ip1(n5822), .ip2(n12394), .ip3(n8537), .op(n10380) );
  or2_1 U8353 ( .ip1(\CORTEXM0DS_INST/vis_pc [2]), .ip2(n10380), .op(n6961) );
  nand2_1 U8354 ( .ip1(\CORTEXM0DS_INST/vis_pc [2]), .ip2(n10380), .op(n10375)
         );
  nand3_1 U8355 ( .ip1(n12091), .ip2(n6961), .ip3(n10375), .op(n7335) );
  inv_1 U8356 ( .ip(n12618), .op(n10969) );
  nand2_1 U8357 ( .ip1(\CORTEXM0DS_INST/u_logic/Dw8vx4 ), .ip2(n10969), .op(
        n7015) );
  inv_1 U8358 ( .ip(n7015), .op(n7054) );
  nand2_1 U8359 ( .ip1(\CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip2(n7054), .op(
        n6964) );
  nand2_1 U8360 ( .ip1(\CORTEXM0DS_INST/u_logic/Dw8vx4 ), .ip2(n11715), .op(
        n7052) );
  inv_1 U8361 ( .ip(n7052), .op(n9503) );
  nand2_1 U8362 ( .ip1(n9503), .ip2(n6962), .op(n6963) );
  nand2_1 U8363 ( .ip1(n6964), .ip2(n6963), .op(n7020) );
  nor2_1 U8364 ( .ip1(n6965), .ip2(n7015), .op(n6966) );
  or2_1 U8365 ( .ip1(n9503), .ip2(n6966), .op(n6969) );
  or2_1 U8366 ( .ip1(n6967), .ip2(n6966), .op(n6968) );
  nand2_1 U8367 ( .ip1(n6969), .ip2(n6968), .op(n6978) );
  nor2_1 U8368 ( .ip1(n11145), .ip2(n7015), .op(n6970) );
  or2_1 U8369 ( .ip1(n9503), .ip2(n6970), .op(n6973) );
  or2_1 U8370 ( .ip1(n6971), .ip2(n6970), .op(n6972) );
  nand2_1 U8371 ( .ip1(n6973), .ip2(n6972), .op(n6980) );
  nand2_1 U8372 ( .ip1(n6978), .ip2(n6980), .op(n9420) );
  nand2_1 U8373 ( .ip1(n9420), .ip2(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .op(
        n6974) );
  xor2_1 U8374 ( .ip1(n7020), .ip2(n6974), .op(n9338) );
  nand2_1 U8375 ( .ip1(n11730), .ip2(n12625), .op(n10599) );
  nand2_1 U8376 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n10599), .op(
        n7000) );
  nand3_1 U8377 ( .ip1(n11214), .ip2(n7000), .ip3(n7094), .op(n6975) );
  nand2_1 U8378 ( .ip1(\CORTEXM0DS_INST/u_logic/Dw8vx4 ), .ip2(n6975), .op(
        n11811) );
  inv_1 U8379 ( .ip(n11811), .op(n11821) );
  nand2_1 U8380 ( .ip1(n9338), .ip2(n11821), .op(n10148) );
  inv_1 U8381 ( .ip(n10148), .op(n11607) );
  inv_1 U8382 ( .ip(n6976), .op(n9296) );
  nor2_1 U8383 ( .ip1(n9296), .ip2(n9420), .op(n6984) );
  inv_1 U8384 ( .ip(n9263), .op(n9258) );
  inv_1 U8385 ( .ip(n6980), .op(n6979) );
  nor2_1 U8386 ( .ip1(n6979), .ip2(n6978), .op(n9433) );
  inv_1 U8387 ( .ip(n9433), .op(n9418) );
  nor2_1 U8388 ( .ip1(n9258), .ip2(n9418), .op(n6983) );
  inv_1 U8389 ( .ip(n9264), .op(n9257) );
  nor2_1 U8390 ( .ip1(n6980), .ip2(n11754), .op(n6977) );
  xor2_1 U8391 ( .ip1(n6978), .ip2(n6977), .op(n9345) );
  nand2_1 U8392 ( .ip1(n9345), .ip2(n6979), .op(n9416) );
  nor2_1 U8393 ( .ip1(n9257), .ip2(n9416), .op(n6982) );
  nor2_1 U8394 ( .ip1(n6980), .ip2(n9345), .op(n9435) );
  and2_1 U8395 ( .ip1(n9282), .ip2(n9435), .op(n6981) );
  nor4_1 U8396 ( .ip1(n6984), .ip2(n6983), .ip3(n6982), .ip4(n6981), .op(n9339) );
  inv_1 U8397 ( .ip(n9339), .op(n6998) );
  inv_1 U8398 ( .ip(n9416), .op(n9429) );
  and2_1 U8399 ( .ip1(n9283), .ip2(n9429), .op(n6988) );
  inv_1 U8400 ( .ip(n9281), .op(n7628) );
  nor2_1 U8401 ( .ip1(n7628), .ip2(n9420), .op(n6987) );
  and2_1 U8402 ( .ip1(n9284), .ip2(n9433), .op(n6986) );
  and2_1 U8403 ( .ip1(n9275), .ip2(n9435), .op(n6985) );
  nor4_1 U8404 ( .ip1(n6988), .ip2(n6987), .ip3(n6986), .ip4(n6985), .op(n9292) );
  inv_1 U8405 ( .ip(n9338), .op(n9443) );
  nand2_1 U8406 ( .ip1(n11821), .ip2(n9443), .op(n11614) );
  nor2_1 U8407 ( .ip1(n9292), .ip2(n11614), .op(n6997) );
  nor2_1 U8408 ( .ip1(n11736), .ip2(n6989), .op(n12389) );
  nor4_1 U8409 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip3(n12095), .ip4(n10547), .op(
        n7062) );
  nor3_1 U8410 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n12615), .ip3(
        n10949), .op(n8622) );
  not_ab_or_c_or_d U8411 ( .ip1(n12389), .ip2(n11191), .ip3(n7062), .ip4(n8622), .op(n6990) );
  inv_1 U8412 ( .ip(\CORTEXM0DS_INST/u_logic/Dw8vx4 ), .op(n9514) );
  nor2_1 U8413 ( .ip1(n6990), .ip2(n9514), .op(n11807) );
  inv_1 U8414 ( .ip(n11807), .op(n11839) );
  inv_1 U8415 ( .ip(\CORTEXM0DS_INST/u_logic/N6hvx4 ), .op(n7305) );
  nor4_1 U8416 ( .ip1(\CORTEXM0DS_INST/u_logic/Z7hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/L9hvx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/B5hvx4 ), .ip4(n7305), .op(n11800) );
  inv_1 U8417 ( .ip(n11800), .op(n8803) );
  nor2_1 U8418 ( .ip1(n11839), .ip2(n8803), .op(n11787) );
  inv_1 U8419 ( .ip(\CORTEXM0DS_INST/u_logic/Xahvx4 ), .op(n11865) );
  nor2_1 U8420 ( .ip1(\CORTEXM0DS_INST/u_logic/N6hvx4 ), .ip2(n11865), .op(
        n10171) );
  inv_1 U8421 ( .ip(n10171), .op(n6991) );
  inv_1 U8422 ( .ip(\CORTEXM0DS_INST/u_logic/Z7hvx4 ), .op(n10209) );
  nor3_1 U8423 ( .ip1(\CORTEXM0DS_INST/u_logic/L9hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/B5hvx4 ), .ip3(n10209), .op(n12682) );
  nand2_1 U8424 ( .ip1(n11807), .ip2(n12682), .op(n9976) );
  nor2_1 U8425 ( .ip1(n6991), .ip2(n9976), .op(n9977) );
  nor2_1 U8426 ( .ip1(\CORTEXM0DS_INST/u_logic/N6hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Xahvx4 ), .op(n12683) );
  inv_1 U8427 ( .ip(n12683), .op(n12685) );
  inv_1 U8428 ( .ip(\CORTEXM0DS_INST/u_logic/L9hvx4 ), .op(n10208) );
  inv_1 U8429 ( .ip(\CORTEXM0DS_INST/u_logic/B5hvx4 ), .op(n10168) );
  nor4_1 U8430 ( .ip1(n12685), .ip2(n10208), .ip3(n10209), .ip4(n10168), .op(
        n11866) );
  nand2_1 U8431 ( .ip1(n11866), .ip2(n11807), .op(n11810) );
  inv_1 U8432 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [3]), .op(n11894) );
  nor2_1 U8433 ( .ip1(n11810), .ip2(n11894), .op(n6992) );
  not_ab_or_c_or_d U8434 ( .ip1(n11787), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [3]), .ip3(n9977), .ip4(n6992), .op(
        n6995) );
  nand2_1 U8435 ( .ip1(\CORTEXM0DS_INST/u_logic/B5hvx4 ), .ip2(n10209), .op(
        n7304) );
  nor3_1 U8436 ( .ip1(\CORTEXM0DS_INST/u_logic/L9hvx4 ), .ip2(n7305), .ip3(
        n7304), .op(n11801) );
  nand2_1 U8437 ( .ip1(n11807), .ip2(n11801), .op(n11841) );
  inv_1 U8438 ( .ip(n11841), .op(n10265) );
  nand2_1 U8439 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [3]), .ip2(n10265), 
        .op(n6994) );
  nor2_1 U8440 ( .ip1(\CORTEXM0DS_INST/u_logic/L9hvx4 ), .ip2(n7304), .op(
        n11867) );
  nand2_1 U8441 ( .ip1(n11867), .ip2(n10171), .op(n8536) );
  nor2_1 U8442 ( .ip1(n11839), .ip2(n8536), .op(n11610) );
  nand2_1 U8443 ( .ip1(n11610), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [3]), 
        .op(n6993) );
  nand4_1 U8444 ( .ip1(n4203), .ip2(n6995), .ip3(n6994), .ip4(n6993), .op(
        n6996) );
  not_ab_or_c_or_d U8445 ( .ip1(n11607), .ip2(n6998), .ip3(n6997), .ip4(n6996), 
        .op(n10398) );
  nor2_1 U8446 ( .ip1(\CORTEXM0DS_INST/u_logic/Zph2z4 [1]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zph2z4 [0]), .op(n7118) );
  not_ab_or_c_or_d U8447 ( .ip1(n7118), .ip2(n7000), .ip3(n6999), .ip4(n12095), 
        .op(n7002) );
  nor2_1 U8448 ( .ip1(n12338), .ip2(n10770), .op(n8609) );
  nor3_1 U8449 ( .ip1(n7001), .ip2(n10779), .ip3(n8609), .op(n10043) );
  inv_1 U8450 ( .ip(n10043), .op(n9933) );
  nor2_1 U8451 ( .ip1(n7002), .ip2(n9933), .op(n7061) );
  nor3_1 U8452 ( .ip1(n11181), .ip2(n10865), .ip3(n11038), .op(n7003) );
  nor2_1 U8453 ( .ip1(n7003), .ip2(n9933), .op(n10050) );
  nand2_1 U8454 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(n7054), .op(
        n7014) );
  nand2_1 U8455 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [4]), .op(n7012)
         );
  and2_1 U8456 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [4]), .op(n7009)
         );
  nand2_1 U8457 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [4]), .op(n7007)
         );
  nand2_1 U8458 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [4]), .op(n7006)
         );
  nand2_1 U8459 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [4]), .op(n7005)
         );
  nand2_1 U8460 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [4]), .op(n7004)
         );
  not_ab_or_c_or_d U8461 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [4]), .ip2(n8925), 
        .ip3(n7009), .ip4(n7008), .op(n7011) );
  nand2_1 U8462 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [4]), .op(n7010)
         );
  nand3_1 U8463 ( .ip1(n7012), .ip2(n7011), .ip3(n7010), .op(n7356) );
  nand2_1 U8464 ( .ip1(n9503), .ip2(n7356), .op(n7013) );
  nand2_1 U8465 ( .ip1(n7014), .ip2(n7013), .op(n7800) );
  inv_1 U8466 ( .ip(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .op(n11079) );
  nor2_1 U8467 ( .ip1(n11079), .ip2(n7015), .op(n7016) );
  or2_1 U8468 ( .ip1(n9503), .ip2(n7016), .op(n7019) );
  or2_1 U8469 ( .ip1(n7017), .ip2(n7016), .op(n7018) );
  nand2_1 U8470 ( .ip1(n7019), .ip2(n7018), .op(n7024) );
  nor2_1 U8471 ( .ip1(n9420), .ip2(n7020), .op(n7022) );
  nand2_1 U8472 ( .ip1(n7024), .ip2(n7022), .op(n7021) );
  nor2_1 U8473 ( .ip1(n7800), .ip2(n7021), .op(n9464) );
  nor2_1 U8474 ( .ip1(n9464), .ip2(n11754), .op(n9256) );
  and2_1 U8475 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n7021), .op(
        n7328) );
  xor2_1 U8476 ( .ip1(n7800), .ip2(n7328), .op(n9465) );
  or2_1 U8477 ( .ip1(n11754), .ip2(n7022), .op(n7023) );
  xor2_1 U8478 ( .ip1(n7024), .ip2(n7023), .op(n7091) );
  nor2_1 U8479 ( .ip1(n9465), .ip2(n7091), .op(n9476) );
  inv_1 U8480 ( .ip(n9476), .op(n10048) );
  nand2_1 U8481 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [5]), .op(n7033)
         );
  and2_1 U8482 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [5]), .op(n7030)
         );
  nand2_1 U8483 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [5]), .op(n7028)
         );
  nand2_1 U8484 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [5]), .op(n7027)
         );
  nand2_1 U8485 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [5]), .op(n7026)
         );
  nand2_1 U8486 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [5]), .op(n7025)
         );
  not_ab_or_c_or_d U8487 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [5]), .ip2(n8925), 
        .ip3(n7030), .ip4(n7029), .op(n7032) );
  nand2_1 U8488 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [5]), .op(n7031)
         );
  nand3_1 U8489 ( .ip1(n7033), .ip2(n7032), .ip3(n7031), .op(n7677) );
  nand2_1 U8490 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [7]), .op(n7042)
         );
  and2_1 U8491 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [7]), .op(n7039)
         );
  nand2_1 U8492 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [7]), .op(n7037)
         );
  nand2_1 U8493 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [7]), .op(n7036)
         );
  nand2_1 U8494 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [7]), .op(n7035)
         );
  nand2_1 U8495 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [7]), .op(n7034)
         );
  not_ab_or_c_or_d U8496 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [7]), .ip2(n8917), 
        .ip3(n7039), .ip4(n7038), .op(n7041) );
  nand2_1 U8497 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [7]), .op(n7040)
         );
  nand3_1 U8498 ( .ip1(n7042), .ip2(n7041), .ip3(n7040), .op(n9499) );
  nand2_1 U8499 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [6]), .op(n7051)
         );
  and2_1 U8500 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [6]), .op(n7048)
         );
  nand2_1 U8501 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [6]), .op(n7046)
         );
  nand2_1 U8502 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [6]), .op(n7045)
         );
  nand2_1 U8503 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [6]), .op(n7044)
         );
  nand2_1 U8504 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [6]), .op(n7043)
         );
  not_ab_or_c_or_d U8505 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [6]), .ip2(n8903), 
        .ip3(n7048), .ip4(n7047), .op(n7050) );
  nand2_1 U8506 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [6]), .op(n7049)
         );
  nand3_1 U8507 ( .ip1(n7051), .ip2(n7050), .ip3(n7049), .op(n9498) );
  nor3_1 U8508 ( .ip1(n7677), .ip2(n9499), .ip3(n9498), .op(n7053) );
  nor2_1 U8509 ( .ip1(n7053), .ip2(n7052), .op(n7056) );
  or2_1 U8510 ( .ip1(n11008), .ip2(n7056), .op(n7059) );
  and4_1 U8511 ( .ip1(n11754), .ip2(n11079), .ip3(n7055), .ip4(n7054), .op(
        n7057) );
  or2_1 U8512 ( .ip1(n7057), .ip2(n7056), .op(n7058) );
  nand2_1 U8513 ( .ip1(n7059), .ip2(n7058), .op(n9505) );
  nor2_1 U8514 ( .ip1(n9505), .ip2(n11730), .op(n9361) );
  or2_1 U8515 ( .ip1(n9361), .ip2(n10043), .op(n10047) );
  nor3_1 U8516 ( .ip1(n9256), .ip2(n10048), .ip3(n10047), .op(n9872) );
  nor2_1 U8517 ( .ip1(n10050), .ip2(n9872), .op(n10395) );
  nand3_1 U8518 ( .ip1(n9869), .ip2(n10043), .ip3(
        \CORTEXM0DS_INST/u_logic/Mcgvx4 ), .op(n7060) );
  nand2_1 U8519 ( .ip1(n10395), .ip2(n7060), .op(n7725) );
  nor2_1 U8520 ( .ip1(n7061), .ip2(n7725), .op(n10382) );
  or2_1 U8521 ( .ip1(n10398), .ip2(n10382), .op(n7333) );
  inv_1 U8522 ( .ip(n7091), .op(n9466) );
  nand2_1 U8523 ( .ip1(n9466), .ip2(n9465), .op(n9479) );
  nor2_1 U8524 ( .ip1(n9361), .ip2(n9479), .op(n7801) );
  nand2_1 U8525 ( .ip1(n7801), .ip2(n9933), .op(n9873) );
  nor2_1 U8526 ( .ip1(n9256), .ip2(n9873), .op(n7331) );
  inv_1 U8527 ( .ip(n7062), .op(n7766) );
  or3_1 U8528 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Zph2z4 [0]), .op(n7063) );
  inv_1 U8529 ( .ip(\CORTEXM0DS_INST/u_logic/Zph2z4 [1]), .op(n7127) );
  not_ab_or_c_or_d U8530 ( .ip1(n7766), .ip2(n7063), .ip3(n7127), .ip4(n9933), 
        .op(n7064) );
  nor2_1 U8531 ( .ip1(n7331), .ip2(n7064), .op(n10846) );
  inv_1 U8532 ( .ip(n10846), .op(n11003) );
  nor2_1 U8533 ( .ip1(n7774), .ip2(n9418), .op(n7068) );
  inv_1 U8534 ( .ip(n9369), .op(n9393) );
  nor2_1 U8535 ( .ip1(n9393), .ip2(n9420), .op(n7067) );
  inv_1 U8536 ( .ip(n9367), .op(n8083) );
  nor2_1 U8537 ( .ip1(n8083), .ip2(n9416), .op(n7066) );
  inv_1 U8538 ( .ip(n9435), .op(n9392) );
  nor2_1 U8539 ( .ip1(n8014), .ip2(n9392), .op(n7065) );
  nor4_1 U8540 ( .ip1(n7068), .ip2(n7067), .ip3(n7066), .ip4(n7065), .op(n7315) );
  nor2_1 U8541 ( .ip1(n7315), .ip2(n10148), .op(n7071) );
  inv_1 U8542 ( .ip(n11810), .op(n11609) );
  nand2_1 U8543 ( .ip1(n11609), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [19]), 
        .op(n7069) );
  nand2_1 U8544 ( .ip1(n4185), .ip2(n7069), .op(n7070) );
  not_ab_or_c_or_d U8545 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [19]), .ip2(
        n11610), .ip3(n7071), .ip4(n7070), .op(n10394) );
  inv_1 U8546 ( .ip(n10394), .op(n10079) );
  nor3_1 U8547 ( .ip1(n9466), .ip2(n9465), .ip3(n10047), .op(n10053) );
  inv_1 U8548 ( .ip(n9256), .op(n9386) );
  nand3_1 U8549 ( .ip1(n10547), .ip2(n12096), .ip3(
        \CORTEXM0DS_INST/u_logic/Zph2z4 [0]), .op(n7090) );
  nor3_1 U8550 ( .ip1(\CORTEXM0DS_INST/u_logic/Zph2z4 [1]), .ip2(n9933), .ip3(
        n7090), .op(n7076) );
  nand2_1 U8551 ( .ip1(n10538), .ip2(n6210), .op(n7072) );
  or2_1 U8552 ( .ip1(n7072), .ip2(n9933), .op(n7075) );
  nand2_1 U8553 ( .ip1(n11202), .ip2(n10937), .op(n7073) );
  or2_1 U8554 ( .ip1(n7073), .ip2(n9933), .op(n7074) );
  nand2_1 U8555 ( .ip1(n7075), .ip2(n7074), .op(n7796) );
  not_ab_or_c_or_d U8556 ( .ip1(n10053), .ip2(n9386), .ip3(n7076), .ip4(n7796), 
        .op(n10996) );
  nand2_1 U8557 ( .ip1(n9429), .ip2(n9432), .op(n7080) );
  inv_1 U8558 ( .ip(n9420), .op(n9431) );
  nand2_1 U8559 ( .ip1(n9431), .ip2(n9428), .op(n7079) );
  inv_1 U8560 ( .ip(n9389), .op(n9434) );
  nand2_1 U8561 ( .ip1(n9433), .ip2(n9434), .op(n7078) );
  inv_1 U8562 ( .ip(n9391), .op(n9368) );
  nand2_1 U8563 ( .ip1(n9435), .ip2(n9368), .op(n7077) );
  nand4_1 U8564 ( .ip1(n7080), .ip2(n7079), .ip3(n7078), .ip4(n7077), .op(
        n7316) );
  nor2_1 U8565 ( .ip1(n9338), .ip2(n7316), .op(n9414) );
  nor2_1 U8566 ( .ip1(n9417), .ip2(n9418), .op(n7084) );
  and2_1 U8567 ( .ip1(n9276), .ip2(n9431), .op(n7083) );
  inv_1 U8568 ( .ip(n9269), .op(n9421) );
  nor2_1 U8569 ( .ip1(n9421), .ip2(n9416), .op(n7082) );
  nor2_1 U8570 ( .ip1(n9419), .ip2(n9392), .op(n7081) );
  nor4_1 U8571 ( .ip1(n7084), .ip2(n7083), .ip3(n7082), .ip4(n7081), .op(n9291) );
  and2_1 U8572 ( .ip1(n9338), .ip2(n9291), .op(n9426) );
  nor3_1 U8573 ( .ip1(n9414), .ip2(n9426), .ip3(n11811), .op(n7089) );
  nand2_1 U8574 ( .ip1(n11609), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [11]), 
        .op(n7087) );
  nand2_1 U8575 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [11]), .ip2(n11787), 
        .op(n7086) );
  nand2_1 U8576 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [11]), .ip2(n10265), 
        .op(n7085) );
  nand4_1 U8577 ( .ip1(n4190), .ip2(n7087), .ip3(n7086), .ip4(n7085), .op(
        n7088) );
  not_ab_or_c_or_d U8578 ( .ip1(n11610), .ip2(
        \CORTEXM0DS_INST/u_logic/Czh2z4 [11]), .ip3(n7089), .ip4(n7088), .op(
        n10396) );
  nor2_1 U8579 ( .ip1(n10996), .ip2(n10396), .op(n7114) );
  nor2_1 U8580 ( .ip1(n9933), .ip2(n7127), .op(n7767) );
  inv_1 U8581 ( .ip(n7090), .op(n7093) );
  nand2_1 U8582 ( .ip1(n7091), .ip2(n9465), .op(n9469) );
  nor2_1 U8583 ( .ip1(n9469), .ip2(n10047), .op(n7092) );
  nor3_1 U8584 ( .ip1(n11730), .ip2(n12625), .ip3(n9933), .op(n10054) );
  not_ab_or_c_or_d U8585 ( .ip1(n7767), .ip2(n7093), .ip3(n7092), .ip4(n10054), 
        .op(n10994) );
  nor3_1 U8586 ( .ip1(\CORTEXM0DS_INST/u_logic/Z7hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/B5hvx4 ), .ip3(n10208), .op(n10166) );
  nand3_1 U8587 ( .ip1(\CORTEXM0DS_INST/u_logic/N6hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Xahvx4 ), .ip3(n10166), .op(n12017) );
  or2_1 U8588 ( .ip1(n11839), .ip2(n12017), .op(n10267) );
  nand2_1 U8589 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n9753), .op(
        n7095) );
  nand2_1 U8590 ( .ip1(n7095), .ip2(n7094), .op(n7096) );
  nand2_1 U8591 ( .ip1(n7096), .ip2(n9329), .op(n7115) );
  nor2_1 U8592 ( .ip1(n7115), .ip2(n11811), .op(n10109) );
  inv_1 U8593 ( .ip(n9464), .op(n9500) );
  nand2_1 U8594 ( .ip1(n11754), .ip2(n11751), .op(n10055) );
  nand2_1 U8595 ( .ip1(n9500), .ip2(n10055), .op(n9325) );
  nor2_1 U8596 ( .ip1(n11730), .ip2(n9325), .op(n9357) );
  nor2_1 U8597 ( .ip1(n9338), .ip2(n9325), .op(n7099) );
  nand2_1 U8598 ( .ip1(n9338), .ip2(n9325), .op(n7097) );
  nand2_1 U8599 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n7097), .op(
        n7098) );
  nor2_1 U8600 ( .ip1(n7099), .ip2(n7098), .op(n9312) );
  mux2_1 U8601 ( .ip1(n9357), .ip2(n9312), .s(n9420), .op(n7110) );
  nand2_1 U8602 ( .ip1(n10109), .ip2(n7110), .op(n7112) );
  nor2_1 U8603 ( .ip1(n9294), .ip2(n9416), .op(n7104) );
  inv_1 U8604 ( .ip(n9332), .op(n9295) );
  nor2_1 U8605 ( .ip1(n9295), .ip2(n9418), .op(n7103) );
  nor2_1 U8606 ( .ip1(n8832), .ip2(n9420), .op(n7102) );
  inv_1 U8607 ( .ip(n7100), .op(n9293) );
  nor2_1 U8608 ( .ip1(n9293), .ip2(n9392), .op(n7101) );
  nor4_1 U8609 ( .ip1(n7104), .ip2(n7103), .ip3(n7102), .ip4(n7101), .op(n9340) );
  nand2_1 U8610 ( .ip1(n9429), .ip2(n9303), .op(n7108) );
  nand2_1 U8611 ( .ip1(n9431), .ip2(n9351), .op(n7107) );
  nand2_1 U8612 ( .ip1(n9433), .ip2(n9304), .op(n7106) );
  inv_1 U8613 ( .ip(n8888), .op(n9330) );
  nand2_1 U8614 ( .ip1(n9435), .ip2(n9330), .op(n7105) );
  nand4_1 U8615 ( .ip1(n7108), .ip2(n7107), .ip3(n7106), .ip4(n7105), .op(
        n9399) );
  nor2_1 U8616 ( .ip1(n9399), .ip2(n9443), .op(n7109) );
  not_ab_or_c_or_d U8617 ( .ip1(n9340), .ip2(n9443), .ip3(n7110), .ip4(n7109), 
        .op(n9314) );
  nand2_1 U8618 ( .ip1(n9314), .ip2(n11821), .op(n7111) );
  and4_1 U8619 ( .ip1(n4175), .ip2(n10267), .ip3(n7112), .ip4(n7111), .op(
        n10399) );
  nor2_1 U8620 ( .ip1(n10994), .ip2(n10399), .op(n7113) );
  not_ab_or_c_or_d U8621 ( .ip1(n11003), .ip2(n10079), .ip3(n7114), .ip4(n7113), .op(n7332) );
  nor2_1 U8622 ( .ip1(n9514), .ip2(n7115), .op(n9362) );
  nor2_1 U8623 ( .ip1(\interconnect_ip_inst/i_ahb_U_mux_hsel_prev [1]), .ip2(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [2]), .op(n7116) );
  nor2_1 U8624 ( .ip1(\interconnect_ip_inst/i_ahb_U_mux_hsel_prev [4]), .ip2(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [3]), .op(n8403) );
  nand3_1 U8625 ( .ip1(n7116), .ip2(n8403), .ip3(
        \interconnect_ip_inst/i_ahb_hresp_none_0_ ), .op(n7117) );
  nand2_1 U8626 ( .ip1(n450), .ip2(n7117), .op(n12602) );
  and2_1 U8627 ( .ip1(n12602), .ip2(n11807), .op(n7327) );
  nor2_1 U8628 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n7118), .op(
        n7119) );
  not_ab_or_c_or_d U8629 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n10587), .ip3(n4150), .ip4(n7119), .op(n7326) );
  inv_1 U8630 ( .ip(n10538), .op(n9934) );
  nor2_1 U8631 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n9934), .op(
        n7723) );
  or2_1 U8632 ( .ip1(\CORTEXM0DS_INST/u_logic/Zph2z4 [0]), .ip2(n7723), .op(
        n7121) );
  inv_1 U8633 ( .ip(n8993), .op(n12082) );
  or2_1 U8634 ( .ip1(n12082), .ip2(n7723), .op(n7120) );
  nand2_1 U8635 ( .ip1(n7121), .ip2(n7120), .op(n7122) );
  or2_1 U8636 ( .ip1(\CORTEXM0DS_INST/u_logic/Zph2z4 [1]), .ip2(n7122), .op(
        n7124) );
  or2_1 U8637 ( .ip1(n4130), .ip2(n7122), .op(n7123) );
  nand2_1 U8638 ( .ip1(n7124), .ip2(n7123), .op(n7129) );
  nand2_1 U8639 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [23]), .ip2(n11609), 
        .op(n7126) );
  nand2_1 U8640 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [23]), .ip2(n11610), 
        .op(n7125) );
  nand3_1 U8641 ( .ip1(n7126), .ip2(n3027), .ip3(n7125), .op(n10416) );
  inv_1 U8642 ( .ip(n10416), .op(n9952) );
  nor4_1 U8643 ( .ip1(\CORTEXM0DS_INST/u_logic/Zph2z4 [0]), .ip2(n9952), .ip3(
        n7127), .ip4(n8993), .op(n7128) );
  nor2_1 U8644 ( .ip1(n7129), .ip2(n7128), .op(n7322) );
  nand2_1 U8645 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [1]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [1]), .op(n7131) );
  nand2_1 U8646 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [0]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [0]), .op(n7130) );
  nand2_1 U8647 ( .ip1(n7131), .ip2(n7130), .op(n7238) );
  nand2_1 U8648 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [3]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [3]), .op(n7133) );
  nand2_1 U8649 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [2]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [2]), .op(n7132) );
  nand2_1 U8650 ( .ip1(n7133), .ip2(n7132), .op(n7237) );
  nor2_1 U8651 ( .ip1(n7238), .ip2(n7237), .op(n7250) );
  inv_1 U8652 ( .ip(n7250), .op(n7138) );
  nand2_1 U8653 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [5]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [5]), .op(n7135) );
  nand2_1 U8654 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [4]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [4]), .op(n7134) );
  nand2_1 U8655 ( .ip1(n7135), .ip2(n7134), .op(n7220) );
  nand2_1 U8656 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [7]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [7]), .op(n7137) );
  nand2_1 U8657 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [6]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [6]), .op(n7136) );
  nand2_1 U8658 ( .ip1(n7137), .ip2(n7136), .op(n7219) );
  or2_1 U8659 ( .ip1(n7220), .ip2(n7219), .op(n7241) );
  nor2_1 U8660 ( .ip1(n7138), .ip2(n7241), .op(n7272) );
  nor2_1 U8661 ( .ip1(n7139), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [23]), .op(
        n7141) );
  not_ab_or_c_or_d U8662 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [23]), .ip2(
        n7139), .ip3(\CORTEXM0DS_INST/u_logic/Zuh2z4 [22]), .ip4(n10204), .op(
        n7140) );
  or2_1 U8663 ( .ip1(n7141), .ip2(n7140), .op(n7142) );
  nand3_1 U8664 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [11]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [11]), .ip3(n7142), .op(n7143) );
  and3_1 U8665 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [10]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [10]), .ip3(n7143), .op(n9887) );
  mux2_1 U8666 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [23]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [21]), .s(n9887), .op(n7152) );
  inv_1 U8667 ( .ip(n7152), .op(n7159) );
  inv_1 U8668 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [19]), .op(n7303) );
  nor2_1 U8669 ( .ip1(n11794), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [19]), 
        .op(n7146) );
  not_ab_or_c_or_d U8670 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [19]), .ip2(
        n11794), .ip3(\CORTEXM0DS_INST/u_logic/Zuh2z4 [18]), .ip4(n7144), .op(
        n7145) );
  or2_1 U8671 ( .ip1(n7146), .ip2(n7145), .op(n7147) );
  nand3_1 U8672 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [9]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [9]), .ip3(n7147), .op(n7148) );
  and3_1 U8673 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [8]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [8]), .ip3(n7148), .op(n9889) );
  mux2_1 U8674 ( .ip1(n7303), .ip2(n11794), .s(n9889), .op(n7158) );
  nand2_1 U8675 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [9]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [9]), .op(n7150) );
  nand2_1 U8676 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [8]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [8]), .op(n7149) );
  nand2_1 U8677 ( .ip1(n7150), .ip2(n7149), .op(n7189) );
  nor2_1 U8678 ( .ip1(n7152), .ip2(n7158), .op(n7154) );
  mux2_1 U8679 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [18]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [16]), .s(n9889), .op(n7182) );
  inv_1 U8680 ( .ip(n7182), .op(n7151) );
  mux2_1 U8681 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [22]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [20]), .s(n9887), .op(n7183) );
  not_ab_or_c_or_d U8682 ( .ip1(n7158), .ip2(n7152), .ip3(n7151), .ip4(n7183), 
        .op(n7153) );
  or2_1 U8683 ( .ip1(n7154), .ip2(n7153), .op(n7157) );
  nand2_1 U8684 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [11]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [11]), .op(n7156) );
  nand2_1 U8685 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [10]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [10]), .op(n7155) );
  nand2_1 U8686 ( .ip1(n7156), .ip2(n7155), .op(n7190) );
  nand2_1 U8687 ( .ip1(n7157), .ip2(n7190), .op(n9888) );
  and2_1 U8688 ( .ip1(n7189), .ip2(n9888), .op(n7734) );
  mux2_1 U8689 ( .ip1(n7159), .ip2(n7158), .s(n7734), .op(n7198) );
  inv_1 U8690 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [29]), .op(n7160) );
  nor2_1 U8691 ( .ip1(n7160), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [31]), .op(
        n7162) );
  not_ab_or_c_or_d U8692 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [31]), .ip2(
        n7160), .ip3(\CORTEXM0DS_INST/u_logic/Zuh2z4 [30]), .ip4(n10202), .op(
        n7161) );
  or2_1 U8693 ( .ip1(n7162), .ip2(n7161), .op(n7163) );
  nand3_1 U8694 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [15]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [15]), .ip3(n7163), .op(n7164) );
  and3_1 U8695 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [14]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [14]), .ip3(n7164), .op(n9880) );
  mux2_1 U8696 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [31]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [29]), .s(n9880), .op(n7181) );
  inv_1 U8697 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [25]), .op(n11789) );
  nor2_1 U8698 ( .ip1(n11789), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [27]), 
        .op(n7166) );
  not_ab_or_c_or_d U8699 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [27]), .ip2(
        n11789), .ip3(\CORTEXM0DS_INST/u_logic/Zuh2z4 [26]), .ip4(n10186), 
        .op(n7165) );
  or2_1 U8700 ( .ip1(n7166), .ip2(n7165), .op(n7167) );
  nand3_1 U8701 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [13]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [13]), .ip3(n7167), .op(n7168) );
  nand3_1 U8702 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [12]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [12]), .ip3(n7168), .op(n9882) );
  mux2_1 U8703 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [25]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [27]), .s(n9882), .op(n7180) );
  inv_1 U8704 ( .ip(n7180), .op(n7170) );
  nor2_1 U8705 ( .ip1(n7181), .ip2(n7170), .op(n7172) );
  mux2_1 U8706 ( .ip1(n10186), .ip2(n7169), .s(n9882), .op(n7185) );
  mux2_1 U8707 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [30]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [28]), .s(n9880), .op(n7264) );
  not_ab_or_c_or_d U8708 ( .ip1(n7170), .ip2(n7181), .ip3(n7185), .ip4(n7264), 
        .op(n7171) );
  or2_1 U8709 ( .ip1(n7172), .ip2(n7171), .op(n7175) );
  and2_1 U8710 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [13]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [13]), .op(n7174) );
  and2_1 U8711 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [12]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [12]), .op(n7173) );
  nor2_1 U8712 ( .ip1(n7174), .ip2(n7173), .op(n7193) );
  or2_1 U8713 ( .ip1(n7175), .ip2(n7193), .op(n7179) );
  nand2_1 U8714 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [15]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [15]), .op(n7177) );
  nand2_1 U8715 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [14]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [14]), .op(n7176) );
  nand2_1 U8716 ( .ip1(n7177), .ip2(n7176), .op(n7194) );
  or2_1 U8717 ( .ip1(n7194), .ip2(n7193), .op(n7178) );
  nand2_1 U8718 ( .ip1(n7179), .ip2(n7178), .op(n9883) );
  mux2_1 U8719 ( .ip1(n7181), .ip2(n7180), .s(n9883), .op(n7196) );
  mux2_1 U8720 ( .ip1(n7183), .ip2(n7182), .s(n7734), .op(n7261) );
  inv_1 U8721 ( .ip(n7261), .op(n7188) );
  inv_1 U8722 ( .ip(n7264), .op(n7184) );
  nand2_1 U8723 ( .ip1(n7194), .ip2(n7184), .op(n7186) );
  inv_1 U8724 ( .ip(n7185), .op(n7260) );
  mux2_1 U8725 ( .ip1(n7186), .ip2(n7260), .s(n9883), .op(n7187) );
  not_ab_or_c_or_d U8726 ( .ip1(n7198), .ip2(n7196), .ip3(n7188), .ip4(n7187), 
        .op(n7192) );
  nor2_1 U8727 ( .ip1(n7190), .ip2(n7189), .op(n7191) );
  or2_1 U8728 ( .ip1(n7192), .ip2(n7191), .op(n7257) );
  nand2_1 U8729 ( .ip1(n7257), .ip2(n7196), .op(n7200) );
  inv_1 U8730 ( .ip(n7193), .op(n7195) );
  nor2_1 U8731 ( .ip1(n7195), .ip2(n7194), .op(n7256) );
  nor3_1 U8732 ( .ip1(n7198), .ip2(n7196), .ip3(n7256), .op(n7197) );
  nor2_1 U8733 ( .ip1(n7197), .ip2(n7257), .op(n10138) );
  inv_1 U8734 ( .ip(n10138), .op(n7733) );
  or2_1 U8735 ( .ip1(n7733), .ip2(n7198), .op(n7199) );
  nand2_1 U8736 ( .ip1(n7200), .ip2(n7199), .op(n7273) );
  nor2_1 U8737 ( .ip1(n7202), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [15]), .op(
        n7204) );
  not_ab_or_c_or_d U8738 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [15]), .ip2(
        n7202), .ip3(\CORTEXM0DS_INST/u_logic/Zuh2z4 [14]), .ip4(n7201), .op(
        n7203) );
  or2_1 U8739 ( .ip1(n7204), .ip2(n7203), .op(n7205) );
  nand3_1 U8740 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [7]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [7]), .ip3(n7205), .op(n7206) );
  and3_1 U8741 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [6]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [6]), .ip3(n7206), .op(n9902) );
  mux2_1 U8742 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [15]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [13]), .s(n9902), .op(n7222) );
  inv_1 U8743 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [9]), .op(n7212) );
  nor2_1 U8744 ( .ip1(n7212), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [11]), .op(
        n7209) );
  inv_1 U8745 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [8]), .op(n7207) );
  not_ab_or_c_or_d U8746 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [11]), .ip2(
        n7212), .ip3(\CORTEXM0DS_INST/u_logic/Zuh2z4 [10]), .ip4(n7207), .op(
        n7208) );
  or2_1 U8747 ( .ip1(n7209), .ip2(n7208), .op(n7210) );
  nand3_1 U8748 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [5]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [5]), .ip3(n7210), .op(n7211) );
  and3_1 U8749 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [4]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [4]), .ip3(n7211), .op(n9893) );
  mux2_1 U8750 ( .ip1(n7213), .ip2(n7212), .s(n9893), .op(n7215) );
  inv_1 U8751 ( .ip(n7215), .op(n7221) );
  nor2_1 U8752 ( .ip1(n7222), .ip2(n7215), .op(n7217) );
  mux2_1 U8753 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [10]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [8]), .s(n9893), .op(n7244) );
  inv_1 U8754 ( .ip(n7244), .op(n7214) );
  mux2_1 U8755 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [14]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [12]), .s(n9902), .op(n7245) );
  not_ab_or_c_or_d U8756 ( .ip1(n7215), .ip2(n7222), .ip3(n7214), .ip4(n7245), 
        .op(n7216) );
  or2_1 U8757 ( .ip1(n7217), .ip2(n7216), .op(n7218) );
  nand2_1 U8758 ( .ip1(n7219), .ip2(n7218), .op(n9892) );
  and2_1 U8759 ( .ip1(n7220), .ip2(n9892), .op(n7731) );
  mux2_1 U8760 ( .ip1(n7222), .ip2(n7221), .s(n7731), .op(n7255) );
  nor2_1 U8761 ( .ip1(n11796), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [3]), .op(
        n7225) );
  not_ab_or_c_or_d U8762 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [3]), .ip2(
        n11796), .ip3(\CORTEXM0DS_INST/u_logic/Zuh2z4 [2]), .ip4(n7223), .op(
        n7224) );
  or2_1 U8763 ( .ip1(n7225), .ip2(n7224), .op(n7226) );
  nand3_1 U8764 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [1]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [1]), .ip3(n7226), .op(n7227) );
  and3_1 U8765 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [0]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [0]), .ip3(n7227), .op(n9896) );
  mux2_1 U8766 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [3]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [1]), .s(n9896), .op(n7240) );
  inv_1 U8767 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [5]), .op(n11813) );
  nor2_1 U8768 ( .ip1(n11813), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [7]), .op(
        n7229) );
  inv_1 U8769 ( .ip(\CORTEXM0DS_INST/u_logic/Zuh2z4 [4]), .op(n10203) );
  not_ab_or_c_or_d U8770 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [7]), .ip2(
        n11813), .ip3(\CORTEXM0DS_INST/u_logic/Zuh2z4 [6]), .ip4(n10203), .op(
        n7228) );
  or2_1 U8771 ( .ip1(n7229), .ip2(n7228), .op(n7230) );
  nand3_1 U8772 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [3]), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [3]), .ip3(n7230), .op(n7231) );
  and3_1 U8773 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [2]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [2]), .ip3(n7231), .op(n9891) );
  mux2_1 U8774 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [7]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [5]), .s(n9891), .op(n7239) );
  inv_1 U8775 ( .ip(n7240), .op(n7233) );
  nor2_1 U8776 ( .ip1(n7239), .ip2(n7233), .op(n7235) );
  mux2_1 U8777 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [2]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [0]), .s(n9896), .op(n7243) );
  inv_1 U8778 ( .ip(n7243), .op(n7232) );
  mux2_1 U8779 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [6]), .ip2(
        \CORTEXM0DS_INST/u_logic/Zuh2z4 [4]), .s(n9891), .op(n7242) );
  not_ab_or_c_or_d U8780 ( .ip1(n7233), .ip2(n7239), .ip3(n7232), .ip4(n7242), 
        .op(n7234) );
  or2_1 U8781 ( .ip1(n7235), .ip2(n7234), .op(n7236) );
  nand2_1 U8782 ( .ip1(n7237), .ip2(n7236), .op(n9894) );
  nand2_1 U8783 ( .ip1(n7238), .ip2(n9894), .op(n9890) );
  mux2_1 U8784 ( .ip1(n7240), .ip2(n7239), .s(n9890), .op(n7254) );
  or2_1 U8785 ( .ip1(n7241), .ip2(n7250), .op(n7253) );
  inv_1 U8786 ( .ip(n7254), .op(n7247) );
  nor2_1 U8787 ( .ip1(n7255), .ip2(n7247), .op(n7249) );
  mux2_1 U8788 ( .ip1(n7243), .ip2(n7242), .s(n9890), .op(n7258) );
  inv_1 U8789 ( .ip(n7258), .op(n7246) );
  mux2_1 U8790 ( .ip1(n7245), .ip2(n7244), .s(n7731), .op(n7259) );
  not_ab_or_c_or_d U8791 ( .ip1(n7247), .ip2(n7255), .ip3(n7246), .ip4(n7259), 
        .op(n7248) );
  or2_1 U8792 ( .ip1(n7249), .ip2(n7248), .op(n7251) );
  or2_1 U8793 ( .ip1(n7251), .ip2(n7250), .op(n7252) );
  nand2_1 U8794 ( .ip1(n7253), .ip2(n7252), .op(n9895) );
  mux2_1 U8795 ( .ip1(n7255), .ip2(n7254), .s(n9895), .op(n7274) );
  inv_1 U8796 ( .ip(n7274), .op(n7268) );
  and2_1 U8797 ( .ip1(n7257), .ip2(n7256), .op(n7271) );
  nor3_1 U8798 ( .ip1(n7273), .ip2(n7268), .ip3(n7271), .op(n7270) );
  mux2_1 U8799 ( .ip1(n7259), .ip2(n7258), .s(n9895), .op(n7277) );
  nor2_1 U8800 ( .ip1(n9883), .ip2(n10138), .op(n7735) );
  and2_1 U8801 ( .ip1(n7260), .ip2(n9883), .op(n7262) );
  mux2_1 U8802 ( .ip1(n7262), .ip2(n7261), .s(n10138), .op(n7263) );
  or2_1 U8803 ( .ip1(n7735), .ip2(n7263), .op(n7266) );
  or2_1 U8804 ( .ip1(n7264), .ip2(n7263), .op(n7265) );
  nand2_1 U8805 ( .ip1(n7266), .ip2(n7265), .op(n7275) );
  nand2_1 U8806 ( .ip1(n7277), .ip2(n7275), .op(n7267) );
  not_ab_or_c_or_d U8807 ( .ip1(n7268), .ip2(n7273), .ip3(n7271), .ip4(n7267), 
        .op(n7269) );
  or2_1 U8808 ( .ip1(n7270), .ip2(n7269), .op(n10137) );
  nor2_1 U8809 ( .ip1(n7272), .ip2(n10137), .op(n9884) );
  nor2_1 U8810 ( .ip1(\CORTEXM0DS_INST/u_logic/Krgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Eqgvx4 ), .op(n8596) );
  nor2_1 U8811 ( .ip1(\CORTEXM0DS_INST/u_logic/Qsgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Wtgvx4 ), .op(n7298) );
  nand2_1 U8812 ( .ip1(n7272), .ip2(n7271), .op(n7283) );
  nor2_1 U8813 ( .ip1(\CORTEXM0DS_INST/u_logic/R3hvx4 ), .ip2(n7283), .op(
        n7294) );
  nand2_1 U8814 ( .ip1(n7298), .ip2(n7294), .op(n9879) );
  nand2_1 U8815 ( .ip1(n8596), .ip2(n9879), .op(n12440) );
  or2_1 U8816 ( .ip1(n9884), .ip2(n12440), .op(n7301) );
  inv_1 U8817 ( .ip(n9884), .op(n10140) );
  mux2_1 U8818 ( .ip1(n7274), .ip2(n7273), .s(n10140), .op(n7284) );
  inv_1 U8819 ( .ip(\CORTEXM0DS_INST/u_logic/Txh2z4 [1]), .op(n7278) );
  nor2_1 U8820 ( .ip1(n7284), .ip2(n7278), .op(n7280) );
  inv_1 U8821 ( .ip(n7275), .op(n7276) );
  mux2_1 U8822 ( .ip1(n7277), .ip2(n7276), .s(n10140), .op(n7291) );
  inv_1 U8823 ( .ip(\CORTEXM0DS_INST/u_logic/Txh2z4 [0]), .op(n10170) );
  not_ab_or_c_or_d U8824 ( .ip1(n7278), .ip2(n7284), .ip3(n7291), .ip4(n10170), 
        .op(n7279) );
  or2_1 U8825 ( .ip1(n7280), .ip2(n7279), .op(n7281) );
  inv_1 U8826 ( .ip(\CORTEXM0DS_INST/u_logic/R3hvx4 ), .op(n11690) );
  or2_1 U8827 ( .ip1(n7281), .ip2(n11690), .op(n7282) );
  nand2_1 U8828 ( .ip1(n7283), .ip2(n7282), .op(n7299) );
  mux2_1 U8829 ( .ip1(n7284), .ip2(\CORTEXM0DS_INST/u_logic/Txh2z4 [1]), .s(
        n7299), .op(n8582) );
  inv_1 U8830 ( .ip(\CORTEXM0DS_INST/u_logic/Uth2z4 [1]), .op(n11828) );
  inv_1 U8831 ( .ip(\CORTEXM0DS_INST/u_logic/Wtgvx4 ), .op(n11852) );
  or2_1 U8832 ( .ip1(\CORTEXM0DS_INST/u_logic/Qsgvx4 ), .ip2(n11852), .op(
        n7289) );
  nor2_1 U8833 ( .ip1(n11828), .ip2(\CORTEXM0DS_INST/u_logic/Psh2z4 [1]), .op(
        n7286) );
  inv_1 U8834 ( .ip(\CORTEXM0DS_INST/u_logic/Uth2z4 [0]), .op(n10167) );
  not_ab_or_c_or_d U8835 ( .ip1(\CORTEXM0DS_INST/u_logic/Psh2z4 [1]), .ip2(
        n11828), .ip3(\CORTEXM0DS_INST/u_logic/Psh2z4 [0]), .ip4(n10167), .op(
        n7285) );
  or2_1 U8836 ( .ip1(n7286), .ip2(n7285), .op(n7287) );
  or2_1 U8837 ( .ip1(n7287), .ip2(n11852), .op(n7288) );
  nand2_1 U8838 ( .ip1(n7289), .ip2(n7288), .op(n10146) );
  mux2_1 U8839 ( .ip1(n7290), .ip2(n11828), .s(n10146), .op(n8583) );
  nor3_1 U8840 ( .ip1(n8582), .ip2(n8583), .ip3(n7294), .op(n7296) );
  inv_1 U8841 ( .ip(n7291), .op(n7292) );
  mux2_1 U8842 ( .ip1(n7292), .ip2(n10170), .s(n7299), .op(n8578) );
  mux2_1 U8843 ( .ip1(\CORTEXM0DS_INST/u_logic/Psh2z4 [0]), .ip2(
        \CORTEXM0DS_INST/u_logic/Uth2z4 [0]), .s(n10146), .op(n8581) );
  nand2_1 U8844 ( .ip1(n8578), .ip2(n8581), .op(n7293) );
  not_ab_or_c_or_d U8845 ( .ip1(n8583), .ip2(n8582), .ip3(n7294), .ip4(n7293), 
        .op(n7295) );
  nor2_1 U8846 ( .ip1(n7296), .ip2(n7295), .op(n10145) );
  inv_1 U8847 ( .ip(n10145), .op(n7297) );
  nor2_1 U8848 ( .ip1(n7298), .ip2(n7297), .op(n9910) );
  nor2_1 U8849 ( .ip1(n7299), .ip2(n9910), .op(n9903) );
  or2_1 U8850 ( .ip1(n9903), .ip2(n12440), .op(n7300) );
  nand2_1 U8851 ( .ip1(n7301), .ip2(n7300), .op(n12465) );
  nand3_1 U8852 ( .ip1(\CORTEXM0DS_INST/u_logic/N6hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Xahvx4 ), .ip3(n12682), .op(n11825) );
  nor2_1 U8853 ( .ip1(n11839), .ip2(n11825), .op(n10152) );
  inv_1 U8854 ( .ip(n8536), .op(n11799) );
  and2_1 U8855 ( .ip1(n11866), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [15]), 
        .op(n7313) );
  nand4_1 U8856 ( .ip1(\CORTEXM0DS_INST/u_logic/N6hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Z7hvx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/B5hvx4 ), .ip4(n10208), .op(n7302) );
  nor2_1 U8857 ( .ip1(\CORTEXM0DS_INST/u_logic/Xahvx4 ), .ip2(n7302), .op(
        n11824) );
  nand2_1 U8858 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [3]), .ip2(n11824), 
        .op(n7311) );
  nor2_1 U8859 ( .ip1(n11865), .ip2(n7302), .op(n11833) );
  nor2_1 U8860 ( .ip1(\CORTEXM0DS_INST/u_logic/Xahvx4 ), .ip2(n7305), .op(
        n8540) );
  inv_1 U8861 ( .ip(n8540), .op(n10207) );
  nor3_1 U8862 ( .ip1(n10208), .ip2(n7304), .ip3(n10207), .op(n11827) );
  inv_1 U8863 ( .ip(n11827), .op(n11795) );
  nor2_1 U8864 ( .ip1(n7303), .ip2(n11795), .op(n7308) );
  nor4_1 U8865 ( .ip1(n7305), .ip2(n11865), .ip3(n10208), .ip4(n7304), .op(
        n11823) );
  inv_1 U8866 ( .ip(n11823), .op(n11790) );
  nor2_1 U8867 ( .ip1(n7306), .ip2(n11790), .op(n7307) );
  not_ab_or_c_or_d U8868 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [11]), .ip2(
        n11833), .ip3(n7308), .ip4(n7307), .op(n7310) );
  nand2_1 U8869 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [15]), .ip2(n11800), 
        .op(n7309) );
  nand3_1 U8870 ( .ip1(n7311), .ip2(n7310), .ip3(n7309), .op(n7312) );
  not_ab_or_c_or_d U8871 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [15]), .ip2(
        n11799), .ip3(n7313), .ip4(n7312), .op(n7314) );
  nor2_1 U8872 ( .ip1(n7314), .ip2(n11839), .op(n7319) );
  inv_1 U8873 ( .ip(n7315), .op(n9376) );
  mux2_1 U8874 ( .ip1(n7316), .ip2(n9376), .s(n9443), .op(n7317) );
  inv_1 U8875 ( .ip(n7317), .op(n9470) );
  nor2_1 U8876 ( .ip1(n9470), .ip2(n11811), .op(n7318) );
  not_ab_or_c_or_d U8877 ( .ip1(n12465), .ip2(n10152), .ip3(n7319), .ip4(n7318), .op(n7320) );
  nand2_1 U8878 ( .ip1(n3002), .ip2(n7320), .op(n10414) );
  nor2_1 U8879 ( .ip1(\CORTEXM0DS_INST/u_logic/Zph2z4 [1]), .ip2(n10414), .op(
        n7321) );
  or2_1 U8880 ( .ip1(n7322), .ip2(n7321), .op(n7324) );
  nand2_1 U8881 ( .ip1(n10414), .ip2(n9748), .op(n7323) );
  nand2_1 U8882 ( .ip1(n7324), .ip2(n7323), .op(n7325) );
  nor4_1 U8883 ( .ip1(n9362), .ip2(n7327), .ip3(n7326), .ip4(n7325), .op(n9871) );
  nor2_1 U8884 ( .ip1(n9933), .ip2(n7327), .op(n7802) );
  nor2_1 U8885 ( .ip1(n7328), .ip2(n7800), .op(n7329) );
  inv_1 U8886 ( .ip(n9469), .op(n9485) );
  nor2_1 U8887 ( .ip1(n7329), .ip2(n9485), .op(n7799) );
  nor2_1 U8888 ( .ip1(n7799), .ip2(n10047), .op(n7330) );
  nor4_1 U8889 ( .ip1(n9871), .ip2(n7802), .ip3(n7331), .ip4(n7330), .op(
        n11002) );
  inv_1 U8890 ( .ip(n11002), .op(n10371) );
  nand3_1 U8891 ( .ip1(n7333), .ip2(n7332), .ip3(n10371), .op(n11388) );
  nand2_1 U8892 ( .ip1(n10859), .ip2(n11388), .op(n7334) );
  nand4_1 U8893 ( .ip1(n10573), .ip2(n7336), .ip3(n7335), .ip4(n7334), .op(
        \CORTEXM0DS_INST/u_logic/Bmhvx4 ) );
  nand2_1 U8894 ( .ip1(\CORTEXM0DS_INST/u_logic/E1dvx4 ), .ip2(n2120), .op(
        n7348) );
  nand2_1 U8895 ( .ip1(\CORTEXM0DS_INST/vis_pc [1]), .ip2(n12321), .op(n7347)
         );
  nand2_1 U8896 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [2]), .ip2(n12320), .op(n7346) );
  inv_1 U8897 ( .ip(n9180), .op(n11718) );
  nand2_1 U8898 ( .ip1(n11718), .ip2(n12314), .op(n7344) );
  xor2_1 U8899 ( .ip1(n7338), .ip2(n7337), .op(n10392) );
  nand2_1 U8900 ( .ip1(n10392), .ip2(n12300), .op(n7343) );
  or2_1 U8901 ( .ip1(n7339), .ip2(\CORTEXM0DS_INST/vis_pc [1]), .op(n7341) );
  nand3_1 U8902 ( .ip1(n12599), .ip2(n7341), .ip3(n7340), .op(n7342) );
  nand3_1 U8903 ( .ip1(n7344), .ip2(n7343), .ip3(n7342), .op(n1851) );
  nand2_1 U8904 ( .ip1(n12691), .ip2(n1851), .op(n7345) );
  nand4_1 U8905 ( .ip1(n7348), .ip2(n7347), .ip3(n7346), .ip4(n7345), .op(
        n6081) );
  nand2_1 U8906 ( .ip1(\CORTEXM0DS_INST/vis_pc [3]), .ip2(n12321), .op(n7391)
         );
  nand2_1 U8907 ( .ip1(\CORTEXM0DS_INST/u_logic/Y3dvx4 ), .ip2(n2120), .op(
        n7390) );
  nand2_1 U8908 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [4]), .ip2(n12320), .op(n7389) );
  nand2_1 U8909 ( .ip1(\CORTEXM0DS_INST/u_logic/P39vx4 ), .ip2(n8295), .op(
        n7364) );
  nand2_1 U8910 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(n7670), .op(
        n7363) );
  inv_1 U8911 ( .ip(\CORTEXM0DS_INST/cm0_r10 [4]), .op(n7366) );
  nor2_1 U8912 ( .ip1(n7349), .ip2(n7366), .op(n7351) );
  and2_1 U8913 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [2]), .op(n7350)
         );
  not_ab_or_c_or_d U8914 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [4]), .ip2(n8914), 
        .ip3(n7351), .ip4(n7350), .op(n7360) );
  nand2_1 U8915 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [4]), .ip2(n8910), .op(n7354)
         );
  nand2_1 U8916 ( .ip1(n8853), .ip2(\CORTEXM0DS_INST/u_logic/Y3dvx4 ), .op(
        n7353) );
  nand2_1 U8917 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [4]), .op(n7352)
         );
  nand3_1 U8918 ( .ip1(n7354), .ip2(n7353), .ip3(n7352), .op(n7355) );
  not_ab_or_c_or_d U8919 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [4]), 
        .ip3(n7356), .ip4(n7355), .op(n7359) );
  nand2_1 U8920 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [2]), .op(n7358)
         );
  nand2_1 U8921 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [4]), .op(n7357)
         );
  nand2_1 U8922 ( .ip1(n8011), .ip2(n12671), .op(n7362) );
  nand2_1 U8923 ( .ip1(\CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip2(n7682), .op(
        n7361) );
  mux2_1 U8924 ( .ip1(n8013), .ip2(n8297), .s(n7365), .op(n9169) );
  and2_1 U8925 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [4]), .op(n7379)
         );
  nor2_1 U8926 ( .ip1(n7367), .ip2(n7366), .op(n7373) );
  nand2_1 U8927 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [2]), .op(n7371)
         );
  nand2_1 U8928 ( .ip1(n8946), .ip2(n9264), .op(n7370) );
  nand2_1 U8929 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/Y3dvx4 ), .op(
        n7369) );
  nand2_1 U8930 ( .ip1(\CORTEXM0DS_INST/u_logic/O2dvx4 ), .ip2(n8948), .op(
        n7368) );
  not_ab_or_c_or_d U8931 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [4]), .ip2(n8957), 
        .ip3(n7373), .ip4(n7372), .op(n7377) );
  nand2_1 U8932 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [4]), .op(n7376)
         );
  nand2_1 U8933 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [4]), .op(n7375)
         );
  nand2_1 U8934 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [2]), .op(n7374)
         );
  nand4_1 U8935 ( .ip1(n7377), .ip2(n7376), .ip3(n7375), .ip4(n7374), .op(
        n7378) );
  not_ab_or_c_or_d U8936 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [4]), .ip2(n8966), 
        .ip3(n7379), .ip4(n7378), .op(n9174) );
  nor2_1 U8937 ( .ip1(n8974), .ip2(n9174), .op(n7701) );
  fulladder U8938 ( .a(n9066), .b(n7381), .ci(n7380), .co(n7700), .s(n6940) );
  nor2_1 U8939 ( .ip1(n7383), .ip2(n7382), .op(n7715) );
  xor2_1 U8940 ( .ip1(n7716), .ip2(n7715), .op(n11397) );
  inv_1 U8941 ( .ip(n7384), .op(n7385) );
  inv_1 U8942 ( .ip(\CORTEXM0DS_INST/vis_pc [3]), .op(n10376) );
  nor2_1 U8943 ( .ip1(n7385), .ip2(n10376), .op(n12226) );
  not_ab_or_c_or_d U8944 ( .ip1(n7385), .ip2(n10376), .ip3(n12226), .ip4(
        n12305), .op(n7387) );
  nor2_1 U8945 ( .ip1(n9174), .ip2(n12295), .op(n7386) );
  not_ab_or_c_or_d U8946 ( .ip1(n12300), .ip2(n11397), .ip3(n7387), .ip4(n7386), .op(\CORTEXM0DS_INST/u_logic/Yuovx4 ) );
  inv_1 U8947 ( .ip(\CORTEXM0DS_INST/u_logic/Yuovx4 ), .op(n1944) );
  nand2_1 U8948 ( .ip1(n12691), .ip2(n1944), .op(n7388) );
  nand4_1 U8949 ( .ip1(n7391), .ip2(n7390), .ip3(n7389), .ip4(n7388), .op(
        n6090) );
  inv_1 U8950 ( .ip(\CORTEXM0DS_INST/vis_pc [10]), .op(n12133) );
  nand4_1 U8951 ( .ip1(\CORTEXM0DS_INST/vis_pc [9]), .ip2(
        \CORTEXM0DS_INST/vis_pc [11]), .ip3(\CORTEXM0DS_INST/vis_pc [7]), 
        .ip4(\CORTEXM0DS_INST/vis_pc [8]), .op(n9802) );
  nor2_1 U8952 ( .ip1(n12133), .ip2(n9802), .op(n8394) );
  inv_1 U8953 ( .ip(\CORTEXM0DS_INST/vis_pc [5]), .op(n12244) );
  nor3_1 U8954 ( .ip1(n7392), .ip2(n8537), .ip3(n10376), .op(n7393) );
  nand3_1 U8955 ( .ip1(\CORTEXM0DS_INST/vis_pc [1]), .ip2(
        \CORTEXM0DS_INST/vis_pc [4]), .ip3(n7393), .op(n10350) );
  nor2_1 U8956 ( .ip1(n12244), .ip2(n10350), .op(n10349) );
  nand2_1 U8957 ( .ip1(\CORTEXM0DS_INST/vis_pc [6]), .ip2(n10349), .op(n10335)
         );
  inv_1 U8958 ( .ip(n5822), .op(n10860) );
  nand2_1 U8959 ( .ip1(n12091), .ip2(n10860), .op(n10861) );
  nor2_1 U8960 ( .ip1(n10335), .ip2(n10861), .op(n10319) );
  nand2_1 U8961 ( .ip1(n8394), .ip2(n10319), .op(n7394) );
  nand2_1 U8962 ( .ip1(n12091), .ip2(n7394), .op(n10302) );
  mux2_1 U8963 ( .ip1(n7394), .ip2(n10302), .s(\CORTEXM0DS_INST/vis_pc [12]), 
        .op(n7810) );
  nor2_1 U8964 ( .ip1(n12376), .ip2(n7823), .op(n8294) );
  nand2_1 U8965 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [13]), .op(n7397)
         );
  nand2_1 U8966 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [13]), .op(n7396)
         );
  nand2_1 U8967 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [13]), .op(n7395)
         );
  nand3_1 U8968 ( .ip1(n7397), .ip2(n7396), .ip3(n7395), .op(n7414) );
  nand2_1 U8969 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [13]), .ip2(n8925), .op(n7412)
         );
  nand2_1 U8970 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [13]), .op(n7401)
         );
  nand2_1 U8971 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [13]), .op(n7400)
         );
  nand2_1 U8972 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [13]), .op(n7399)
         );
  nand2_1 U8973 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [13]), .op(n7398)
         );
  nand2_1 U8974 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [11]), .op(n7405)
         );
  nand2_1 U8975 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [11]), .op(n7404)
         );
  nand2_1 U8976 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [13]), .op(n7403)
         );
  nand2_1 U8977 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [13]), .op(n7402)
         );
  not_ab_or_c_or_d U8978 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [13]), 
        .ip3(n7407), .ip4(n7406), .op(n7411) );
  and2_1 U8979 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [13]), .op(n7409)
         );
  inv_1 U8980 ( .ip(\CORTEXM0DS_INST/u_logic/Ngdvx4 ), .op(n8298) );
  nor2_1 U8981 ( .ip1(n8909), .ip2(n8298), .op(n7408) );
  not_ab_or_c_or_d U8982 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [13]), .ip2(n8917), 
        .ip3(n7409), .ip4(n7408), .op(n7410) );
  nand3_1 U8983 ( .ip1(n7412), .ip2(n7411), .ip3(n7410), .op(n7413) );
  not_ab_or_c_or_d U8984 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [13]), 
        .ip3(n7414), .ip4(n7413), .op(n11285) );
  nor2_1 U8985 ( .ip1(n11285), .ip2(n8292), .op(n7415) );
  not_ab_or_c_or_d U8986 ( .ip1(\CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip2(n8295), 
        .ip3(n8294), .ip4(n7415), .op(n7416) );
  mux2_1 U8987 ( .ip1(n8297), .ip2(n8013), .s(n7416), .op(n9137) );
  and2_1 U8988 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [13]), .op(n7428)
         );
  and2_1 U8989 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [13]), .op(n7422)
         );
  nand2_1 U8990 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [11]), .op(n7420)
         );
  inv_1 U8991 ( .ip(n9417), .op(n9270) );
  nand2_1 U8992 ( .ip1(n8946), .ip2(n9270), .op(n7419) );
  nand2_1 U8993 ( .ip1(\CORTEXM0DS_INST/u_logic/Cfdvx4 ), .ip2(n8948), .op(
        n7418) );
  nand2_1 U8994 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/Ngdvx4 ), .op(
        n7417) );
  not_ab_or_c_or_d U8995 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [13]), .ip2(n8956), 
        .ip3(n7422), .ip4(n7421), .op(n7426) );
  nand2_1 U8996 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [13]), .op(n7425)
         );
  nand2_1 U8997 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [13]), .op(n7424)
         );
  nand2_1 U8998 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [11]), .op(n7423)
         );
  nand4_1 U8999 ( .ip1(n7426), .ip2(n7425), .ip3(n7424), .ip4(n7423), .op(
        n7427) );
  not_ab_or_c_or_d U9000 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [13]), .ip2(n8966), 
        .ip3(n7428), .ip4(n7427), .op(n9804) );
  nor2_1 U9001 ( .ip1(n8974), .ip2(n9804), .op(n8312) );
  nand2_1 U9002 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [12]), .op(n7431)
         );
  nand2_1 U9003 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [12]), .op(n7430)
         );
  nand2_1 U9004 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [12]), .op(n7429)
         );
  nand3_1 U9005 ( .ip1(n7431), .ip2(n7430), .ip3(n7429), .op(n7450) );
  inv_1 U9006 ( .ip(\CORTEXM0DS_INST/u_logic/Cfdvx4 ), .op(n12148) );
  nor2_1 U9007 ( .ip1(n8909), .ip2(n12148), .op(n7432) );
  or2_1 U9008 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [12]), .ip2(n7432), .op(n7434)
         );
  or2_1 U9009 ( .ip1(n8915), .ip2(n7432), .op(n7433) );
  nand2_1 U9010 ( .ip1(n7434), .ip2(n7433), .op(n7448) );
  nand2_1 U9011 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [12]), .op(n7438)
         );
  nand2_1 U9012 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [12]), .op(n7437)
         );
  nand2_1 U9013 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [12]), .op(n7436)
         );
  nand2_1 U9014 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [12]), .op(n7435)
         );
  nand2_1 U9015 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [10]), .op(n7442)
         );
  nand2_1 U9016 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [10]), .op(n7441)
         );
  nand2_1 U9017 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [12]), .op(n7440)
         );
  nand2_1 U9018 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [12]), .op(n7439)
         );
  not_ab_or_c_or_d U9019 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [12]), 
        .ip3(n7444), .ip4(n7443), .op(n7447) );
  nand2_1 U9020 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [12]), .op(n7446)
         );
  nand2_1 U9021 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [12]), .op(n7445)
         );
  not_ab_or_c_or_d U9022 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [12]), 
        .ip3(n7450), .ip4(n7449), .op(n11269) );
  nor2_1 U9023 ( .ip1(n11269), .ip2(n8292), .op(n7451) );
  not_ab_or_c_or_d U9024 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n8295), 
        .ip3(n8294), .ip4(n7451), .op(n7452) );
  mux2_1 U9025 ( .ip1(n8297), .ip2(n8013), .s(n7452), .op(n9143) );
  and2_1 U9026 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [12]), .op(n7464)
         );
  and2_1 U9027 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [12]), .op(n7458)
         );
  nand2_1 U9028 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [10]), .op(n7456)
         );
  nand2_1 U9029 ( .ip1(n8946), .ip2(n9269), .op(n7455) );
  nand2_1 U9030 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/Cfdvx4 ), .op(
        n7454) );
  nand2_1 U9031 ( .ip1(\CORTEXM0DS_INST/u_logic/Rddvx4 ), .ip2(n8948), .op(
        n7453) );
  not_ab_or_c_or_d U9032 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [12]), .ip2(n8966), 
        .ip3(n7458), .ip4(n7457), .op(n7462) );
  nand2_1 U9033 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [12]), .op(n7461)
         );
  nand2_1 U9034 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [12]), .op(n7460)
         );
  nand2_1 U9035 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [10]), .op(n7459)
         );
  nand4_1 U9036 ( .ip1(n7462), .ip2(n7461), .ip3(n7460), .ip4(n7459), .op(
        n7463) );
  not_ab_or_c_or_d U9037 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [12]), .ip2(n8944), 
        .ip3(n7464), .ip4(n7463), .op(n12141) );
  nor2_1 U9038 ( .ip1(n8974), .ip2(n12141), .op(n7722) );
  nand2_1 U9039 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [11]), .op(n7467)
         );
  nand2_1 U9040 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [11]), .op(n7466)
         );
  nand2_1 U9041 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [11]), .op(n7465)
         );
  nand3_1 U9042 ( .ip1(n7467), .ip2(n7466), .ip3(n7465), .op(n7484) );
  nand2_1 U9043 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [11]), .ip2(n8902), .op(n7482)
         );
  nand2_1 U9044 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [11]), .op(n7471)
         );
  nand2_1 U9045 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [11]), .op(n7470)
         );
  nand2_1 U9046 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [11]), .op(n7469)
         );
  nand2_1 U9047 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [11]), .op(n7468)
         );
  nand2_1 U9048 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [9]), .op(n7475)
         );
  nand2_1 U9049 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [9]), .op(n7474)
         );
  nand2_1 U9050 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [11]), .op(n7473)
         );
  nand2_1 U9051 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [11]), .op(n7472)
         );
  not_ab_or_c_or_d U9052 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [11]), 
        .ip3(n7477), .ip4(n7476), .op(n7481) );
  and2_1 U9053 ( .ip1(n8853), .ip2(\CORTEXM0DS_INST/u_logic/Rddvx4 ), .op(
        n7479) );
  and2_1 U9054 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [11]), .op(n7478)
         );
  not_ab_or_c_or_d U9055 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [11]), .ip2(n8917), 
        .ip3(n7479), .ip4(n7478), .op(n7480) );
  nand3_1 U9056 ( .ip1(n7482), .ip2(n7481), .ip3(n7480), .op(n7483) );
  not_ab_or_c_or_d U9057 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [11]), 
        .ip3(n7484), .ip4(n7483), .op(n11260) );
  nor2_1 U9058 ( .ip1(n11260), .ip2(n8292), .op(n7485) );
  not_ab_or_c_or_d U9059 ( .ip1(n8295), .ip2(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), 
        .ip3(n8294), .ip4(n7485), .op(n7486) );
  mux2_1 U9060 ( .ip1(n8297), .ip2(n8013), .s(n7486), .op(n9145) );
  and2_1 U9061 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [11]), .op(n7498)
         );
  and2_1 U9062 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [11]), .op(n7492)
         );
  nand2_1 U9063 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [9]), .op(n7490)
         );
  nand2_1 U9064 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/Rddvx4 ), .op(
        n7489) );
  nand2_1 U9065 ( .ip1(n8946), .ip2(n9276), .op(n7488) );
  nand2_1 U9066 ( .ip1(\CORTEXM0DS_INST/u_logic/Gcdvx4 ), .ip2(n8948), .op(
        n7487) );
  not_ab_or_c_or_d U9067 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [11]), .ip2(n8966), 
        .ip3(n7492), .ip4(n7491), .op(n7496) );
  nand2_1 U9068 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [11]), .op(n7495)
         );
  nand2_1 U9069 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [11]), .op(n7494)
         );
  nand2_1 U9070 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [9]), .op(n7493)
         );
  nand4_1 U9071 ( .ip1(n7496), .ip2(n7495), .ip3(n7494), .ip4(n7493), .op(
        n7497) );
  not_ab_or_c_or_d U9072 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [11]), .ip2(n8956), 
        .ip3(n7498), .ip4(n7497), .op(n12134) );
  nor2_1 U9073 ( .ip1(n8974), .ip2(n12134), .op(n7719) );
  nand2_1 U9074 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [10]), .ip2(n8914), .op(n7501)
         );
  nand2_1 U9075 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [10]), .op(n7500)
         );
  nand2_1 U9076 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [10]), .op(n7499)
         );
  nand3_1 U9077 ( .ip1(n7501), .ip2(n7500), .ip3(n7499), .op(n7520) );
  and2_1 U9078 ( .ip1(n8853), .ip2(\CORTEXM0DS_INST/u_logic/Gcdvx4 ), .op(
        n7502) );
  or2_1 U9079 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [10]), .ip2(n7502), .op(n7504)
         );
  or2_1 U9080 ( .ip1(n8915), .ip2(n7502), .op(n7503) );
  nand2_1 U9081 ( .ip1(n7504), .ip2(n7503), .op(n7518) );
  nand2_1 U9082 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [10]), .op(n7508)
         );
  nand2_1 U9083 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [10]), .op(n7507)
         );
  nand2_1 U9084 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [10]), .op(n7506)
         );
  nand2_1 U9085 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [10]), .op(n7505)
         );
  nand2_1 U9086 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [8]), .op(n7512)
         );
  nand2_1 U9087 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [10]), .op(n7511)
         );
  nand2_1 U9088 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [10]), .op(n7510)
         );
  nand2_1 U9089 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [10]), .op(n7509)
         );
  not_ab_or_c_or_d U9090 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [8]), 
        .ip3(n7514), .ip4(n7513), .op(n7517) );
  nand2_1 U9091 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [10]), .op(n7516)
         );
  nand2_1 U9092 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [10]), .op(n7515)
         );
  not_ab_or_c_or_d U9093 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [10]), 
        .ip3(n7520), .ip4(n7519), .op(n11255) );
  nor2_1 U9094 ( .ip1(n11255), .ip2(n8292), .op(n7522) );
  inv_1 U9095 ( .ip(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .op(n12580) );
  nor2_1 U9096 ( .ip1(n12580), .ip2(n8008), .op(n7521) );
  not_ab_or_c_or_d U9097 ( .ip1(n7575), .ip2(\CORTEXM0DS_INST/u_logic/Wv9vx4 ), 
        .ip3(n7522), .ip4(n7521), .op(n7523) );
  mux2_1 U9098 ( .ip1(n8297), .ip2(n8013), .s(n7523), .op(n9061) );
  and2_1 U9099 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [10]), .op(n7535)
         );
  and2_1 U9100 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [10]), .op(n7529)
         );
  nand2_1 U9101 ( .ip1(n8946), .ip2(n9275), .op(n7527) );
  nand2_1 U9102 ( .ip1(\CORTEXM0DS_INST/u_logic/Wadvx4 ), .ip2(n8948), .op(
        n7526) );
  nand2_1 U9103 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/Gcdvx4 ), .op(
        n7525) );
  nand2_1 U9104 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [8]), .op(n7524)
         );
  not_ab_or_c_or_d U9105 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [10]), .ip2(n8966), 
        .ip3(n7529), .ip4(n7528), .op(n7533) );
  nand2_1 U9106 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [10]), .op(n7532)
         );
  nand2_1 U9107 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [10]), .op(n7531)
         );
  nand2_1 U9108 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [8]), .op(n7530)
         );
  nand4_1 U9109 ( .ip1(n7533), .ip2(n7532), .ip3(n7531), .ip4(n7530), .op(
        n7534) );
  not_ab_or_c_or_d U9110 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [10]), .ip2(n8945), 
        .ip3(n7535), .ip4(n7534), .op(n12123) );
  nor2_1 U9111 ( .ip1(n8974), .ip2(n12123), .op(n7703) );
  nand2_1 U9112 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n8295), .op(
        n7561) );
  nand2_1 U9113 ( .ip1(\CORTEXM0DS_INST/u_logic/Su9vx4 ), .ip2(n7575), .op(
        n7560) );
  nor2_1 U9114 ( .ip1(n7536), .ip2(n9582), .op(n7651) );
  nand2_1 U9115 ( .ip1(\CORTEXM0DS_INST/u_logic/Ks9vx4 ), .ip2(n7651), .op(
        n7559) );
  nand2_1 U9116 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [9]), .op(n7540)
         );
  nand2_1 U9117 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [9]), .op(n7539)
         );
  nand2_1 U9118 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [9]), .op(n7538)
         );
  nand2_1 U9119 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [9]), .op(n7537)
         );
  nand2_1 U9120 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [7]), .op(n7544)
         );
  nand2_1 U9121 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [7]), .op(n7543)
         );
  nand2_1 U9122 ( .ip1(n8853), .ip2(\CORTEXM0DS_INST/u_logic/Wadvx4 ), .op(
        n7542) );
  nand2_1 U9123 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [9]), .op(n7541)
         );
  not_ab_or_c_or_d U9124 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [9]), 
        .ip3(n7546), .ip4(n7545), .op(n7557) );
  nand2_1 U9125 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [9]), .op(n7549)
         );
  nand2_1 U9126 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [9]), .op(n7548)
         );
  nand2_1 U9127 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [9]), .op(n7547)
         );
  nand3_1 U9128 ( .ip1(n7549), .ip2(n7548), .ip3(n7547), .op(n7555) );
  nand2_1 U9129 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [9]), .op(n7553)
         );
  nand2_1 U9130 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [9]), .op(n7552)
         );
  nand2_1 U9131 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [9]), .op(n7551)
         );
  nand2_1 U9132 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [9]), .op(n7550)
         );
  not_ab_or_c_or_d U9133 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [9]), 
        .ip3(n7555), .ip4(n7554), .op(n7556) );
  nand2_1 U9134 ( .ip1(n7557), .ip2(n7556), .op(n12659) );
  nand2_1 U9135 ( .ip1(n8011), .ip2(n12659), .op(n7558) );
  mux2_1 U9136 ( .ip1(n8013), .ip2(n8297), .s(n7562), .op(n9050) );
  and2_1 U9137 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [9]), .op(n7574)
         );
  and2_1 U9138 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [9]), .op(n7568)
         );
  nand2_1 U9139 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [7]), .op(n7566)
         );
  nand2_1 U9140 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/Wadvx4 ), .op(
        n7565) );
  nand2_1 U9141 ( .ip1(n8946), .ip2(n9284), .op(n7564) );
  nand2_1 U9142 ( .ip1(\CORTEXM0DS_INST/u_logic/M9dvx4 ), .ip2(n8948), .op(
        n7563) );
  not_ab_or_c_or_d U9143 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [9]), .ip2(n8966), 
        .ip3(n7568), .ip4(n7567), .op(n7572) );
  nand2_1 U9144 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [9]), .op(n7571)
         );
  nand2_1 U9145 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [9]), .op(n7570)
         );
  nand2_1 U9146 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [7]), .op(n7569)
         );
  nand4_1 U9147 ( .ip1(n7572), .ip2(n7571), .ip3(n7570), .ip4(n7569), .op(
        n7573) );
  not_ab_or_c_or_d U9148 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [9]), .ip2(n8944), 
        .ip3(n7574), .ip4(n7573), .op(n9055) );
  nor2_1 U9149 ( .ip1(n8974), .ip2(n9055), .op(n7705) );
  nand2_1 U9150 ( .ip1(\CORTEXM0DS_INST/u_logic/R89vx4 ), .ip2(n8295), .op(
        n7599) );
  nand2_1 U9151 ( .ip1(\CORTEXM0DS_INST/u_logic/Ot9vx4 ), .ip2(n7575), .op(
        n7598) );
  nand2_1 U9152 ( .ip1(\CORTEXM0DS_INST/u_logic/Gr9vx4 ), .ip2(n7651), .op(
        n7597) );
  nand2_1 U9153 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [8]), .op(n7579)
         );
  nand2_1 U9154 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [8]), .op(n7578)
         );
  nand2_1 U9155 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [8]), .op(n7577)
         );
  nand2_1 U9156 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [8]), .op(n7576)
         );
  and4_1 U9157 ( .ip1(n7579), .ip2(n7578), .ip3(n7577), .ip4(n7576), .op(n7595) );
  and2_1 U9158 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [8]), .op(n7581)
         );
  inv_1 U9159 ( .ip(\CORTEXM0DS_INST/u_logic/M9dvx4 ), .op(n12118) );
  nor2_1 U9160 ( .ip1(n8909), .ip2(n12118), .op(n7580) );
  not_ab_or_c_or_d U9161 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [8]), .ip2(n8925), 
        .ip3(n7581), .ip4(n7580), .op(n7594) );
  nand2_1 U9162 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [8]), .op(n7585)
         );
  nand2_1 U9163 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [8]), .op(n7584)
         );
  nand2_1 U9164 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [8]), .op(n7583)
         );
  nand2_1 U9165 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [8]), .op(n7582)
         );
  nand2_1 U9166 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [6]), .op(n7589)
         );
  nand2_1 U9167 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [6]), .op(n7588)
         );
  nand2_1 U9168 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [8]), .op(n7587)
         );
  nand2_1 U9169 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [8]), .op(n7586)
         );
  not_ab_or_c_or_d U9170 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [8]), 
        .ip3(n7591), .ip4(n7590), .op(n7593) );
  nand2_1 U9171 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [8]), .op(n7592)
         );
  nand2_1 U9172 ( .ip1(n8011), .ip2(n12658), .op(n7596) );
  mux2_1 U9173 ( .ip1(n8013), .ip2(n8297), .s(n7600), .op(n9136) );
  and2_1 U9174 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [8]), .op(n7612)
         );
  and2_1 U9175 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [8]), .op(n7606)
         );
  nand2_1 U9176 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [6]), .op(n7604)
         );
  nand2_1 U9177 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/M9dvx4 ), .op(
        n7603) );
  nand2_1 U9178 ( .ip1(n8946), .ip2(n9283), .op(n7602) );
  nand2_1 U9179 ( .ip1(\CORTEXM0DS_INST/u_logic/C8dvx4 ), .ip2(n8948), .op(
        n7601) );
  not_ab_or_c_or_d U9180 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [8]), .ip2(n8958), 
        .ip3(n7606), .ip4(n7605), .op(n7610) );
  nand2_1 U9181 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [8]), .op(n7609)
         );
  nand2_1 U9182 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [8]), .op(n7608)
         );
  nand2_1 U9183 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [6]), .op(n7607)
         );
  nand4_1 U9184 ( .ip1(n7610), .ip2(n7609), .ip3(n7608), .ip4(n7607), .op(
        n7611) );
  not_ab_or_c_or_d U9185 ( .ip1(n8966), .ip2(\CORTEXM0DS_INST/cm0_r12 [8]), 
        .ip3(n7612), .ip4(n7611), .op(n12114) );
  nor2_1 U9186 ( .ip1(n8974), .ip2(n12114), .op(n7707) );
  and2_1 U9187 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [7]), .op(n7614)
         );
  and2_1 U9188 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [7]), .op(n7613)
         );
  not_ab_or_c_or_d U9189 ( .ip1(\CORTEXM0DS_INST/vis_msp [5]), .ip2(n8922), 
        .ip3(n7614), .ip4(n7613), .op(n7622) );
  nand2_1 U9190 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [7]), .op(n7617)
         );
  nand2_1 U9191 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [7]), .op(n7616)
         );
  nand2_1 U9192 ( .ip1(n8853), .ip2(\CORTEXM0DS_INST/u_logic/C8dvx4 ), .op(
        n7615) );
  nand3_1 U9193 ( .ip1(n7617), .ip2(n7616), .ip3(n7615), .op(n7618) );
  not_ab_or_c_or_d U9194 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [7]), 
        .ip3(n9499), .ip4(n7618), .op(n7621) );
  nand2_1 U9195 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [5]), .op(n7620)
         );
  nand2_1 U9196 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [7]), .op(n7619)
         );
  nand2_1 U9197 ( .ip1(n8011), .ip2(n12681), .op(n7626) );
  nand2_1 U9198 ( .ip1(\CORTEXM0DS_INST/u_logic/Ks9vx4 ), .ip2(n7670), .op(
        n7625) );
  nand2_1 U9199 ( .ip1(\CORTEXM0DS_INST/u_logic/K79vx4 ), .ip2(n8295), .op(
        n7624) );
  nand2_1 U9200 ( .ip1(\CORTEXM0DS_INST/u_logic/Cq9vx4 ), .ip2(n7651), .op(
        n7623) );
  mux2_1 U9201 ( .ip1(n8013), .ip2(n8297), .s(n7627), .op(n9026) );
  and2_1 U9202 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [7]), .op(n7636)
         );
  nor2_1 U9203 ( .ip1(n7628), .ip2(n8887), .op(n7630) );
  and2_1 U9204 ( .ip1(n8948), .ip2(\CORTEXM0DS_INST/u_logic/S6dvx4 ), .op(
        n7629) );
  not_ab_or_c_or_d U9205 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/C8dvx4 ), 
        .ip3(n7630), .ip4(n7629), .op(n7634) );
  nand2_1 U9206 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [7]), .op(n7633)
         );
  nand2_1 U9207 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [7]), .op(n7632)
         );
  nand2_1 U9208 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [5]), .op(n7631)
         );
  not_ab_or_c_or_d U9209 ( .ip1(n8966), .ip2(\CORTEXM0DS_INST/cm0_r12 [7]), 
        .ip3(n7636), .ip4(n7635), .op(n7640) );
  nand2_1 U9210 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [7]), .op(n7639)
         );
  nand2_1 U9211 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [7]), .op(n7638)
         );
  nand2_1 U9212 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [5]), .op(n7637)
         );
  and4_1 U9213 ( .ip1(n7640), .ip2(n7639), .ip3(n7638), .ip4(n7637), .op(
        n12296) );
  nor2_1 U9214 ( .ip1(n8974), .ip2(n12296), .op(n7709) );
  and2_1 U9215 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [6]), .op(n7642)
         );
  inv_1 U9216 ( .ip(\CORTEXM0DS_INST/cm0_r14 [6]), .op(n7657) );
  nor2_1 U9217 ( .ip1(n8143), .ip2(n7657), .op(n7641) );
  not_ab_or_c_or_d U9218 ( .ip1(\CORTEXM0DS_INST/vis_msp [4]), .ip2(n8922), 
        .ip3(n7642), .ip4(n7641), .op(n7650) );
  nand2_1 U9219 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [6]), .op(n7645)
         );
  nand2_1 U9220 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [6]), .op(n7644)
         );
  nand2_1 U9221 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [6]), .op(n7643)
         );
  nand3_1 U9222 ( .ip1(n7645), .ip2(n7644), .ip3(n7643), .op(n7646) );
  not_ab_or_c_or_d U9223 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [6]), 
        .ip3(n9498), .ip4(n7646), .op(n7649) );
  nand2_1 U9224 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [4]), .op(n7648)
         );
  nand2_1 U9225 ( .ip1(n8853), .ip2(\CORTEXM0DS_INST/u_logic/S6dvx4 ), .op(
        n7647) );
  nand2_1 U9226 ( .ip1(n8011), .ip2(n12677), .op(n7655) );
  nand2_1 U9227 ( .ip1(\CORTEXM0DS_INST/u_logic/Gr9vx4 ), .ip2(n7670), .op(
        n7654) );
  nand2_1 U9228 ( .ip1(\CORTEXM0DS_INST/u_logic/D69vx4 ), .ip2(n8295), .op(
        n7653) );
  nand2_1 U9229 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(n7651), .op(
        n7652) );
  mux2_1 U9230 ( .ip1(n8013), .ip2(n8297), .s(n7656), .op(n11406) );
  nor2_1 U9231 ( .ip1(n8154), .ip2(n7657), .op(n7669) );
  and2_1 U9232 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [6]), .op(n7663)
         );
  nand2_1 U9233 ( .ip1(n8946), .ip2(n9282), .op(n7661) );
  nand2_1 U9234 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/S6dvx4 ), .op(
        n7660) );
  nand2_1 U9235 ( .ip1(\CORTEXM0DS_INST/u_logic/I5dvx4 ), .ip2(n8948), .op(
        n7659) );
  nand2_1 U9236 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [4]), .op(n7658)
         );
  not_ab_or_c_or_d U9237 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [6]), 
        .ip3(n7663), .ip4(n7662), .op(n7667) );
  nand2_1 U9238 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [6]), .op(n7666)
         );
  nand2_1 U9239 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [6]), .op(n7665)
         );
  nand2_1 U9240 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [4]), .op(n7664)
         );
  nand4_1 U9241 ( .ip1(n7667), .ip2(n7666), .ip3(n7665), .ip4(n7664), .op(
        n7668) );
  not_ab_or_c_or_d U9242 ( .ip1(n8966), .ip2(\CORTEXM0DS_INST/cm0_r12 [6]), 
        .ip3(n7669), .ip4(n7668), .op(n12240) );
  nor2_1 U9243 ( .ip1(n8974), .ip2(n12240), .op(n7711) );
  nand2_1 U9244 ( .ip1(\CORTEXM0DS_INST/u_logic/Cq9vx4 ), .ip2(n7670), .op(
        n7686) );
  nand2_1 U9245 ( .ip1(\CORTEXM0DS_INST/u_logic/W49vx4 ), .ip2(n8295), .op(
        n7685) );
  inv_1 U9246 ( .ip(\CORTEXM0DS_INST/u_logic/I5dvx4 ), .op(n12234) );
  nor2_1 U9247 ( .ip1(n8909), .ip2(n12234), .op(n7672) );
  and2_1 U9248 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [3]), .op(n7671)
         );
  not_ab_or_c_or_d U9249 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [5]), 
        .ip3(n7672), .ip4(n7671), .op(n7681) );
  nand2_1 U9250 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [5]), .ip2(n8910), .op(n7675)
         );
  nand2_1 U9251 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [5]), .op(n7674)
         );
  nand2_1 U9252 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [5]), .op(n7673)
         );
  nand3_1 U9253 ( .ip1(n7675), .ip2(n7674), .ip3(n7673), .op(n7676) );
  not_ab_or_c_or_d U9254 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [5]), 
        .ip3(n7677), .ip4(n7676), .op(n7680) );
  nand2_1 U9255 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [3]), .op(n7679)
         );
  nand2_1 U9256 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [5]), .op(n7678)
         );
  nand2_1 U9257 ( .ip1(n8011), .ip2(n12675), .op(n7684) );
  nand2_1 U9258 ( .ip1(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .ip2(n7682), .op(
        n7683) );
  mux2_1 U9259 ( .ip1(n8013), .ip2(n8297), .s(n7687), .op(n9080) );
  and2_1 U9260 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [5]), .op(n7695)
         );
  nor2_1 U9261 ( .ip1(n7975), .ip2(n12234), .op(n7689) );
  nor2_1 U9262 ( .ip1(n9258), .ip2(n8887), .op(n7688) );
  not_ab_or_c_or_d U9263 ( .ip1(\CORTEXM0DS_INST/u_logic/Y3dvx4 ), .ip2(n8948), 
        .ip3(n7689), .ip4(n7688), .op(n7693) );
  nand2_1 U9264 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [5]), .op(n7692)
         );
  nand2_1 U9265 ( .ip1(n8966), .ip2(\CORTEXM0DS_INST/cm0_r12 [5]), .op(n7691)
         );
  nand2_1 U9266 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [3]), .op(n7690)
         );
  not_ab_or_c_or_d U9267 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [5]), .ip2(n8956), 
        .ip3(n7695), .ip4(n7694), .op(n7699) );
  nand2_1 U9268 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [5]), .op(n7698)
         );
  nand2_1 U9269 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [5]), .op(n7697)
         );
  nand2_1 U9270 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [3]), .op(n7696)
         );
  and2_1 U9271 ( .ip1(n8969), .ip2(n12233), .op(n7714) );
  fulladder U9272 ( .a(n9169), .b(n7701), .ci(n7700), .co(n7713), .s(n7716) );
  fulladder U9273 ( .a(n9061), .b(n7703), .ci(n7702), .co(n7718), .s(n9020) );
  fulladder U9274 ( .a(n9050), .b(n7705), .ci(n7704), .co(n7702), .s(n8528) );
  inv_1 U9275 ( .ip(n8528), .op(n7717) );
  fulladder U9276 ( .a(n9136), .b(n7707), .ci(n7706), .co(n7704), .s(n9220) );
  fulladder U9277 ( .a(n9026), .b(n7709), .ci(n7708), .co(n7706), .s(n9030) );
  fulladder U9278 ( .a(n11406), .b(n7711), .ci(n7710), .co(n7708), .s(n7712)
         );
  inv_1 U9279 ( .ip(n7712), .op(n9214) );
  fulladder U9280 ( .a(n9080), .b(n7714), .ci(n7713), .co(n7710), .s(n9216) );
  and2_1 U9281 ( .ip1(n7716), .ip2(n7715), .op(n9215) );
  nand2_1 U9282 ( .ip1(n9216), .ip2(n9215), .op(n9213) );
  nor2_1 U9283 ( .ip1(n9214), .ip2(n9213), .op(n9029) );
  and2_1 U9284 ( .ip1(n9030), .ip2(n9029), .op(n9219) );
  nand2_1 U9285 ( .ip1(n9220), .ip2(n9219), .op(n8527) );
  nor2_1 U9286 ( .ip1(n7717), .ip2(n8527), .op(n9019) );
  nand2_1 U9287 ( .ip1(n9020), .ip2(n9019), .op(n9217) );
  fulladder U9288 ( .a(n9145), .b(n7719), .ci(n7718), .co(n7721), .s(n7720) );
  inv_1 U9289 ( .ip(n7720), .op(n9218) );
  nor2_1 U9290 ( .ip1(n9217), .ip2(n9218), .op(n9221) );
  fulladder U9291 ( .a(n9143), .b(n7722), .ci(n7721), .co(n8311), .s(n9222) );
  nand2_1 U9292 ( .ip1(n9221), .ip2(n9222), .op(n8383) );
  xor2_1 U9293 ( .ip1(n8382), .ip2(n8383), .op(n9229) );
  inv_1 U9294 ( .ip(n9229), .op(n11292) );
  nand2_1 U9295 ( .ip1(n11292), .ip2(n10572), .op(n7809) );
  nor2_1 U9296 ( .ip1(n7723), .ip2(n10490), .op(n7724) );
  not_ab_or_c_or_d U9297 ( .ip1(\CORTEXM0DS_INST/u_logic/Zph2z4 [1]), .ip2(
        n11212), .ip3(n7724), .ip4(n9933), .op(n7726) );
  or2_1 U9298 ( .ip1(n7726), .ip2(n7725), .op(n10323) );
  inv_1 U9299 ( .ip(n11614), .op(n10184) );
  nand2_1 U9300 ( .ip1(n9429), .ip2(n9368), .op(n7730) );
  nand2_1 U9301 ( .ip1(n9431), .ip2(n9434), .op(n7729) );
  nand2_1 U9302 ( .ip1(n9433), .ip2(n9369), .op(n7728) );
  nand2_1 U9303 ( .ip1(n9435), .ip2(n9367), .op(n7727) );
  nand4_1 U9304 ( .ip1(n7730), .ip2(n7729), .ip3(n7728), .ip4(n7727), .op(
        n9998) );
  nand2_1 U9305 ( .ip1(n10184), .ip2(n9998), .op(n7751) );
  and2_1 U9306 ( .ip1(n9890), .ip2(n9895), .op(n7732) );
  nor2_1 U9307 ( .ip1(n7731), .ip2(n9895), .op(n9901) );
  nor2_1 U9308 ( .ip1(n7732), .ip2(n9901), .op(n7737) );
  nor2_1 U9309 ( .ip1(n7734), .ip2(n7733), .op(n9886) );
  nor2_1 U9310 ( .ip1(n7735), .ip2(n9886), .op(n7736) );
  mux2_1 U9311 ( .ip1(n7737), .ip2(n7736), .s(n10140), .op(n7738) );
  nand2_1 U9312 ( .ip1(n9903), .ip2(n7738), .op(n7739) );
  not_ab_or_c_or_d U9313 ( .ip1(n9879), .ip2(n7739), .ip3(
        \CORTEXM0DS_INST/u_logic/Krgvx4 ), .ip4(
        \CORTEXM0DS_INST/u_logic/Eqgvx4 ), .op(n12464) );
  inv_1 U9314 ( .ip(n10152), .op(n10266) );
  nor2_1 U9315 ( .ip1(n12464), .ip2(n10266), .op(n7744) );
  nand2_1 U9316 ( .ip1(n11610), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [13]), 
        .op(n7742) );
  nand2_1 U9317 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [13]), .ip2(n11787), 
        .op(n7741) );
  nand2_1 U9318 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [13]), .ip2(n10265), 
        .op(n7740) );
  nand4_1 U9319 ( .ip1(n2976), .ip2(n7742), .ip3(n7741), .ip4(n7740), .op(
        n7743) );
  not_ab_or_c_or_d U9320 ( .ip1(n11609), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [13]), .ip3(n7744), .ip4(n7743), .op(
        n7750) );
  inv_1 U9321 ( .ip(n9419), .op(n9430) );
  nand2_1 U9322 ( .ip1(n9429), .ip2(n9430), .op(n7748) );
  nand2_1 U9323 ( .ip1(n9433), .ip2(n9428), .op(n7747) );
  nand2_1 U9324 ( .ip1(n9431), .ip2(n9270), .op(n7746) );
  nand2_1 U9325 ( .ip1(n9435), .ip2(n9432), .op(n7745) );
  nand4_1 U9326 ( .ip1(n7748), .ip2(n7747), .ip3(n7746), .ip4(n7745), .op(
        n9978) );
  nand2_1 U9327 ( .ip1(n11607), .ip2(n9978), .op(n7749) );
  nand3_1 U9328 ( .ip1(n7751), .ip2(n7750), .ip3(n7749), .op(n10362) );
  nand2_1 U9329 ( .ip1(n10323), .ip2(n10362), .op(n7807) );
  inv_1 U9330 ( .ip(n9312), .op(n9346) );
  nand2_1 U9331 ( .ip1(n9325), .ip2(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .op(
        n9347) );
  mux2_1 U9332 ( .ip1(n9346), .ip2(n9347), .s(n9435), .op(n7752) );
  inv_1 U9333 ( .ip(n7752), .op(n7762) );
  nand2_1 U9334 ( .ip1(n10109), .ip2(n7762), .op(n7764) );
  nor2_1 U9335 ( .ip1(n9293), .ip2(n9416), .op(n7756) );
  nor2_1 U9336 ( .ip1(n9296), .ip2(n9418), .op(n7755) );
  nor2_1 U9337 ( .ip1(n9295), .ip2(n9420), .op(n7754) );
  nor2_1 U9338 ( .ip1(n9257), .ip2(n9392), .op(n7753) );
  nor4_1 U9339 ( .ip1(n7756), .ip2(n7755), .ip3(n7754), .ip4(n7753), .op(n9987) );
  nand2_1 U9340 ( .ip1(n9429), .ip2(n9330), .op(n7760) );
  nand2_1 U9341 ( .ip1(n9433), .ip2(n9329), .op(n7759) );
  nand2_1 U9342 ( .ip1(n9431), .ip2(n9304), .op(n7758) );
  nand2_1 U9343 ( .ip1(n9435), .ip2(n9331), .op(n7757) );
  nand4_1 U9344 ( .ip1(n7760), .ip2(n7759), .ip3(n7758), .ip4(n7757), .op(
        n9311) );
  nor2_1 U9345 ( .ip1(n9311), .ip2(n9443), .op(n7761) );
  not_ab_or_c_or_d U9346 ( .ip1(n9987), .ip2(n9443), .ip3(n7762), .ip4(n7761), 
        .op(n9315) );
  nand2_1 U9347 ( .ip1(n9315), .ip2(n11821), .op(n7763) );
  nand4_1 U9348 ( .ip1(n3067), .ip2(n10267), .ip3(n7764), .ip4(n7763), .op(
        n10360) );
  nand2_1 U9349 ( .ip1(n7766), .ip2(n7765), .op(n7768) );
  nand2_1 U9350 ( .ip1(n7768), .ip2(n7767), .op(n7769) );
  nand2_1 U9351 ( .ip1(n7769), .ip2(n9873), .op(n10322) );
  nor2_1 U9352 ( .ip1(n9350), .ip2(n9420), .op(n7773) );
  nor2_1 U9353 ( .ip1(n9319), .ip2(n9418), .op(n7772) );
  nor2_1 U9354 ( .ip1(n9318), .ip2(n9416), .op(n7771) );
  nor2_1 U9355 ( .ip1(n9317), .ip2(n9392), .op(n7770) );
  nor4_1 U9356 ( .ip1(n7773), .ip2(n7772), .ip3(n7771), .ip4(n7770), .op(n9383) );
  nor2_1 U9357 ( .ip1(n9383), .ip2(n11614), .op(n7782) );
  inv_1 U9358 ( .ip(n8014), .op(n9401) );
  nand2_1 U9359 ( .ip1(n9429), .ip2(n9401), .op(n7778) );
  nand2_1 U9360 ( .ip1(n9433), .ip2(n9403), .op(n7777) );
  inv_1 U9361 ( .ip(n7774), .op(n9370) );
  nand2_1 U9362 ( .ip1(n9431), .ip2(n9370), .op(n7776) );
  nand2_1 U9363 ( .ip1(n9435), .ip2(n9402), .op(n7775) );
  nand4_1 U9364 ( .ip1(n7778), .ip2(n7777), .ip3(n7776), .ip4(n7775), .op(
        n9999) );
  nand2_1 U9365 ( .ip1(n11607), .ip2(n9999), .op(n7780) );
  nand2_1 U9366 ( .ip1(n11609), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [21]), 
        .op(n7779) );
  nand3_1 U9367 ( .ip1(n7780), .ip2(n3101), .ip3(n7779), .op(n7781) );
  not_ab_or_c_or_d U9368 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [21]), .ip2(
        n11610), .ip3(n7782), .ip4(n7781), .op(n10357) );
  and2_1 U9369 ( .ip1(n9386), .ip2(n10053), .op(n7783) );
  nor2_1 U9370 ( .ip1(n10054), .ip2(n7783), .op(n10310) );
  nor2_1 U9371 ( .ip1(n10357), .ip2(n10310), .op(n7798) );
  nand2_1 U9372 ( .ip1(n9429), .ip2(n9275), .op(n7787) );
  nand2_1 U9373 ( .ip1(n9431), .ip2(n9284), .op(n7786) );
  nand2_1 U9374 ( .ip1(n9433), .ip2(n9276), .op(n7785) );
  nand2_1 U9375 ( .ip1(n9435), .ip2(n9269), .op(n7784) );
  nand4_1 U9376 ( .ip1(n7787), .ip2(n7786), .ip3(n7785), .ip4(n7784), .op(
        n9982) );
  inv_1 U9377 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [5]), .op(n11643) );
  nor2_1 U9378 ( .ip1(n11643), .ip2(n11841), .op(n7795) );
  nand2_1 U9379 ( .ip1(n9429), .ip2(n9282), .op(n7791) );
  nand2_1 U9380 ( .ip1(n9431), .ip2(n9263), .op(n7790) );
  nand2_1 U9381 ( .ip1(n9433), .ip2(n9281), .op(n7789) );
  nand2_1 U9382 ( .ip1(n9435), .ip2(n9283), .op(n7788) );
  nand4_1 U9383 ( .ip1(n7791), .ip2(n7790), .ip3(n7789), .ip4(n7788), .op(
        n9994) );
  nand2_1 U9384 ( .ip1(n11607), .ip2(n9994), .op(n7793) );
  nand2_1 U9385 ( .ip1(n11610), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [5]), 
        .op(n7792) );
  nand3_1 U9386 ( .ip1(n7793), .ip2(n3084), .ip3(n7792), .op(n7794) );
  not_ab_or_c_or_d U9387 ( .ip1(n10184), .ip2(n9982), .ip3(n7795), .ip4(n7794), 
        .op(n10356) );
  inv_1 U9388 ( .ip(n10055), .op(n9874) );
  nor3_1 U9389 ( .ip1(n9469), .ip2(n10047), .ip3(n9874), .op(n10052) );
  nor2_1 U9390 ( .ip1(n10052), .ip2(n7796), .op(n10296) );
  nor2_1 U9391 ( .ip1(n10356), .ip2(n10296), .op(n7797) );
  not_ab_or_c_or_d U9392 ( .ip1(n10360), .ip2(n10322), .ip3(n7798), .ip4(n7797), .op(n7806) );
  not_ab_or_c_or_d U9393 ( .ip1(n9874), .ip2(n7800), .ip3(n7799), .ip4(n9361), 
        .op(n9387) );
  nor2_1 U9394 ( .ip1(n7801), .ip2(n9387), .op(n9451) );
  inv_1 U9395 ( .ip(n9451), .op(n7805) );
  nor2_1 U9396 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(n10975) );
  nor2_1 U9397 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n11038), .op(
        n8614) );
  nor2_1 U9398 ( .ip1(n6210), .ip2(n10587), .op(n7803) );
  inv_1 U9399 ( .ip(n7802), .op(n9867) );
  not_ab_or_c_or_d U9400 ( .ip1(n10975), .ip2(n8614), .ip3(n7803), .ip4(n9867), 
        .op(n7804) );
  not_ab_or_c_or_d U9401 ( .ip1(n7805), .ip2(n9933), .ip3(n7804), .ip4(n9871), 
        .op(n10330) );
  inv_1 U9402 ( .ip(n10330), .op(n10314) );
  nand3_1 U9403 ( .ip1(n7807), .ip2(n7806), .ip3(n10314), .op(n11290) );
  nand2_1 U9404 ( .ip1(n10859), .ip2(n11290), .op(n7808) );
  nand4_1 U9405 ( .ip1(n7810), .ip2(n10573), .ip3(n7809), .ip4(n7808), .op(
        \CORTEXM0DS_INST/u_logic/Nehvx4 ) );
  nand2_1 U9406 ( .ip1(\CORTEXM0DS_INST/u_logic/W1evx4 ), .ip2(n2120), .op(
        n8401) );
  nand2_1 U9407 ( .ip1(\CORTEXM0DS_INST/vis_pc [27]), .ip2(n12321), .op(n8400)
         );
  nand2_1 U9408 ( .ip1(\CORTEXM0DS_INST/vis_apsr [0]), .ip2(n12320), .op(n8399) );
  inv_1 U9409 ( .ip(n12691), .op(n12317) );
  and2_1 U9410 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [27]), .op(n7818)
         );
  nor2_1 U9411 ( .ip1(n9319), .ip2(n8887), .op(n7812) );
  inv_1 U9412 ( .ip(\CORTEXM0DS_INST/u_logic/Azdvx4 ), .op(n12263) );
  nor2_1 U9413 ( .ip1(n12051), .ip2(n12263), .op(n7811) );
  not_ab_or_c_or_d U9414 ( .ip1(\CORTEXM0DS_INST/u_logic/L0evx4 ), .ip2(n8947), 
        .ip3(n7812), .ip4(n7811), .op(n7816) );
  nand2_1 U9415 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [27]), .op(n7815)
         );
  nand2_1 U9416 ( .ip1(n8966), .ip2(\CORTEXM0DS_INST/cm0_r12 [27]), .op(n7814)
         );
  nand2_1 U9417 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [25]), .op(n7813)
         );
  not_ab_or_c_or_d U9418 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [27]), 
        .ip3(n7818), .ip4(n7817), .op(n7822) );
  nand2_1 U9419 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [27]), .op(n7821)
         );
  nand2_1 U9420 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [27]), .op(n7820)
         );
  nand2_1 U9421 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [25]), .op(n7819)
         );
  or2_1 U9422 ( .ip1(n7823), .ip2(n12376), .op(n7825) );
  or2_1 U9423 ( .ip1(n8008), .ip2(n12376), .op(n7824) );
  nand2_1 U9424 ( .ip1(n7825), .ip2(n7824), .op(n7826) );
  mux2_1 U9425 ( .ip1(n8297), .ip2(n8013), .s(n7826), .op(n8942) );
  mux2_1 U9426 ( .ip1(n7827), .ip2(n8942), .s(n8292), .op(n8943) );
  inv_1 U9427 ( .ip(n8943), .op(n8342) );
  inv_1 U9428 ( .ip(n8942), .op(n8341) );
  nand2_1 U9429 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [27]), .op(n7830)
         );
  nand2_1 U9430 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [27]), .op(n7829)
         );
  nand2_1 U9431 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [27]), .op(n7828)
         );
  nand3_1 U9432 ( .ip1(n7830), .ip2(n7829), .ip3(n7828), .op(n7849) );
  inv_1 U9433 ( .ip(\CORTEXM0DS_INST/u_logic/L0evx4 ), .op(n12275) );
  nor2_1 U9434 ( .ip1(n8909), .ip2(n12275), .op(n7831) );
  or2_1 U9435 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [27]), .ip2(n7831), .op(n7833)
         );
  or2_1 U9436 ( .ip1(n8941), .ip2(n7831), .op(n7832) );
  nand2_1 U9437 ( .ip1(n7833), .ip2(n7832), .op(n7847) );
  nand2_1 U9438 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [27]), .op(n7837)
         );
  nand2_1 U9439 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [27]), .op(n7836)
         );
  nand2_1 U9440 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [27]), .op(n7835)
         );
  nand2_1 U9441 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [27]), .op(n7834)
         );
  nand2_1 U9442 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [25]), .op(n7841)
         );
  nand2_1 U9443 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [27]), .op(n7840)
         );
  nand2_1 U9444 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [27]), .op(n7839)
         );
  nand2_1 U9445 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [27]), .op(n7838)
         );
  not_ab_or_c_or_d U9446 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [25]), 
        .ip3(n7843), .ip4(n7842), .op(n7846) );
  nand2_1 U9447 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [27]), .op(n7845)
         );
  nand2_1 U9448 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [27]), .op(n7844)
         );
  not_ab_or_c_or_d U9449 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [27]), 
        .ip3(n7849), .ip4(n7848), .op(n9853) );
  mux2_1 U9450 ( .ip1(n8342), .ip2(n8341), .s(n9853), .op(n9193) );
  or2_1 U9451 ( .ip1(n12274), .ip2(n9193), .op(n7850) );
  nand2_1 U9452 ( .ip1(n8969), .ip2(n7850), .op(n8318) );
  nand2_1 U9453 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [26]), .ip2(n8916), .op(n7853)
         );
  nand2_1 U9454 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [26]), .op(n7852)
         );
  nand2_1 U9455 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [26]), .op(n7851)
         );
  nand3_1 U9456 ( .ip1(n7853), .ip2(n7852), .ip3(n7851), .op(n7870) );
  and2_1 U9457 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [24]), .op(n7855)
         );
  and2_1 U9458 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [26]), .op(n7854)
         );
  not_ab_or_c_or_d U9459 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [26]), .ip2(n8917), 
        .ip3(n7855), .ip4(n7854), .op(n7868) );
  nand2_1 U9460 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [26]), .op(n7858)
         );
  nand2_1 U9461 ( .ip1(n8853), .ip2(\CORTEXM0DS_INST/u_logic/Azdvx4 ), .op(
        n7857) );
  nand2_1 U9462 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [26]), .op(n7856)
         );
  nand3_1 U9463 ( .ip1(n7858), .ip2(n7857), .ip3(n7856), .op(n7864) );
  nand2_1 U9464 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [26]), .op(n7862)
         );
  nand2_1 U9465 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [26]), .op(n7861)
         );
  nand2_1 U9466 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [26]), .op(n7860)
         );
  nand2_1 U9467 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [26]), .op(n7859)
         );
  not_ab_or_c_or_d U9468 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [26]), 
        .ip3(n7864), .ip4(n7863), .op(n7867) );
  nand2_1 U9469 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [24]), .op(n7866)
         );
  nand2_1 U9470 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [26]), .op(n7865)
         );
  not_ab_or_c_or_d U9471 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [26]), 
        .ip3(n7870), .ip4(n7869), .op(n9850) );
  mux2_1 U9472 ( .ip1(n8943), .ip2(n8942), .s(n9850), .op(n11427) );
  and2_1 U9473 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [26]), .op(n7882)
         );
  and2_1 U9474 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [26]), .op(n7876)
         );
  nand2_1 U9475 ( .ip1(n8946), .ip2(n9377), .op(n7874) );
  nand2_1 U9476 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [24]), .op(n7873)
         );
  nand2_1 U9477 ( .ip1(\CORTEXM0DS_INST/u_logic/Pxdvx4 ), .ip2(n8948), .op(
        n7872) );
  nand2_1 U9478 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/Azdvx4 ), .op(
        n7871) );
  not_ab_or_c_or_d U9479 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [26]), .ip2(n8966), 
        .ip3(n7876), .ip4(n7875), .op(n7880) );
  nand2_1 U9480 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [26]), .op(n7879)
         );
  nand2_1 U9481 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [26]), .op(n7878)
         );
  nand2_1 U9482 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [24]), .op(n7877)
         );
  nand4_1 U9483 ( .ip1(n7880), .ip2(n7879), .ip3(n7878), .ip4(n7877), .op(
        n7881) );
  not_ab_or_c_or_d U9484 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [26]), .ip2(n8957), 
        .ip3(n7882), .ip4(n7881), .op(n12259) );
  nor2_1 U9485 ( .ip1(n11427), .ip2(n12259), .op(n11435) );
  nand2_1 U9486 ( .ip1(n11435), .ip2(n8969), .op(n8315) );
  nand2_1 U9487 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [25]), .op(n7885)
         );
  nand2_1 U9488 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [25]), .op(n7884)
         );
  nand2_1 U9489 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [25]), .op(n7883)
         );
  nand3_1 U9490 ( .ip1(n7885), .ip2(n7884), .ip3(n7883), .op(n7904) );
  inv_1 U9491 ( .ip(\CORTEXM0DS_INST/u_logic/Pxdvx4 ), .op(n12254) );
  nor2_1 U9492 ( .ip1(n8909), .ip2(n12254), .op(n7886) );
  or2_1 U9493 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [25]), .ip2(n7886), .op(n7888)
         );
  or2_1 U9494 ( .ip1(n8915), .ip2(n7886), .op(n7887) );
  nand2_1 U9495 ( .ip1(n7888), .ip2(n7887), .op(n7902) );
  nand2_1 U9496 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [25]), .op(n7892)
         );
  nand2_1 U9497 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [25]), .op(n7891)
         );
  nand2_1 U9498 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [25]), .op(n7890)
         );
  nand2_1 U9499 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [25]), .op(n7889)
         );
  nand2_1 U9500 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [23]), .op(n7896)
         );
  nand2_1 U9501 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [23]), .op(n7895)
         );
  nand2_1 U9502 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [25]), .op(n7894)
         );
  nand2_1 U9503 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [25]), .op(n7893)
         );
  not_ab_or_c_or_d U9504 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [25]), 
        .ip3(n7898), .ip4(n7897), .op(n7901) );
  nand2_1 U9505 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [25]), .op(n7900)
         );
  nand2_1 U9506 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [25]), .op(n7899)
         );
  ab_or_c_or_d U9507 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [25]), .ip3(
        n7904), .ip4(n7903), .op(n11423) );
  mux2_1 U9508 ( .ip1(n8341), .ip2(n8342), .s(n11423), .op(n9100) );
  and2_1 U9509 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [25]), .op(n7912)
         );
  inv_1 U9510 ( .ip(\CORTEXM0DS_INST/u_logic/Ewdvx4 ), .op(n12316) );
  nor2_1 U9511 ( .ip1(n12051), .ip2(n12316), .op(n7906) );
  nor2_1 U9512 ( .ip1(n9350), .ip2(n8887), .op(n7905) );
  not_ab_or_c_or_d U9513 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [23]), 
        .ip3(n7906), .ip4(n7905), .op(n7910) );
  nand2_1 U9514 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [25]), .op(n7909)
         );
  nand2_1 U9515 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [25]), .op(n7908)
         );
  nand2_1 U9516 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/Pxdvx4 ), .op(
        n7907) );
  not_ab_or_c_or_d U9517 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [25]), 
        .ip3(n7912), .ip4(n7911), .op(n7916) );
  nand2_1 U9518 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [25]), .op(n7915)
         );
  nand2_1 U9519 ( .ip1(n8966), .ip2(\CORTEXM0DS_INST/cm0_r12 [25]), .op(n7914)
         );
  nand2_1 U9520 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [23]), .op(n7913)
         );
  inv_1 U9521 ( .ip(n12253), .op(n9099) );
  nor2_1 U9522 ( .ip1(n8974), .ip2(n9099), .op(n8359) );
  nand2_1 U9523 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [24]), .op(n7919)
         );
  nand2_1 U9524 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [24]), .op(n7918)
         );
  nand2_1 U9525 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [24]), .op(n7917)
         );
  nand3_1 U9526 ( .ip1(n7919), .ip2(n7918), .ip3(n7917), .op(n7938) );
  nor2_1 U9527 ( .ip1(n8909), .ip2(n12316), .op(n7920) );
  or2_1 U9528 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [24]), .ip2(n7920), .op(n7922)
         );
  or2_1 U9529 ( .ip1(n8924), .ip2(n7920), .op(n7921) );
  nand2_1 U9530 ( .ip1(n7922), .ip2(n7921), .op(n7936) );
  nand2_1 U9531 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [24]), .op(n7926)
         );
  nand2_1 U9532 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [24]), .op(n7925)
         );
  nand2_1 U9533 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [24]), .op(n7924)
         );
  nand2_1 U9534 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [24]), .op(n7923)
         );
  nand2_1 U9535 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [22]), .op(n7930)
         );
  nand2_1 U9536 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [22]), .op(n7929)
         );
  nand2_1 U9537 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [24]), .op(n7928)
         );
  nand2_1 U9538 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [24]), .op(n7927)
         );
  not_ab_or_c_or_d U9539 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [24]), 
        .ip3(n7932), .ip4(n7931), .op(n7935) );
  nand2_1 U9540 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [24]), .op(n7934)
         );
  nand2_1 U9541 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [24]), .op(n7933)
         );
  ab_or_c_or_d U9542 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [24]), .ip3(
        n7938), .ip4(n7937), .op(n11413) );
  mux2_1 U9543 ( .ip1(n8341), .ip2(n8342), .s(n11413), .op(n9047) );
  and2_1 U9544 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [24]), .op(n7950)
         );
  and2_1 U9545 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [24]), .op(n7944)
         );
  nand2_1 U9546 ( .ip1(n8946), .ip2(n9402), .op(n7942) );
  nand2_1 U9547 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/Ewdvx4 ), .op(
        n7941) );
  nand2_1 U9548 ( .ip1(\CORTEXM0DS_INST/u_logic/Tudvx4 ), .ip2(n8948), .op(
        n7940) );
  nand2_1 U9549 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [22]), .op(n7939)
         );
  not_ab_or_c_or_d U9550 ( .ip1(n8966), .ip2(\CORTEXM0DS_INST/cm0_r12 [24]), 
        .ip3(n7944), .ip4(n7943), .op(n7948) );
  nand2_1 U9551 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [24]), .op(n7947)
         );
  nand2_1 U9552 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [24]), .op(n7946)
         );
  nand2_1 U9553 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [22]), .op(n7945)
         );
  nand4_1 U9554 ( .ip1(n7948), .ip2(n7947), .ip3(n7946), .ip4(n7945), .op(
        n7949) );
  not_ab_or_c_or_d U9555 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [24]), .ip2(n8957), 
        .ip3(n7950), .ip4(n7949), .op(n9046) );
  nor2_1 U9556 ( .ip1(n8974), .ip2(n9046), .op(n8361) );
  inv_1 U9557 ( .ip(\CORTEXM0DS_INST/cm0_r14 [23]), .op(n7974) );
  nor2_1 U9558 ( .ip1(n8143), .ip2(n7974), .op(n7952) );
  inv_1 U9559 ( .ip(\CORTEXM0DS_INST/u_logic/Tudvx4 ), .op(n12107) );
  nor2_1 U9560 ( .ip1(n8909), .ip2(n12107), .op(n7951) );
  not_ab_or_c_or_d U9561 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [23]), 
        .ip3(n7952), .ip4(n7951), .op(n7970) );
  nand2_1 U9562 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [23]), .op(n7956)
         );
  nand2_1 U9563 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [23]), .op(n7955)
         );
  nand2_1 U9564 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [23]), .op(n7954)
         );
  nand2_1 U9565 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [23]), .op(n7953)
         );
  and4_1 U9566 ( .ip1(n7956), .ip2(n7955), .ip3(n7954), .ip4(n7953), .op(n7969) );
  nand2_1 U9567 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [23]), .op(n7960)
         );
  nand2_1 U9568 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [23]), .op(n7959)
         );
  nand2_1 U9569 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [23]), .op(n7958)
         );
  nand2_1 U9570 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [23]), .op(n7957)
         );
  nand2_1 U9571 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [21]), .op(n7964)
         );
  nand2_1 U9572 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [21]), .op(n7963)
         );
  nand2_1 U9573 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [23]), .op(n7962)
         );
  nand2_1 U9574 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [23]), .op(n7961)
         );
  not_ab_or_c_or_d U9575 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [23]), 
        .ip3(n7966), .ip4(n7965), .op(n7968) );
  nand2_1 U9576 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [23]), .op(n7967)
         );
  nor2_1 U9577 ( .ip1(n12376), .ip2(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .op(
        n7971) );
  not_ab_or_c_or_d U9578 ( .ip1(n12376), .ip2(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip3(n7971), .ip4(n8008), .op(n7972) );
  not_ab_or_c_or_d U9579 ( .ip1(n8011), .ip2(n12678), .ip3(n8294), .ip4(n7972), 
        .op(n7973) );
  mux2_1 U9580 ( .ip1(n8297), .ip2(n8013), .s(n7973), .op(n9056) );
  nor2_1 U9581 ( .ip1(n8154), .ip2(n7974), .op(n7987) );
  inv_1 U9582 ( .ip(\CORTEXM0DS_INST/u_logic/Itdvx4 ), .op(n12223) );
  nor2_1 U9583 ( .ip1(n12051), .ip2(n12223), .op(n7977) );
  nor2_1 U9584 ( .ip1(n7975), .ip2(n12107), .op(n7976) );
  not_ab_or_c_or_d U9585 ( .ip1(n8946), .ip2(n9403), .ip3(n7977), .ip4(n7976), 
        .op(n7981) );
  nand2_1 U9586 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [23]), .op(n7980)
         );
  nand2_1 U9587 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [23]), .op(n7979)
         );
  nand2_1 U9588 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [21]), .op(n7978)
         );
  and4_1 U9589 ( .ip1(n7981), .ip2(n7980), .ip3(n7979), .ip4(n7978), .op(n7985) );
  nand2_1 U9590 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [23]), .op(n7984)
         );
  nand2_1 U9591 ( .ip1(n8966), .ip2(\CORTEXM0DS_INST/cm0_r12 [23]), .op(n7983)
         );
  nand2_1 U9592 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [21]), .op(n7982)
         );
  nand4_1 U9593 ( .ip1(n7985), .ip2(n7984), .ip3(n7983), .ip4(n7982), .op(
        n7986) );
  not_ab_or_c_or_d U9594 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [23]), .ip2(n8956), 
        .ip3(n7987), .ip4(n7986), .op(n12099) );
  nor2_1 U9595 ( .ip1(n8974), .ip2(n12099), .op(n8363) );
  nand2_1 U9596 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [22]), .op(n7991)
         );
  nand2_1 U9597 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [22]), .op(n7990)
         );
  nand2_1 U9598 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [22]), .op(n7989)
         );
  nand2_1 U9599 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [22]), .op(n7988)
         );
  and4_1 U9600 ( .ip1(n7991), .ip2(n7990), .ip3(n7989), .ip4(n7988), .op(n8007) );
  and2_1 U9601 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [22]), .op(n7993)
         );
  nor2_1 U9602 ( .ip1(n8909), .ip2(n12223), .op(n7992) );
  not_ab_or_c_or_d U9603 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [22]), .ip2(n8941), 
        .ip3(n7993), .ip4(n7992), .op(n8006) );
  nand2_1 U9604 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [22]), .op(n7997)
         );
  nand2_1 U9605 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [22]), .op(n7996)
         );
  nand2_1 U9606 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [22]), .op(n7995)
         );
  nand2_1 U9607 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [22]), .op(n7994)
         );
  nand2_1 U9608 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [20]), .op(n8001)
         );
  nand2_1 U9609 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [20]), .op(n8000)
         );
  nand2_1 U9610 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [22]), .op(n7999)
         );
  nand2_1 U9611 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [22]), .op(n7998)
         );
  not_ab_or_c_or_d U9612 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [22]), 
        .ip3(n8003), .ip4(n8002), .op(n8005) );
  nand2_1 U9613 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [22]), .op(n8004)
         );
  nor2_1 U9614 ( .ip1(n12376), .ip2(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .op(
        n8009) );
  not_ab_or_c_or_d U9615 ( .ip1(n12376), .ip2(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip3(n8009), .ip4(n8008), .op(n8010) );
  not_ab_or_c_or_d U9616 ( .ip1(n8011), .ip2(n12676), .ip3(n8294), .ip4(n8010), 
        .op(n8012) );
  mux2_1 U9617 ( .ip1(n8297), .ip2(n8013), .s(n8012), .op(n9139) );
  and2_1 U9618 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [22]), .op(n8022)
         );
  inv_1 U9619 ( .ip(\CORTEXM0DS_INST/u_logic/Xrdvx4 ), .op(n12213) );
  nor2_1 U9620 ( .ip1(n12051), .ip2(n12213), .op(n8016) );
  nor2_1 U9621 ( .ip1(n8014), .ip2(n8887), .op(n8015) );
  not_ab_or_c_or_d U9622 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/Itdvx4 ), 
        .ip3(n8016), .ip4(n8015), .op(n8020) );
  nand2_1 U9623 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [22]), .op(n8019)
         );
  nand2_1 U9624 ( .ip1(n8966), .ip2(\CORTEXM0DS_INST/cm0_r12 [22]), .op(n8018)
         );
  nand2_1 U9625 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [20]), .op(n8017)
         );
  not_ab_or_c_or_d U9626 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [22]), 
        .ip3(n8022), .ip4(n8021), .op(n8026) );
  nand2_1 U9627 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [22]), .op(n8025)
         );
  nand2_1 U9628 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [22]), .op(n8024)
         );
  nand2_1 U9629 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [20]), .op(n8023)
         );
  inv_1 U9630 ( .ip(n12222), .op(n9102) );
  nor2_1 U9631 ( .ip1(n8974), .ip2(n9102), .op(n8365) );
  nand2_1 U9632 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [21]), .op(n8029)
         );
  nand2_1 U9633 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [21]), .op(n8028)
         );
  nand2_1 U9634 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [21]), .op(n8027)
         );
  nand3_1 U9635 ( .ip1(n8029), .ip2(n8028), .ip3(n8027), .op(n8046) );
  nand2_1 U9636 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [21]), .ip2(n8933), .op(n8044)
         );
  nand2_1 U9637 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [21]), .op(n8033)
         );
  nand2_1 U9638 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [21]), .op(n8032)
         );
  nand2_1 U9639 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [21]), .op(n8031)
         );
  nand2_1 U9640 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [21]), .op(n8030)
         );
  nand2_1 U9641 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [19]), .op(n8037)
         );
  nand2_1 U9642 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [19]), .op(n8036)
         );
  nand2_1 U9643 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [21]), .op(n8035)
         );
  nand2_1 U9644 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [21]), .op(n8034)
         );
  not_ab_or_c_or_d U9645 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [21]), 
        .ip3(n8039), .ip4(n8038), .op(n8043) );
  nor2_1 U9646 ( .ip1(n8909), .ip2(n12213), .op(n8041) );
  and2_1 U9647 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [21]), .op(n8040)
         );
  not_ab_or_c_or_d U9648 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [21]), .ip2(n8903), 
        .ip3(n8041), .ip4(n8040), .op(n8042) );
  nand3_1 U9649 ( .ip1(n8044), .ip2(n8043), .ip3(n8042), .op(n8045) );
  not_ab_or_c_or_d U9650 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [21]), 
        .ip3(n8046), .ip4(n8045), .op(n9109) );
  nor2_1 U9651 ( .ip1(n9109), .ip2(n8292), .op(n8047) );
  not_ab_or_c_or_d U9652 ( .ip1(n8295), .ip2(\CORTEXM0DS_INST/u_logic/Wv9vx4 ), 
        .ip3(n8294), .ip4(n8047), .op(n8048) );
  mux2_1 U9653 ( .ip1(n8297), .ip2(n8013), .s(n8048), .op(n9142) );
  and2_1 U9654 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [21]), .op(n8060)
         );
  and2_1 U9655 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [21]), .op(n8054)
         );
  nand2_1 U9656 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [19]), .op(n8052)
         );
  nand2_1 U9657 ( .ip1(n8946), .ip2(n9370), .op(n8051) );
  nand2_1 U9658 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/Xrdvx4 ), .op(
        n8050) );
  nand2_1 U9659 ( .ip1(\CORTEXM0DS_INST/u_logic/Mqdvx4 ), .ip2(n8948), .op(
        n8049) );
  not_ab_or_c_or_d U9660 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [21]), .ip2(n8957), 
        .ip3(n8054), .ip4(n8053), .op(n8058) );
  nand2_1 U9661 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [21]), .op(n8057)
         );
  nand2_1 U9662 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [21]), .op(n8056)
         );
  nand2_1 U9663 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [19]), .op(n8055)
         );
  nand4_1 U9664 ( .ip1(n8058), .ip2(n8057), .ip3(n8056), .ip4(n8055), .op(
        n8059) );
  not_ab_or_c_or_d U9665 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [21]), .ip2(n8966), 
        .ip3(n8060), .ip4(n8059), .op(n11366) );
  nor2_1 U9666 ( .ip1(n8974), .ip2(n11366), .op(n8367) );
  nand2_1 U9667 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [20]), .op(n8063)
         );
  nand2_1 U9668 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [20]), .op(n8062)
         );
  nand2_1 U9669 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [20]), .op(n8061)
         );
  nand3_1 U9670 ( .ip1(n8063), .ip2(n8062), .ip3(n8061), .op(n8080) );
  nand2_1 U9671 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [20]), .ip2(n8902), .op(n8078)
         );
  nand2_1 U9672 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [20]), .op(n8067)
         );
  nand2_1 U9673 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [20]), .op(n8066)
         );
  nand2_1 U9674 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [20]), .op(n8065)
         );
  nand2_1 U9675 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [20]), .op(n8064)
         );
  nand2_1 U9676 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [18]), .op(n8071)
         );
  nand2_1 U9677 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [18]), .op(n8070)
         );
  nand2_1 U9678 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [20]), .op(n8069)
         );
  nand2_1 U9679 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [20]), .op(n8068)
         );
  not_ab_or_c_or_d U9680 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [20]), 
        .ip3(n8073), .ip4(n8072), .op(n8077) );
  and2_1 U9681 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [20]), .op(n8075)
         );
  inv_1 U9682 ( .ip(\CORTEXM0DS_INST/u_logic/Mqdvx4 ), .op(n12202) );
  nor2_1 U9683 ( .ip1(n8909), .ip2(n12202), .op(n8074) );
  not_ab_or_c_or_d U9684 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [20]), .ip2(n8903), 
        .ip3(n8075), .ip4(n8074), .op(n8076) );
  nand3_1 U9685 ( .ip1(n8078), .ip2(n8077), .ip3(n8076), .op(n8079) );
  not_ab_or_c_or_d U9686 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [20]), 
        .ip3(n8080), .ip4(n8079), .op(n11356) );
  nor2_1 U9687 ( .ip1(n11356), .ip2(n8292), .op(n8081) );
  not_ab_or_c_or_d U9688 ( .ip1(n8295), .ip2(\CORTEXM0DS_INST/u_logic/Su9vx4 ), 
        .ip3(n8294), .ip4(n8081), .op(n8082) );
  mux2_1 U9689 ( .ip1(n8297), .ip2(n8013), .s(n8082), .op(n9144) );
  and2_1 U9690 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [20]), .op(n8091)
         );
  inv_1 U9691 ( .ip(\CORTEXM0DS_INST/u_logic/Bpdvx4 ), .op(n12193) );
  nor2_1 U9692 ( .ip1(n12051), .ip2(n12193), .op(n8085) );
  nor2_1 U9693 ( .ip1(n8083), .ip2(n8887), .op(n8084) );
  not_ab_or_c_or_d U9694 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/Mqdvx4 ), 
        .ip3(n8085), .ip4(n8084), .op(n8089) );
  nand2_1 U9695 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [20]), .op(n8088)
         );
  nand2_1 U9696 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [20]), .op(n8087)
         );
  nand2_1 U9697 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [18]), .op(n8086)
         );
  not_ab_or_c_or_d U9698 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [20]), .ip2(n8966), 
        .ip3(n8091), .ip4(n8090), .op(n8095) );
  nand2_1 U9699 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [20]), .op(n8094)
         );
  nand2_1 U9700 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [20]), .op(n8093)
         );
  nand2_1 U9701 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [18]), .op(n8092)
         );
  inv_1 U9702 ( .ip(n12201), .op(n9097) );
  nor2_1 U9703 ( .ip1(n8974), .ip2(n9097), .op(n8369) );
  nand2_1 U9704 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [19]), .op(n8098)
         );
  nand2_1 U9705 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [19]), .op(n8097)
         );
  nand2_1 U9706 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [19]), .op(n8096)
         );
  nand3_1 U9707 ( .ip1(n8098), .ip2(n8097), .ip3(n8096), .op(n8115) );
  nand2_1 U9708 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [19]), .ip2(n8903), .op(n8113)
         );
  nand2_1 U9709 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [19]), .op(n8102)
         );
  nand2_1 U9710 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [19]), .op(n8101)
         );
  nand2_1 U9711 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [19]), .op(n8100)
         );
  nand2_1 U9712 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [19]), .op(n8099)
         );
  nand2_1 U9713 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [17]), .op(n8106)
         );
  nand2_1 U9714 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [19]), .op(n8105)
         );
  nand2_1 U9715 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [19]), .op(n8104)
         );
  nand2_1 U9716 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [19]), .op(n8103)
         );
  not_ab_or_c_or_d U9717 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [17]), 
        .ip3(n8108), .ip4(n8107), .op(n8112) );
  nor2_1 U9718 ( .ip1(n8909), .ip2(n12193), .op(n8110) );
  and2_1 U9719 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [19]), .op(n8109)
         );
  not_ab_or_c_or_d U9720 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [19]), .ip2(n8925), 
        .ip3(n8110), .ip4(n8109), .op(n8111) );
  nand3_1 U9721 ( .ip1(n8113), .ip2(n8112), .ip3(n8111), .op(n8114) );
  not_ab_or_c_or_d U9722 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [19]), 
        .ip3(n8115), .ip4(n8114), .op(n9108) );
  nor2_1 U9723 ( .ip1(n9108), .ip2(n8292), .op(n8116) );
  not_ab_or_c_or_d U9724 ( .ip1(n8295), .ip2(\CORTEXM0DS_INST/u_logic/Ot9vx4 ), 
        .ip3(n8294), .ip4(n8116), .op(n8117) );
  mux2_1 U9725 ( .ip1(n8297), .ip2(n8013), .s(n8117), .op(n9141) );
  and2_1 U9726 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [19]), .op(n8129)
         );
  and2_1 U9727 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [19]), .op(n8123)
         );
  nand2_1 U9728 ( .ip1(n8946), .ip2(n9369), .op(n8121) );
  nand2_1 U9729 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/Bpdvx4 ), .op(
        n8120) );
  nand2_1 U9730 ( .ip1(\CORTEXM0DS_INST/u_logic/Qndvx4 ), .ip2(n8948), .op(
        n8119) );
  nand2_1 U9731 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [17]), .op(n8118)
         );
  not_ab_or_c_or_d U9732 ( .ip1(n8966), .ip2(\CORTEXM0DS_INST/cm0_r12 [19]), 
        .ip3(n8123), .ip4(n8122), .op(n8127) );
  nand2_1 U9733 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [19]), .op(n8126)
         );
  nand2_1 U9734 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [19]), .op(n8125)
         );
  nand2_1 U9735 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [17]), .op(n8124)
         );
  nand4_1 U9736 ( .ip1(n8127), .ip2(n8126), .ip3(n8125), .ip4(n8124), .op(
        n8128) );
  not_ab_or_c_or_d U9737 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [19]), 
        .ip3(n8129), .ip4(n8128), .op(n11342) );
  nor2_1 U9738 ( .ip1(n8974), .ip2(n11342), .op(n8371) );
  nand2_1 U9739 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [18]), .op(n8132)
         );
  nand2_1 U9740 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [18]), .op(n8131)
         );
  nand2_1 U9741 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [18]), .op(n8130)
         );
  nand3_1 U9742 ( .ip1(n8132), .ip2(n8131), .ip3(n8130), .op(n8150) );
  nand2_1 U9743 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [18]), .ip2(n8903), .op(n8148)
         );
  nand2_1 U9744 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [18]), .op(n8136)
         );
  nand2_1 U9745 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [18]), .op(n8135)
         );
  nand2_1 U9746 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [18]), .op(n8134)
         );
  nand2_1 U9747 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [18]), .op(n8133)
         );
  nand2_1 U9748 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [16]), .op(n8140)
         );
  nand2_1 U9749 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [16]), .op(n8139)
         );
  nand2_1 U9750 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [18]), .op(n8138)
         );
  nand2_1 U9751 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [18]), .op(n8137)
         );
  not_ab_or_c_or_d U9752 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [18]), 
        .ip3(n8142), .ip4(n8141), .op(n8147) );
  inv_1 U9753 ( .ip(\CORTEXM0DS_INST/cm0_r14 [18]), .op(n8153) );
  nor2_1 U9754 ( .ip1(n8143), .ip2(n8153), .op(n8145) );
  inv_1 U9755 ( .ip(\CORTEXM0DS_INST/u_logic/Qndvx4 ), .op(n12183) );
  nor2_1 U9756 ( .ip1(n8909), .ip2(n12183), .op(n8144) );
  not_ab_or_c_or_d U9757 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [18]), .ip2(n8915), 
        .ip3(n8145), .ip4(n8144), .op(n8146) );
  nand3_1 U9758 ( .ip1(n8148), .ip2(n8147), .ip3(n8146), .op(n8149) );
  not_ab_or_c_or_d U9759 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [18]), 
        .ip3(n8150), .ip4(n8149), .op(n12666) );
  nor2_1 U9760 ( .ip1(n12666), .ip2(n8292), .op(n8151) );
  not_ab_or_c_or_d U9761 ( .ip1(n8295), .ip2(\CORTEXM0DS_INST/u_logic/Ks9vx4 ), 
        .ip3(n8294), .ip4(n8151), .op(n8152) );
  mux2_1 U9762 ( .ip1(n8297), .ip2(n8013), .s(n8152), .op(n9132) );
  nor2_1 U9763 ( .ip1(n8154), .ip2(n8153), .op(n8166) );
  and2_1 U9764 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [18]), .op(n8160)
         );
  nand2_1 U9765 ( .ip1(n8946), .ip2(n9368), .op(n8158) );
  nand2_1 U9766 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/Qndvx4 ), .op(
        n8157) );
  nand2_1 U9767 ( .ip1(\CORTEXM0DS_INST/u_logic/Fmdvx4 ), .ip2(n8948), .op(
        n8156) );
  nand2_1 U9768 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [16]), .op(n8155)
         );
  not_ab_or_c_or_d U9769 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [18]), .ip2(n8966), 
        .ip3(n8160), .ip4(n8159), .op(n8164) );
  nand2_1 U9770 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [18]), .op(n8163)
         );
  nand2_1 U9771 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [18]), .op(n8162)
         );
  nand2_1 U9772 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [16]), .op(n8161)
         );
  nand4_1 U9773 ( .ip1(n8164), .ip2(n8163), .ip3(n8162), .ip4(n8161), .op(
        n8165) );
  not_ab_or_c_or_d U9774 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [18]), 
        .ip3(n8166), .ip4(n8165), .op(n12175) );
  nor2_1 U9775 ( .ip1(n8974), .ip2(n12175), .op(n8373) );
  nand2_1 U9776 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [17]), .op(n8169)
         );
  nand2_1 U9777 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [17]), .op(n8168)
         );
  nand2_1 U9778 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [17]), .op(n8167)
         );
  nand3_1 U9779 ( .ip1(n8169), .ip2(n8168), .ip3(n8167), .op(n8188) );
  inv_1 U9780 ( .ip(\CORTEXM0DS_INST/u_logic/Fmdvx4 ), .op(n12172) );
  nor2_1 U9781 ( .ip1(n8909), .ip2(n12172), .op(n8170) );
  or2_1 U9782 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [17]), .ip2(n8170), .op(n8172)
         );
  or2_1 U9783 ( .ip1(n8933), .ip2(n8170), .op(n8171) );
  nand2_1 U9784 ( .ip1(n8172), .ip2(n8171), .op(n8186) );
  nand2_1 U9785 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [17]), .op(n8176)
         );
  nand2_1 U9786 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [17]), .op(n8175)
         );
  nand2_1 U9787 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [17]), .op(n8174)
         );
  nand2_1 U9788 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [17]), .op(n8173)
         );
  nand2_1 U9789 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [15]), .op(n8180)
         );
  nand2_1 U9790 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [15]), .op(n8179)
         );
  nand2_1 U9791 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [17]), .op(n8178)
         );
  nand2_1 U9792 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [17]), .op(n8177)
         );
  not_ab_or_c_or_d U9793 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [17]), 
        .ip3(n8182), .ip4(n8181), .op(n8185) );
  nand2_1 U9794 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [17]), .op(n8184)
         );
  nand2_1 U9795 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [17]), .op(n8183)
         );
  not_ab_or_c_or_d U9796 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [17]), 
        .ip3(n8188), .ip4(n8187), .op(n11316) );
  nor2_1 U9797 ( .ip1(n11316), .ip2(n8292), .op(n8189) );
  not_ab_or_c_or_d U9798 ( .ip1(n8295), .ip2(\CORTEXM0DS_INST/u_logic/Gr9vx4 ), 
        .ip3(n8294), .ip4(n8189), .op(n8190) );
  mux2_1 U9799 ( .ip1(n8297), .ip2(n8013), .s(n8190), .op(n9140) );
  and2_1 U9800 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [17]), .op(n8202)
         );
  and2_1 U9801 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [17]), .op(n8196)
         );
  nand2_1 U9802 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [15]), .op(n8194)
         );
  nand2_1 U9803 ( .ip1(n8946), .ip2(n9434), .op(n8193) );
  nand2_1 U9804 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/Fmdvx4 ), .op(
        n8192) );
  nand2_1 U9805 ( .ip1(\CORTEXM0DS_INST/u_logic/Ukdvx4 ), .ip2(n8948), .op(
        n8191) );
  not_ab_or_c_or_d U9806 ( .ip1(n8966), .ip2(\CORTEXM0DS_INST/cm0_r12 [17]), 
        .ip3(n8196), .ip4(n8195), .op(n8200) );
  nand2_1 U9807 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [17]), .op(n8199)
         );
  nand2_1 U9808 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [17]), .op(n8198)
         );
  nand2_1 U9809 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [15]), .op(n8197)
         );
  nand4_1 U9810 ( .ip1(n8200), .ip2(n8199), .ip3(n8198), .ip4(n8197), .op(
        n8201) );
  not_ab_or_c_or_d U9811 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [17]), .ip2(n8957), 
        .ip3(n8202), .ip4(n8201), .op(n11319) );
  nor2_1 U9812 ( .ip1(n8974), .ip2(n11319), .op(n8375) );
  nand2_1 U9813 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [16]), .op(n8205)
         );
  nand2_1 U9814 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [16]), .op(n8204)
         );
  nand2_1 U9815 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [16]), .op(n8203)
         );
  nand3_1 U9816 ( .ip1(n8205), .ip2(n8204), .ip3(n8203), .op(n8222) );
  nand2_1 U9817 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [16]), .ip2(n8925), .op(n8220)
         );
  nand2_1 U9818 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [16]), .op(n8209)
         );
  nand2_1 U9819 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [16]), .op(n8208)
         );
  nand2_1 U9820 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [16]), .op(n8207)
         );
  nand2_1 U9821 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [16]), .op(n8206)
         );
  nand2_1 U9822 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [14]), .op(n8213)
         );
  nand2_1 U9823 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [14]), .op(n8212)
         );
  nand2_1 U9824 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [16]), .op(n8211)
         );
  nand2_1 U9825 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [16]), .op(n8210)
         );
  not_ab_or_c_or_d U9826 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [16]), 
        .ip3(n8215), .ip4(n8214), .op(n8219) );
  inv_1 U9827 ( .ip(\CORTEXM0DS_INST/u_logic/Ukdvx4 ), .op(n12163) );
  nor2_1 U9828 ( .ip1(n8909), .ip2(n12163), .op(n8217) );
  and2_1 U9829 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [16]), .op(n8216)
         );
  not_ab_or_c_or_d U9830 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [16]), .ip2(n8917), 
        .ip3(n8217), .ip4(n8216), .op(n8218) );
  nand3_1 U9831 ( .ip1(n8220), .ip2(n8219), .ip3(n8218), .op(n8221) );
  not_ab_or_c_or_d U9832 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [16]), 
        .ip3(n8222), .ip4(n8221), .op(n11308) );
  nor2_1 U9833 ( .ip1(n11308), .ip2(n8292), .op(n8223) );
  not_ab_or_c_or_d U9834 ( .ip1(n8295), .ip2(\CORTEXM0DS_INST/u_logic/Cq9vx4 ), 
        .ip3(n8294), .ip4(n8223), .op(n8224) );
  mux2_1 U9835 ( .ip1(n8297), .ip2(n8013), .s(n8224), .op(n9134) );
  and2_1 U9836 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [16]), .op(n8232)
         );
  inv_1 U9837 ( .ip(n9432), .op(n9390) );
  nor2_1 U9838 ( .ip1(n9390), .ip2(n8887), .op(n8226) );
  inv_1 U9839 ( .ip(\CORTEXM0DS_INST/u_logic/Jjdvx4 ), .op(n8240) );
  nor2_1 U9840 ( .ip1(n12051), .ip2(n8240), .op(n8225) );
  not_ab_or_c_or_d U9841 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [14]), 
        .ip3(n8226), .ip4(n8225), .op(n8230) );
  nand2_1 U9842 ( .ip1(n8966), .ip2(\CORTEXM0DS_INST/cm0_r12 [16]), .op(n8229)
         );
  nand2_1 U9843 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [16]), .op(n8228)
         );
  nand2_1 U9844 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/Ukdvx4 ), .op(
        n8227) );
  not_ab_or_c_or_d U9845 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [16]), .ip2(n8957), 
        .ip3(n8232), .ip4(n8231), .op(n8236) );
  nand2_1 U9846 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [16]), .op(n8235)
         );
  nand2_1 U9847 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [16]), .op(n8234)
         );
  nand2_1 U9848 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [14]), .op(n8233)
         );
  nand4_1 U9849 ( .ip1(n8236), .ip2(n8235), .ip3(n8234), .ip4(n8233), .op(
        n9135) );
  inv_1 U9850 ( .ip(n9135), .op(n12159) );
  nor2_1 U9851 ( .ip1(n8974), .ip2(n12159), .op(n8377) );
  nand2_1 U9852 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [15]), .op(n8239)
         );
  nand2_1 U9853 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [15]), .op(n8238)
         );
  nand2_1 U9854 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [15]), .op(n8237)
         );
  nand3_1 U9855 ( .ip1(n8239), .ip2(n8238), .ip3(n8237), .op(n8257) );
  and2_1 U9856 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [13]), .op(n8242)
         );
  nor2_1 U9857 ( .ip1(n8909), .ip2(n8240), .op(n8241) );
  not_ab_or_c_or_d U9858 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [15]), .ip2(n8910), 
        .ip3(n8242), .ip4(n8241), .op(n8255) );
  nand2_1 U9859 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [15]), .op(n8246)
         );
  nand2_1 U9860 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [15]), .op(n8245)
         );
  nand2_1 U9861 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [15]), .op(n8244)
         );
  nand2_1 U9862 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [15]), .op(n8243)
         );
  nand2_1 U9863 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [15]), .op(n8249)
         );
  nand2_1 U9864 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [15]), .op(n8248)
         );
  nand2_1 U9865 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [15]), .op(n8247)
         );
  nand3_1 U9866 ( .ip1(n8249), .ip2(n8248), .ip3(n8247), .op(n8250) );
  not_ab_or_c_or_d U9867 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [15]), 
        .ip3(n8251), .ip4(n8250), .op(n8254) );
  nand2_1 U9868 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [13]), .op(n8253)
         );
  nand2_1 U9869 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [15]), .op(n8252)
         );
  not_ab_or_c_or_d U9870 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [15]), 
        .ip3(n8257), .ip4(n8256), .op(n9858) );
  nor2_1 U9871 ( .ip1(n9858), .ip2(n8292), .op(n8258) );
  not_ab_or_c_or_d U9872 ( .ip1(n8295), .ip2(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), 
        .ip3(n8294), .ip4(n8258), .op(n8259) );
  mux2_1 U9873 ( .ip1(n8297), .ip2(n8013), .s(n8259), .op(n11540) );
  and2_1 U9874 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [15]), .op(n8271)
         );
  and2_1 U9875 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [15]), .op(n8265)
         );
  nand2_1 U9876 ( .ip1(\CORTEXM0DS_INST/u_logic/Yhdvx4 ), .ip2(n8948), .op(
        n8263) );
  nand2_1 U9877 ( .ip1(n8946), .ip2(n9428), .op(n8262) );
  nand2_1 U9878 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/Jjdvx4 ), .op(
        n8261) );
  nand2_1 U9879 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [13]), .op(n8260)
         );
  not_ab_or_c_or_d U9880 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [15]), .ip2(n8966), 
        .ip3(n8265), .ip4(n8264), .op(n8269) );
  nand2_1 U9881 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [15]), .op(n8268)
         );
  nand2_1 U9882 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [15]), .op(n8267)
         );
  nand2_1 U9883 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [13]), .op(n8266)
         );
  nand4_1 U9884 ( .ip1(n8269), .ip2(n8268), .ip3(n8267), .ip4(n8266), .op(
        n8270) );
  not_ab_or_c_or_d U9885 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [15]), 
        .ip3(n8271), .ip4(n8270), .op(n10964) );
  nor2_1 U9886 ( .ip1(n8974), .ip2(n10964), .op(n8379) );
  nand2_1 U9887 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [14]), .op(n8274)
         );
  nand2_1 U9888 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [14]), .op(n8273)
         );
  nand2_1 U9889 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [14]), .op(n8272)
         );
  nand3_1 U9890 ( .ip1(n8274), .ip2(n8273), .ip3(n8272), .op(n8291) );
  nand2_1 U9891 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [14]), .ip2(n8910), .op(n8289)
         );
  nand2_1 U9892 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [14]), .op(n8278)
         );
  nand2_1 U9893 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [14]), .op(n8277)
         );
  nand2_1 U9894 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [14]), .op(n8276)
         );
  nand2_1 U9895 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [14]), .op(n8275)
         );
  nand2_1 U9896 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [12]), .op(n8282)
         );
  nand2_1 U9897 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [12]), .op(n8281)
         );
  nand2_1 U9898 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [14]), .op(n8280)
         );
  nand2_1 U9899 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [14]), .op(n8279)
         );
  not_ab_or_c_or_d U9900 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [14]), 
        .ip3(n8284), .ip4(n8283), .op(n8288) );
  and2_1 U9901 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [14]), .op(n8286)
         );
  and2_1 U9902 ( .ip1(n8853), .ip2(\CORTEXM0DS_INST/u_logic/Yhdvx4 ), .op(
        n8285) );
  not_ab_or_c_or_d U9903 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [14]), .ip2(n8903), 
        .ip3(n8286), .ip4(n8285), .op(n8287) );
  nand3_1 U9904 ( .ip1(n8289), .ip2(n8288), .ip3(n8287), .op(n8290) );
  not_ab_or_c_or_d U9905 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [14]), 
        .ip3(n8291), .ip4(n8290), .op(n11295) );
  nor2_1 U9906 ( .ip1(n11295), .ip2(n8292), .op(n8293) );
  not_ab_or_c_or_d U9907 ( .ip1(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .ip2(n8295), 
        .ip3(n8294), .ip4(n8293), .op(n8296) );
  mux2_1 U9908 ( .ip1(n8297), .ip2(n8013), .s(n8296), .op(n9147) );
  and2_1 U9909 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [14]), .op(n8306)
         );
  nor2_1 U9910 ( .ip1(n9419), .ip2(n8887), .op(n8300) );
  nor2_1 U9911 ( .ip1(n12051), .ip2(n8298), .op(n8299) );
  not_ab_or_c_or_d U9912 ( .ip1(\CORTEXM0DS_INST/u_logic/Yhdvx4 ), .ip2(n8947), 
        .ip3(n8300), .ip4(n8299), .op(n8304) );
  nand2_1 U9913 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [14]), .op(n8303)
         );
  nand2_1 U9914 ( .ip1(n8966), .ip2(\CORTEXM0DS_INST/cm0_r12 [14]), .op(n8302)
         );
  nand2_1 U9915 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [12]), .op(n8301)
         );
  not_ab_or_c_or_d U9916 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [14]), .ip2(n8957), 
        .ip3(n8306), .ip4(n8305), .op(n8310) );
  nand2_1 U9917 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [14]), .op(n8309)
         );
  nand2_1 U9918 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [14]), .op(n8308)
         );
  nand2_1 U9919 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [12]), .op(n8307)
         );
  nand4_1 U9920 ( .ip1(n8310), .ip2(n8309), .ip3(n8308), .ip4(n8307), .op(
        n9148) );
  inv_1 U9921 ( .ip(n9148), .op(n9810) );
  nor2_1 U9922 ( .ip1(n8974), .ip2(n9810), .op(n8381) );
  fulladder U9923 ( .a(n9137), .b(n8312), .ci(n8311), .co(n8380), .s(n8382) );
  inv_1 U9924 ( .ip(n12259), .op(n11431) );
  nand2_1 U9925 ( .ip1(n11431), .ip2(n8969), .op(n8313) );
  xor2_1 U9926 ( .ip1(n11427), .ip2(n8313), .op(n8391) );
  nand2_1 U9927 ( .ip1(n8392), .ip2(n8391), .op(n8314) );
  nand2_1 U9928 ( .ip1(n8315), .ip2(n8314), .op(n8357) );
  inv_1 U9929 ( .ip(n9193), .op(n9196) );
  and2_1 U9930 ( .ip1(n8969), .ip2(n12274), .op(n8316) );
  xor2_1 U9931 ( .ip1(n9196), .ip2(n8316), .op(n8356) );
  nor2_1 U9932 ( .ip1(n8357), .ip2(n8356), .op(n8317) );
  nor2_1 U9933 ( .ip1(n8318), .ip2(n8317), .op(n8971) );
  nand2_1 U9934 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [28]), .op(n8321)
         );
  nand2_1 U9935 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [28]), .op(n8320)
         );
  nand2_1 U9936 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [28]), .op(n8319)
         );
  nand3_1 U9937 ( .ip1(n8321), .ip2(n8320), .ip3(n8319), .op(n8340) );
  and2_1 U9938 ( .ip1(n8853), .ip2(\CORTEXM0DS_INST/u_logic/W1evx4 ), .op(
        n8322) );
  or2_1 U9939 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [28]), .ip2(n8322), .op(n8324)
         );
  or2_1 U9940 ( .ip1(n8903), .ip2(n8322), .op(n8323) );
  nand2_1 U9941 ( .ip1(n8324), .ip2(n8323), .op(n8338) );
  nand2_1 U9942 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [28]), .op(n8328)
         );
  nand2_1 U9943 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [28]), .op(n8327)
         );
  nand2_1 U9944 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [28]), .op(n8326)
         );
  nand2_1 U9945 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [28]), .op(n8325)
         );
  nand2_1 U9946 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [26]), .op(n8332)
         );
  nand2_1 U9947 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [26]), .op(n8331)
         );
  nand2_1 U9948 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [28]), .op(n8330)
         );
  nand2_1 U9949 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [28]), .op(n8329)
         );
  not_ab_or_c_or_d U9950 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [28]), 
        .ip3(n8334), .ip4(n8333), .op(n8337) );
  nand2_1 U9951 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [28]), .op(n8336)
         );
  nand2_1 U9952 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [28]), .op(n8335)
         );
  not_ab_or_c_or_d U9953 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [28]), 
        .ip3(n8340), .ip4(n8339), .op(n11009) );
  mux2_1 U9954 ( .ip1(n8342), .ip2(n8341), .s(n11009), .op(n9159) );
  inv_1 U9955 ( .ip(n9159), .op(n9163) );
  and2_1 U9956 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [28]), .op(n8350)
         );
  nor2_1 U9957 ( .ip1(n9317), .ip2(n8887), .op(n8344) );
  nor2_1 U9958 ( .ip1(n12051), .ip2(n12275), .op(n8343) );
  not_ab_or_c_or_d U9959 ( .ip1(\CORTEXM0DS_INST/u_logic/W1evx4 ), .ip2(n8947), 
        .ip3(n8344), .ip4(n8343), .op(n8348) );
  nand2_1 U9960 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [28]), .op(n8347)
         );
  nand2_1 U9961 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [28]), .op(n8346)
         );
  nand2_1 U9962 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [26]), .op(n8345)
         );
  not_ab_or_c_or_d U9963 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [28]), 
        .ip3(n8350), .ip4(n8349), .op(n8354) );
  nand2_1 U9964 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [28]), .op(n8353)
         );
  nand2_1 U9965 ( .ip1(n8966), .ip2(\CORTEXM0DS_INST/cm0_r12 [28]), .op(n8352)
         );
  nand2_1 U9966 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [26]), .op(n8351)
         );
  inv_1 U9967 ( .ip(n9160), .op(n8395) );
  nor2_1 U9968 ( .ip1(n8974), .ip2(n8395), .op(n8355) );
  xor2_1 U9969 ( .ip1(n9163), .ip2(n8355), .op(n8970) );
  xor2_1 U9970 ( .ip1(n8971), .ip2(n8970), .op(n8982) );
  xor2_1 U9971 ( .ip1(n8357), .ip2(n8356), .op(n9016) );
  inv_1 U9972 ( .ip(n9016), .op(n8393) );
  fulladder U9973 ( .a(n9100), .b(n8359), .ci(n8358), .co(n8392), .s(n9018) );
  fulladder U9974 ( .a(n9047), .b(n8361), .ci(n8360), .co(n8358), .s(n9241) );
  fulladder U9975 ( .a(n9056), .b(n8363), .ci(n8362), .co(n8360), .s(n9206) );
  inv_1 U9976 ( .ip(n9206), .op(n8389) );
  fulladder U9977 ( .a(n9139), .b(n8365), .ci(n8364), .co(n8362), .s(n9243) );
  fulladder U9978 ( .a(n9142), .b(n8367), .ci(n8366), .co(n8364), .s(n9233) );
  inv_1 U9979 ( .ip(n9233), .op(n8388) );
  fulladder U9980 ( .a(n9144), .b(n8369), .ci(n8368), .co(n8366), .s(n9245) );
  fulladder U9981 ( .a(n9141), .b(n8371), .ci(n8370), .co(n8368), .s(n9247) );
  inv_1 U9982 ( .ip(n9247), .op(n8387) );
  fulladder U9983 ( .a(n9132), .b(n8373), .ci(n8372), .co(n8370), .s(n9210) );
  fulladder U9984 ( .a(n9140), .b(n8375), .ci(n8374), .co(n8372), .s(n9226) );
  inv_1 U9985 ( .ip(n9226), .op(n8386) );
  fulladder U9986 ( .a(n9134), .b(n8377), .ci(n8376), .co(n8374), .s(n9208) );
  fulladder U9987 ( .a(n11540), .b(n8379), .ci(n8378), .co(n8376), .s(n9228)
         );
  inv_1 U9988 ( .ip(n9228), .op(n8385) );
  fulladder U9989 ( .a(n9147), .b(n8381), .ci(n8380), .co(n8378), .s(n9212) );
  inv_1 U9990 ( .ip(n8382), .op(n8384) );
  nor2_1 U9991 ( .ip1(n8384), .ip2(n8383), .op(n9211) );
  nand2_1 U9992 ( .ip1(n9212), .ip2(n9211), .op(n9227) );
  nor2_1 U9993 ( .ip1(n8385), .ip2(n9227), .op(n9207) );
  nand2_1 U9994 ( .ip1(n9208), .ip2(n9207), .op(n9225) );
  nor2_1 U9995 ( .ip1(n8386), .ip2(n9225), .op(n9209) );
  nand2_1 U9996 ( .ip1(n9210), .ip2(n9209), .op(n9246) );
  nor2_1 U9997 ( .ip1(n8387), .ip2(n9246), .op(n9244) );
  nand2_1 U9998 ( .ip1(n9245), .ip2(n9244), .op(n9232) );
  nor2_1 U9999 ( .ip1(n8388), .ip2(n9232), .op(n9242) );
  nand2_1 U10000 ( .ip1(n9243), .ip2(n9242), .op(n9205) );
  nor2_1 U10001 ( .ip1(n8389), .ip2(n9205), .op(n9240) );
  nand2_1 U10002 ( .ip1(n9241), .ip2(n9240), .op(n9017) );
  inv_1 U10003 ( .ip(n9017), .op(n8390) );
  nand2_1 U10004 ( .ip1(n9018), .ip2(n8390), .op(n9251) );
  xnor2_1 U10005 ( .ip1(n8392), .ip2(n8391), .op(n9250) );
  nor2_1 U10006 ( .ip1(n9251), .ip2(n9250), .op(n9015) );
  nand2_1 U10007 ( .ip1(n8393), .ip2(n9015), .op(n8983) );
  xor2_1 U10008 ( .ip1(n8982), .ip2(n8983), .op(n10071) );
  inv_1 U10009 ( .ip(\CORTEXM0DS_INST/vis_pc [27]), .op(n10072) );
  nand2_1 U10010 ( .ip1(n12226), .ip2(\CORTEXM0DS_INST/vis_pc [4]), .op(n12239) );
  nor2_1 U10011 ( .ip1(n12239), .ip2(n12244), .op(n12291) );
  nand2_1 U10012 ( .ip1(n12291), .ip2(\CORTEXM0DS_INST/vis_pc [6]), .op(n12292) );
  nand2_1 U10013 ( .ip1(n8394), .ip2(\CORTEXM0DS_INST/vis_pc [12]), .op(n9937)
         );
  nor2_1 U10014 ( .ip1(n12292), .ip2(n9937), .op(n9807) );
  nand2_1 U10015 ( .ip1(n9807), .ip2(\CORTEXM0DS_INST/vis_pc [13]), .op(n10966) );
  inv_1 U10016 ( .ip(\CORTEXM0DS_INST/vis_pc [14]), .op(n10965) );
  nor2_1 U10017 ( .ip1(n10966), .ip2(n10965), .op(n12155) );
  nand2_1 U10018 ( .ip1(n12155), .ip2(\CORTEXM0DS_INST/vis_pc [15]), .op(
        n12167) );
  inv_1 U10019 ( .ip(\CORTEXM0DS_INST/vis_pc [16]), .op(n12166) );
  nor2_1 U10020 ( .ip1(n12167), .ip2(n12166), .op(n12176) );
  nand3_1 U10021 ( .ip1(\CORTEXM0DS_INST/vis_pc [17]), .ip2(
        \CORTEXM0DS_INST/vis_pc [18]), .ip3(n12176), .op(n12197) );
  inv_1 U10022 ( .ip(\CORTEXM0DS_INST/vis_pc [19]), .op(n12196) );
  nor2_1 U10023 ( .ip1(n12197), .ip2(n12196), .op(n12205) );
  nand2_1 U10024 ( .ip1(n12205), .ip2(\CORTEXM0DS_INST/vis_pc [20]), .op(
        n12218) );
  inv_1 U10025 ( .ip(\CORTEXM0DS_INST/vis_pc [21]), .op(n12217) );
  nor2_1 U10026 ( .ip1(n12218), .ip2(n12217), .op(n12216) );
  nand2_1 U10027 ( .ip1(n12216), .ip2(\CORTEXM0DS_INST/vis_pc [22]), .op(
        n12308) );
  inv_1 U10028 ( .ip(\CORTEXM0DS_INST/vis_pc [23]), .op(n12307) );
  nor2_1 U10029 ( .ip1(n12308), .ip2(n12307), .op(n12306) );
  nand2_1 U10030 ( .ip1(n12306), .ip2(\CORTEXM0DS_INST/vis_pc [24]), .op(
        n12258) );
  inv_1 U10031 ( .ip(\CORTEXM0DS_INST/vis_pc [25]), .op(n12257) );
  nor2_1 U10032 ( .ip1(n12258), .ip2(n12257), .op(n12266) );
  nand2_1 U10033 ( .ip1(n12266), .ip2(\CORTEXM0DS_INST/vis_pc [26]), .op(
        n12267) );
  nand3_1 U10034 ( .ip1(\CORTEXM0DS_INST/vis_pc [27]), .ip2(n12266), .ip3(
        \CORTEXM0DS_INST/vis_pc [26]), .op(n9821) );
  inv_1 U10035 ( .ip(n9821), .op(n9814) );
  not_ab_or_c_or_d U10036 ( .ip1(n10072), .ip2(n12267), .ip3(n9814), .ip4(
        n12305), .op(n8397) );
  nor2_1 U10037 ( .ip1(n8395), .ip2(n12295), .op(n8396) );
  not_ab_or_c_or_d U10038 ( .ip1(n12300), .ip2(n10071), .ip3(n8397), .ip4(
        n8396), .op(\CORTEXM0DS_INST/u_logic/V2qvx4 ) );
  or2_1 U10039 ( .ip1(n12317), .ip2(\CORTEXM0DS_INST/u_logic/V2qvx4 ), .op(
        n8398) );
  nand4_1 U10040 ( .ip1(n8401), .ip2(n8400), .ip3(n8399), .ip4(n8398), .op(
        n6079) );
  nor2_1 U10041 ( .ip1(\CORTEXM0DS_INST/u_logic/Z7hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/B5hvx4 ), .op(n8402) );
  nand2_1 U10042 ( .ip1(n8402), .ip2(n10208), .op(n11775) );
  inv_1 U10043 ( .ip(\interconnect_ip_inst/i_ahb_U_mux_hsel_prev [1]), .op(
        n8800) );
  inv_1 U10044 ( .ip(n8403), .op(n8798) );
  nor3_1 U10045 ( .ip1(n8800), .ip2(n8798), .ip3(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [2]), .op(n5920) );
  inv_1 U10046 ( .ip(n5920), .op(n8499) );
  nor4_1 U10047 ( .ip1(n12685), .ip2(n11839), .ip3(n11775), .ip4(n8499), .op(
        n12694) );
  nand2_1 U10048 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n10975), .op(
        n12352) );
  inv_1 U10049 ( .ip(n12352), .op(n9749) );
  nand3_1 U10050 ( .ip1(n11186), .ip2(n10729), .ip3(n12095), .op(n8404) );
  not_ab_or_c_or_d U10051 ( .ip1(n12615), .ip2(n8404), .ip3(n12075), .ip4(
        n10811), .op(n8406) );
  inv_1 U10052 ( .ip(n9664), .op(n10915) );
  nor2_1 U10053 ( .ip1(n10915), .ip2(n9620), .op(n8405) );
  not_ab_or_c_or_d U10054 ( .ip1(n9749), .ip2(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip3(n8406), .ip4(n8405), .op(n8412) );
  inv_1 U10055 ( .ip(n11736), .op(n11085) );
  inv_1 U10056 ( .ip(n11771), .op(n11726) );
  nand2_1 U10057 ( .ip1(n11744), .ip2(n11207), .op(n8408) );
  nor2_1 U10058 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(n10770), .op(
        n10778) );
  nand2_1 U10059 ( .ip1(n10778), .ip2(n10547), .op(n8407) );
  nand2_1 U10060 ( .ip1(n8408), .ip2(n8407), .op(n8409) );
  nand2_1 U10061 ( .ip1(n11726), .ip2(n8409), .op(n8411) );
  nand2_1 U10062 ( .ip1(n12606), .ip2(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .op(
        n8410) );
  nand4_1 U10063 ( .ip1(n8412), .ip2(n11085), .ip3(n8411), .ip4(n8410), .op(
        n2135) );
  nor2_1 U10064 ( .ip1(\CORTEXM0DS_INST/u_logic/Ho8vx4 ), .ip2(n12075), .op(
        n8415) );
  nor2_1 U10065 ( .ip1(n11038), .ip2(n12592), .op(n12279) );
  nand2_1 U10066 ( .ip1(n12279), .ip2(n12588), .op(n12332) );
  inv_1 U10067 ( .ip(n12332), .op(n8414) );
  nor2_1 U10068 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n10506), .op(
        n10827) );
  nand2_1 U10069 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(n10827), .op(
        n10792) );
  inv_1 U10070 ( .ip(n10792), .op(n12339) );
  nor2_1 U10071 ( .ip1(n12096), .ip2(n8826), .op(n8413) );
  not_ab_or_c_or_d U10072 ( .ip1(n8415), .ip2(n8414), .ip3(n12339), .ip4(n8413), .op(n8423) );
  nand2_1 U10073 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Aj9vx4 ), .op(n12073) );
  inv_1 U10074 ( .ip(n12073), .op(n10512) );
  inv_1 U10075 ( .ip(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .op(n12584) );
  nand2_1 U10076 ( .ip1(n10512), .ip2(n12584), .op(n10515) );
  inv_1 U10077 ( .ip(n10515), .op(n9623) );
  nand2_1 U10078 ( .ip1(n12588), .ip2(n9754), .op(n10869) );
  inv_1 U10079 ( .ip(n10869), .op(n8712) );
  inv_1 U10080 ( .ip(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .op(n12530) );
  nand2_1 U10081 ( .ip1(n12530), .ip2(n12588), .op(n10612) );
  inv_1 U10082 ( .ip(n10612), .op(n10455) );
  inv_1 U10083 ( .ip(\CORTEXM0DS_INST/u_logic/R89vx4 ), .op(n12570) );
  not_ab_or_c_or_d U10084 ( .ip1(n10455), .ip2(n12570), .ip3(n11038), .ip4(
        n10782), .op(n8418) );
  nor2_1 U10085 ( .ip1(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Cf9vx4 ), .op(n9566) );
  nand2_1 U10086 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n12530), .op(
        n10749) );
  nor3_1 U10087 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Ho8vx4 ), .ip3(n10749), .op(n10717) );
  nand2_1 U10088 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(n12584), .op(
        n10742) );
  inv_1 U10089 ( .ip(n10742), .op(n10757) );
  inv_1 U10090 ( .ip(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .op(n9754) );
  nand2_1 U10091 ( .ip1(\CORTEXM0DS_INST/u_logic/R89vx4 ), .ip2(n12564), .op(
        n10925) );
  nand3_1 U10092 ( .ip1(n10757), .ip2(n9754), .ip3(n10925), .op(n10693) );
  nor3_1 U10093 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n10693), .ip3(
        n12073), .op(n8416) );
  not_ab_or_c_or_d U10094 ( .ip1(n9566), .ip2(n10512), .ip3(n10717), .ip4(
        n8416), .op(n8417) );
  nand2_1 U10095 ( .ip1(n11736), .ip2(n11771), .op(n11758) );
  nand2_1 U10096 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n12580), .op(
        n10751) );
  inv_1 U10097 ( .ip(n10751), .op(n10871) );
  nand3_1 U10098 ( .ip1(n10871), .ip2(n10512), .ip3(n12075), .op(n10440) );
  nand3_1 U10099 ( .ip1(n8417), .ip2(n11758), .ip3(n10440), .op(n8466) );
  not_ab_or_c_or_d U10100 ( .ip1(n9623), .ip2(n8712), .ip3(n8418), .ip4(n8466), 
        .op(n8422) );
  nand2_1 U10101 ( .ip1(n8419), .ip2(n11715), .op(n8446) );
  nand2_1 U10102 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Mc9vx4 ), .op(n12327) );
  inv_1 U10103 ( .ip(n12327), .op(n10767) );
  nor2_1 U10104 ( .ip1(n10767), .ip2(n10749), .op(n8435) );
  inv_1 U10105 ( .ip(n10701), .op(n10517) );
  nand2_1 U10106 ( .ip1(n10517), .ip2(n12592), .op(n10622) );
  inv_1 U10107 ( .ip(n10622), .op(n8436) );
  not_ab_or_c_or_d U10108 ( .ip1(n10827), .ip2(n9754), .ip3(n8435), .ip4(n8436), .op(n8420) );
  or2_1 U10109 ( .ip1(\CORTEXM0DS_INST/u_logic/Ho8vx4 ), .ip2(n8420), .op(
        n8421) );
  nand4_1 U10110 ( .ip1(n8423), .ip2(n8422), .ip3(n8446), .ip4(n8421), .op(
        n3368) );
  nand2_1 U10111 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Kg9vx4 ), .op(n10605) );
  nor2_1 U10112 ( .ip1(n10782), .ip2(n10605), .op(n10696) );
  nand2_1 U10113 ( .ip1(n10701), .ip2(n11053), .op(n8425) );
  nor2_1 U10114 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n10749), .op(
        n12280) );
  inv_1 U10115 ( .ip(n12280), .op(n8424) );
  nand2_1 U10116 ( .ip1(n10454), .ip2(n12530), .op(n9695) );
  nand2_1 U10117 ( .ip1(n8424), .ip2(n9695), .op(n10932) );
  nand2_1 U10118 ( .ip1(n8425), .ip2(n10932), .op(n9668) );
  or2_1 U10119 ( .ip1(n9668), .ip2(\CORTEXM0DS_INST/u_logic/Ho8vx4 ), .op(
        n8431) );
  nand3_1 U10120 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/R89vx4 ), .op(n8426) );
  nand2_1 U10121 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n8426), .op(
        n8428) );
  nand2_1 U10122 ( .ip1(\CORTEXM0DS_INST/u_logic/K79vx4 ), .ip2(n12570), .op(
        n10882) );
  inv_1 U10123 ( .ip(n10882), .op(n8427) );
  nor2_1 U10124 ( .ip1(n12580), .ip2(n9754), .op(n12278) );
  nand2_1 U10125 ( .ip1(n8427), .ip2(n12278), .op(n10669) );
  nand2_1 U10126 ( .ip1(n9463), .ip2(n10669), .op(n12349) );
  nand3_1 U10127 ( .ip1(n8428), .ip2(n10827), .ip3(n12349), .op(n8429) );
  or2_1 U10128 ( .ip1(n8429), .ip2(\CORTEXM0DS_INST/u_logic/Ho8vx4 ), .op(
        n8430) );
  nand2_1 U10129 ( .ip1(n8431), .ip2(n8430), .op(n8442) );
  nand3_1 U10130 ( .ip1(n10830), .ip2(n10679), .ip3(n11730), .op(n10479) );
  nor2_1 U10131 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n10479), .op(
        n11756) );
  inv_1 U10132 ( .ip(\CORTEXM0DS_INST/u_logic/P39vx4 ), .op(n12550) );
  nand2_1 U10133 ( .ip1(n11756), .ip2(n12550), .op(n10690) );
  nand3_1 U10134 ( .ip1(n8712), .ip2(n10512), .ip3(n12580), .op(n8432) );
  nand3_1 U10135 ( .ip1(n8813), .ip2(n10690), .ip3(n8432), .op(n8441) );
  or2_1 U10136 ( .ip1(n9934), .ip2(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .op(
        n8434) );
  nand2_1 U10137 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n10969), .op(
        n9519) );
  or2_1 U10138 ( .ip1(n9519), .ip2(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .op(
        n8433) );
  nand2_1 U10139 ( .ip1(n8434), .ip2(n8433), .op(n9725) );
  nand2_1 U10140 ( .ip1(n11756), .ip2(n12625), .op(n9680) );
  inv_1 U10141 ( .ip(n9680), .op(n8439) );
  nor2_1 U10142 ( .ip1(n8436), .ip2(n8435), .op(n8437) );
  nor2_1 U10143 ( .ip1(n8437), .ip2(n12329), .op(n8438) );
  not_ab_or_c_or_d U10144 ( .ip1(n9725), .ip2(n10776), .ip3(n8439), .ip4(n8438), .op(n8472) );
  nor2_1 U10145 ( .ip1(n11754), .ip2(n9620), .op(n9827) );
  nand2_1 U10146 ( .ip1(n9827), .ip2(n6210), .op(n9572) );
  nand4_1 U10147 ( .ip1(n8472), .ip2(n11758), .ip3(n9572), .ip4(n10440), .op(
        n8440) );
  nor4_1 U10148 ( .ip1(n10696), .ip2(n8442), .ip3(n8441), .ip4(n8440), .op(
        n12088) );
  nor2_1 U10149 ( .ip1(n9700), .ip2(n11035), .op(n10584) );
  nor3_1 U10150 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n10770), .ip3(
        n10588), .op(n8444) );
  nor2_1 U10151 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n12073), .op(
        n10511) );
  inv_1 U10152 ( .ip(n10511), .op(n11029) );
  nor2_1 U10153 ( .ip1(n12075), .ip2(n11029), .op(n8443) );
  not_ab_or_c_or_d U10154 ( .ip1(n10584), .ip2(n12625), .ip3(n8444), .ip4(
        n8443), .op(n8450) );
  nand2_1 U10155 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(n11730), .op(
        n12621) );
  nor3_1 U10156 ( .ip1(n10771), .ip2(n10770), .ip3(n12621), .op(n8811) );
  inv_1 U10157 ( .ip(n12072), .op(n11161) );
  nand2_1 U10158 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n11161), .op(
        n8447) );
  nor3_1 U10159 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n12614), .ip3(
        n10943), .op(n8445) );
  nor2_1 U10160 ( .ip1(n10027), .ip2(n8445), .op(n12081) );
  nand3_1 U10161 ( .ip1(n8447), .ip2(n12081), .ip3(n8446), .op(n8448) );
  not_ab_or_c_or_d U10162 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(
        n10717), .ip3(n8811), .ip4(n8448), .op(n8449) );
  inv_1 U10163 ( .ip(n10908), .op(n10820) );
  nand2_1 U10164 ( .ip1(n10820), .ip2(n9749), .op(n12080) );
  nand4_1 U10165 ( .ip1(n12088), .ip2(n8450), .ip3(n8449), .ip4(n12080), .op(
        n4626) );
  inv_1 U10166 ( .ip(n11186), .op(n12388) );
  nand2_1 U10167 ( .ip1(n10729), .ip2(n12095), .op(n11213) );
  nor3_1 U10168 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n12388), .ip3(
        n11213), .op(n8810) );
  nor2_1 U10169 ( .ip1(n12075), .ip2(n12530), .op(n10617) );
  nand3_1 U10170 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n10617), .ip3(
        n12588), .op(n10707) );
  inv_1 U10171 ( .ip(n10707), .op(n10753) );
  nor3_1 U10172 ( .ip1(n12614), .ip2(n9620), .ip3(n8451), .op(n8452) );
  not_ab_or_c_or_d U10173 ( .ip1(n8810), .ip2(\CORTEXM0DS_INST/u_logic/Ho8vx4 ), .ip3(n10753), .ip4(n8452), .op(n8471) );
  nor2_1 U10174 ( .ip1(n10547), .ip2(n11729), .op(n10810) );
  nor2_1 U10175 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(n12075), .op(
        n11039) );
  and3_1 U10176 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip3(n11039), .op(n8462) );
  inv_1 U10177 ( .ip(n9827), .op(n12336) );
  inv_1 U10178 ( .ip(n10975), .op(n8549) );
  or2_1 U10179 ( .ip1(n12336), .ip2(n8549), .op(n8454) );
  nand2_1 U10180 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n11754), .op(
        n12071) );
  or2_1 U10181 ( .ip1(n12071), .ip2(n8549), .op(n8453) );
  nand2_1 U10182 ( .ip1(n8454), .ip2(n8453), .op(n8461) );
  nor2_1 U10183 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n12352), .op(
        n11175) );
  nand2_1 U10184 ( .ip1(n11175), .ip2(n11089), .op(n8496) );
  inv_1 U10185 ( .ip(n12621), .op(n8455) );
  nand2_1 U10186 ( .ip1(n8456), .ip2(n8455), .op(n8458) );
  nand2_1 U10187 ( .ip1(n8458), .ip2(n8457), .op(n8459) );
  nand2_1 U10188 ( .ip1(n8459), .ip2(n11038), .op(n8460) );
  nand2_1 U10189 ( .ip1(n8496), .ip2(n8460), .op(n12083) );
  nor4_1 U10190 ( .ip1(n10810), .ip2(n8462), .ip3(n8461), .ip4(n12083), .op(
        n8470) );
  inv_1 U10191 ( .ip(n11206), .op(n8463) );
  nor3_1 U10192 ( .ip1(n10908), .ip2(n9620), .ip3(n8463), .op(n8492) );
  inv_1 U10193 ( .ip(\CORTEXM0DS_INST/u_logic/D69vx4 ), .op(n12558) );
  nor3_1 U10194 ( .ip1(\CORTEXM0DS_INST/u_logic/R89vx4 ), .ip2(n12564), .ip3(
        n12558), .op(n8487) );
  nor2_1 U10195 ( .ip1(n8487), .ip2(n12584), .op(n10870) );
  nor2_1 U10196 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Mc9vx4 ), .op(n9692) );
  nor4_1 U10197 ( .ip1(n10870), .ip2(n9692), .ip3(n10869), .ip4(n12073), .op(
        n8468) );
  nand2_1 U10198 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Ho8vx4 ), .op(n5100) );
  or2_1 U10199 ( .ip1(n5100), .ip2(n12075), .op(n8465) );
  or2_1 U10200 ( .ip1(n12332), .ip2(n12075), .op(n8464) );
  nand2_1 U10201 ( .ip1(n8465), .ip2(n8464), .op(n8467) );
  nor4_1 U10202 ( .ip1(n8492), .ip2(n8468), .ip3(n8467), .ip4(n8466), .op(
        n8469) );
  nand4_1 U10203 ( .ip1(n8472), .ip2(n8471), .ip3(n8470), .ip4(n8469), .op(
        n1744) );
  nor2_1 U10204 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n8738), .op(
        n11074) );
  inv_1 U10205 ( .ip(n8554), .op(n8473) );
  nand2_1 U10206 ( .ip1(n8474), .ip2(n8473), .op(n8483) );
  nand2_1 U10207 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n12584), .op(
        n10758) );
  nor2_1 U10208 ( .ip1(n12592), .ip2(n10749), .op(n10828) );
  nand2_1 U10209 ( .ip1(n10828), .ip2(n12338), .op(n11070) );
  not_ab_or_c_or_d U10210 ( .ip1(n12075), .ip2(n10758), .ip3(n10782), .ip4(
        n11070), .op(n8482) );
  inv_1 U10211 ( .ip(n10899), .op(n8475) );
  or2_1 U10212 ( .ip1(n8475), .ip2(n9620), .op(n8478) );
  inv_1 U10213 ( .ip(n9757), .op(n8476) );
  or2_1 U10214 ( .ip1(n8476), .ip2(n9620), .op(n8477) );
  nand2_1 U10215 ( .ip1(n8478), .ip2(n8477), .op(n8480) );
  nand2_1 U10216 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n10726), .op(
        n9832) );
  nor2_1 U10217 ( .ip1(n10771), .ip2(n9832), .op(n8479) );
  or2_1 U10218 ( .ip1(n10027), .ip2(n8479), .op(n8557) );
  ab_or_c_or_d U10219 ( .ip1(n11175), .ip2(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), 
        .ip3(n8480), .ip4(n8557), .op(n8481) );
  not_ab_or_c_or_d U10220 ( .ip1(n11074), .ip2(n8483), .ip3(n8482), .ip4(n8481), .op(n8498) );
  nor2_1 U10221 ( .ip1(n12075), .ip2(n10782), .op(n10462) );
  nand2_1 U10222 ( .ip1(n10462), .ip2(n12280), .op(n8486) );
  nand3_1 U10223 ( .ip1(\CORTEXM0DS_INST/u_logic/P39vx4 ), .ip2(n11756), .ip3(
        n12625), .op(n8485) );
  nand3_1 U10224 ( .ip1(n9753), .ip2(n10727), .ip3(n12095), .op(n8484) );
  nand3_1 U10225 ( .ip1(n8486), .ip2(n8485), .ip3(n8484), .op(n8494) );
  nand2_1 U10226 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Cf9vx4 ), .op(n8809) );
  nor4_1 U10227 ( .ip1(n12584), .ip2(n8809), .ip3(n10652), .ip4(n10605), .op(
        n11054) );
  nor2_1 U10228 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n10925), .op(
        n10766) );
  inv_1 U10229 ( .ip(n10766), .op(n10746) );
  nand2_1 U10230 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Cf9vx4 ), .op(n11139) );
  inv_1 U10231 ( .ip(n10605), .op(n11068) );
  nand2_1 U10232 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n12338), .op(
        n12330) );
  nor2_1 U10233 ( .ip1(n12329), .ip2(n12330), .op(n11052) );
  nand2_1 U10234 ( .ip1(n11068), .ip2(n11052), .op(n10813) );
  inv_1 U10235 ( .ip(n10813), .op(n12381) );
  nand2_1 U10236 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(n12381), .op(
        n12359) );
  nor4_1 U10237 ( .ip1(\CORTEXM0DS_INST/u_logic/D69vx4 ), .ip2(n10746), .ip3(
        n11139), .ip4(n12359), .op(n8488) );
  or2_1 U10238 ( .ip1(n11054), .ip2(n8488), .op(n8490) );
  nor2_1 U10239 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n12580), .op(
        n10756) );
  nand2_1 U10240 ( .ip1(n8487), .ip2(n10756), .op(n10700) );
  inv_1 U10241 ( .ip(n10700), .op(n9698) );
  or2_1 U10242 ( .ip1(n9698), .ip2(n8488), .op(n8489) );
  nand2_1 U10243 ( .ip1(n8490), .ip2(n8489), .op(n8491) );
  nor2_1 U10244 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n8491), .op(
        n8493) );
  not_ab_or_c_or_d U10245 ( .ip1(n12338), .ip2(n8494), .ip3(n8493), .ip4(n8492), .op(n8497) );
  nand2_1 U10246 ( .ip1(n8495), .ip2(n12034), .op(n10719) );
  nand4_1 U10247 ( .ip1(n8498), .ip2(n8497), .ip3(n10719), .ip4(n8496), .op(
        n3317) );
  inv_1 U10248 ( .ip(\CORTEXM0DS_INST/cm0_xpsr[24] ), .op(n12284) );
  nor3_1 U10249 ( .ip1(\CORTEXM0DS_INST/u_logic/H0gvx4 ), .ip2(n12284), .ip3(
        n12602), .op(n8759) );
  inv_1 U10250 ( .ip(n8759), .op(n12657) );
  nor2_1 U10251 ( .ip1(n12657), .ip2(n8499), .op(n4815) );
  inv_1 U10252 ( .ip(n4815), .op(n12527) );
  inv_1 U10253 ( .ip(n12639), .op(n12090) );
  inv_1 U10254 ( .ip(n1186), .op(n12528) );
  nand3_1 U10255 ( .ip1(n12090), .ip2(n8500), .ip3(n12528), .op(n8502) );
  not_ab_or_c_or_d U10256 ( .ip1(n1709), .ip2(n8502), .ip3(n12641), .ip4(n8501), .op(n12593) );
  inv_1 U10257 ( .ip(n12593), .op(n12574) );
  nor4_1 U10258 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n8537), .ip3(
        n12527), .ip4(n12574), .op(n1144) );
  inv_1 U10259 ( .ip(n1144), .op(n12575) );
  nor2_1 U10260 ( .ip1(n1155), .ip2(n12575), .op(n8504) );
  or2_1 U10261 ( .ip1(\CORTEXM0DS_INST/u_logic/Bwfvx4 ), .ip2(n8504), .op(
        n8506) );
  or2_1 U10262 ( .ip1(\CORTEXM0DS_INST/u_logic/V8evx4 ), .ip2(n8537), .op(
        n8503) );
  not_ab_or_c_or_d U10263 ( .ip1(n12090), .ip2(n8503), .ip3(
        \CORTEXM0DS_INST/u_logic/Xyfvx4 ), .ip4(n12574), .op(n12597) );
  or2_1 U10264 ( .ip1(n12597), .ip2(n8504), .op(n8505) );
  nand2_1 U10265 ( .ip1(n8506), .ip2(n8505), .op(n8509) );
  nand2_1 U10266 ( .ip1(n12593), .ip2(\CORTEXM0DS_INST/u_logic/V8evx4 ), .op(
        n12568) );
  inv_1 U10267 ( .ip(n12568), .op(n12594) );
  nand2_1 U10268 ( .ip1(\CORTEXM0DS_INST/u_logic/G8fvx4 ), .ip2(n12594), .op(
        n8508) );
  nand2_1 U10269 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(n12574), .op(
        n8507) );
  nand4_1 U10270 ( .ip1(n1154), .ip2(n8509), .ip3(n8508), .ip4(n8507), .op(
        n6031) );
  nor2_1 U10271 ( .ip1(n1157), .ip2(n12575), .op(n8510) );
  or2_1 U10272 ( .ip1(\CORTEXM0DS_INST/u_logic/Qufvx4 ), .ip2(n8510), .op(
        n8512) );
  or2_1 U10273 ( .ip1(n12597), .ip2(n8510), .op(n8511) );
  nand2_1 U10274 ( .ip1(n8512), .ip2(n8511), .op(n8515) );
  nand2_1 U10275 ( .ip1(\CORTEXM0DS_INST/u_logic/V6fvx4 ), .ip2(n12594), .op(
        n8514) );
  nand2_1 U10276 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n12574), .op(
        n8513) );
  nand4_1 U10277 ( .ip1(n1076), .ip2(n8515), .ip3(n8514), .ip4(n8513), .op(
        n6016) );
  nand2_1 U10278 ( .ip1(\CORTEXM0DS_INST/u_logic/Ho8vx4 ), .ip2(n12574), .op(
        n8519) );
  nand3_1 U10279 ( .ip1(\CORTEXM0DS_INST/u_logic/Xyfvx4 ), .ip2(n12593), .ip3(
        n12657), .op(n8518) );
  nand2_1 U10280 ( .ip1(\CORTEXM0DS_INST/u_logic/R9fvx4 ), .ip2(n12594), .op(
        n8517) );
  nand2_1 U10281 ( .ip1(n12597), .ip2(\CORTEXM0DS_INST/u_logic/Mxfvx4 ), .op(
        n8516) );
  nand4_1 U10282 ( .ip1(n8519), .ip2(n8518), .ip3(n8517), .ip4(n8516), .op(
        \CORTEXM0DS_INST/u_logic/Llnvx4 ) );
  nand2_1 U10283 ( .ip1(\CORTEXM0DS_INST/vis_pc [2]), .ip2(n12321), .op(n8523)
         );
  nand2_1 U10284 ( .ip1(\CORTEXM0DS_INST/u_logic/O2dvx4 ), .ip2(n2120), .op(
        n8522) );
  nand2_1 U10285 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [3]), .ip2(n12320), .op(
        n8521) );
  or2_1 U10286 ( .ip1(n12317), .ip2(\CORTEXM0DS_INST/u_logic/Ekovx4 ), .op(
        n8520) );
  nand4_1 U10287 ( .ip1(n8523), .ip2(n8522), .ip3(n8521), .ip4(n8520), .op(
        n6091) );
  nand2_1 U10288 ( .ip1(\CORTEXM0DS_INST/vis_pc [8]), .ip2(n12321), .op(n8535)
         );
  nand2_1 U10289 ( .ip1(\CORTEXM0DS_INST/u_logic/Wadvx4 ), .ip2(n2120), .op(
        n8534) );
  nand2_1 U10290 ( .ip1(\CORTEXM0DS_INST/u_logic/Oy8vx4 ), .ip2(n12320), .op(
        n8533) );
  inv_1 U10291 ( .ip(n9055), .op(n8531) );
  inv_1 U10292 ( .ip(\CORTEXM0DS_INST/vis_pc [8]), .op(n8526) );
  inv_1 U10293 ( .ip(\CORTEXM0DS_INST/vis_pc [7]), .op(n12113) );
  nor2_1 U10294 ( .ip1(n12292), .ip2(n12113), .op(n12112) );
  inv_1 U10295 ( .ip(n12112), .op(n8525) );
  nand2_1 U10296 ( .ip1(\CORTEXM0DS_INST/vis_pc [8]), .ip2(n12112), .op(n12121) );
  inv_1 U10297 ( .ip(n12121), .op(n8524) );
  not_ab_or_c_or_d U10298 ( .ip1(n8526), .ip2(n8525), .ip3(n8524), .ip4(n12305), .op(n8530) );
  xor2_1 U10299 ( .ip1(n8528), .ip2(n8527), .op(n10012) );
  nor2_1 U10300 ( .ip1(n10012), .ip2(n12309), .op(n8529) );
  not_ab_or_c_or_d U10301 ( .ip1(n12314), .ip2(n8531), .ip3(n8530), .ip4(n8529), .op(\CORTEXM0DS_INST/u_logic/Xxovx4 ) );
  or2_1 U10302 ( .ip1(\CORTEXM0DS_INST/u_logic/Xxovx4 ), .ip2(n12317), .op(
        n8532) );
  nand4_1 U10303 ( .ip1(n8535), .ip2(n8534), .ip3(n8533), .ip4(n8532), .op(
        n6104) );
  buf_1 U10304 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12737) );
  buf_1 U10305 ( .ip(n12737), .op(n12730) );
  buf_1 U10306 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12725) );
  buf_1 U10307 ( .ip(n12725), .op(n12709) );
  buf_1 U10308 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12735) );
  buf_1 U10309 ( .ip(n12735), .op(n12728) );
  buf_1 U10310 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12733) );
  buf_1 U10311 ( .ip(n12733), .op(n12727) );
  buf_1 U10312 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12711) );
  buf_1 U10313 ( .ip(n12711), .op(n12704) );
  buf_1 U10314 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12717) );
  buf_1 U10315 ( .ip(n12717), .op(n12706) );
  buf_1 U10316 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12710) );
  buf_1 U10317 ( .ip(n12713), .op(n12707) );
  buf_1 U10318 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12724) );
  buf_1 U10319 ( .ip(n12724), .op(n12715) );
  buf_1 U10320 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12729) );
  buf_1 U10321 ( .ip(n12729), .op(n12721) );
  buf_1 U10322 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12720) );
  buf_1 U10323 ( .ip(n12720), .op(n12719) );
  buf_1 U10324 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12716) );
  buf_1 U10325 ( .ip(n12716), .op(n12712) );
  buf_1 U10326 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12732) );
  buf_1 U10327 ( .ip(n12732), .op(n12723) );
  buf_1 U10328 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12722) );
  buf_1 U10329 ( .ip(n12722), .op(n12714) );
  buf_1 U10330 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12726) );
  buf_1 U10331 ( .ip(n12726), .op(n12718) );
  buf_1 U10332 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12739) );
  buf_1 U10333 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12708) );
  buf_1 U10334 ( .ip(n12708), .op(n12699) );
  buf_1 U10335 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12713) );
  buf_1 U10336 ( .ip(n12713), .op(n12698) );
  buf_1 U10337 ( .ip(n12715), .op(n12734) );
  buf_1 U10338 ( .ip(n12715), .op(n12701) );
  buf_1 U10339 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12703) );
  buf_1 U10340 ( .ip(n12726), .op(n12702) );
  buf_1 U10341 ( .ip(\CORTEXM0DS_INST/u_logic/N586 ), .op(n12705) );
  buf_1 U10342 ( .ip(n12705), .op(n12731) );
  buf_1 U10343 ( .ip(n12736), .op(n12700) );
  inv_1 U10344 ( .ip(\CORTEXM0DS_INST/u_logic/Mf8vx4 ), .op(n12635) );
  nor2_1 U10345 ( .ip1(n8536), .ip2(n12635), .op(n12689) );
  buf_1 U10346 ( .ip(n12689), .op(n12695) );
  nor2_1 U10347 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n8537), .op(
        n8539) );
  nor4_1 U10348 ( .ip1(n8539), .ip2(n12527), .ip3(n8538), .ip4(n12574), .op(
        n1148) );
  nor2_1 U10349 ( .ip1(n12095), .ip2(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .op(
        n11660) );
  inv_1 U10350 ( .ip(n10816), .op(n10801) );
  nand4_1 U10351 ( .ip1(n12625), .ip2(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip3(
        n11660), .ip4(n10801), .op(n11862) );
  nor3_1 U10352 ( .ip1(n11863), .ip2(n11846), .ip3(n11862), .op(n8542) );
  nand3_1 U10353 ( .ip1(n11867), .ip2(n8540), .ip3(
        \CORTEXM0DS_INST/u_logic/Mf8vx4 ), .op(n11666) );
  inv_1 U10354 ( .ip(n11666), .op(n9716) );
  nor2_1 U10355 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [11]), .ip2(n9716), 
        .op(n8541) );
  nor4_1 U10356 ( .ip1(n8542), .ip2(n2531), .ip3(n12740), .ip4(n8541), .op(
        \CORTEXM0DS_INST/u_logic/Uzhvx4 ) );
  nor2_1 U10357 ( .ip1(n8543), .ip2(n11862), .op(n8545) );
  nor2_1 U10358 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [13]), .ip2(n9716), 
        .op(n8544) );
  nor4_1 U10359 ( .ip1(n8545), .ip2(n2502), .ip3(n12743), .ip4(n8544), .op(
        \CORTEXM0DS_INST/u_logic/Gzhvx4 ) );
  inv_1 U10360 ( .ip(n11862), .op(n12687) );
  and2_1 U10361 ( .ip1(n8546), .ip2(n12687), .op(n8548) );
  nor2_1 U10362 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [9]), .ip2(n9716), .op(
        n8547) );
  nor4_1 U10363 ( .ip1(n8548), .ip2(n2528), .ip3(n12741), .ip4(n8547), .op(
        \CORTEXM0DS_INST/u_logic/I0ivx4 ) );
  buf_1 U10364 ( .ip(n12699), .op(n12736) );
  buf_1 U10365 ( .ip(n12728), .op(n12738) );
  buf_1 U10366 ( .ip(n12727), .op(n12696) );
  buf_1 U10367 ( .ip(n12707), .op(n12697) );
  nand2_1 U10368 ( .ip1(n11661), .ip2(n10728), .op(n8550) );
  not_ab_or_c_or_d U10369 ( .ip1(n12096), .ip2(n8550), .ip3(n11751), .ip4(
        n8549), .op(n8558) );
  nand3_1 U10370 ( .ip1(n12686), .ip2(n9757), .ip3(n11725), .op(n8552) );
  nor2_1 U10371 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(n11211), .op(
        n10881) );
  nand2_1 U10372 ( .ip1(n10881), .ip2(n11169), .op(n8551) );
  nand2_1 U10373 ( .ip1(n8552), .ip2(n8551), .op(n9836) );
  nor2_1 U10374 ( .ip1(n8553), .ip2(n11183), .op(n8820) );
  nand3_1 U10375 ( .ip1(n8820), .ip2(n10728), .ip3(n8554), .op(n8555) );
  nand3_1 U10376 ( .ip1(n11184), .ip2(n8554), .ip3(n10865), .op(n10500) );
  nand2_1 U10377 ( .ip1(n8555), .ip2(n10500), .op(n8556) );
  nand2_1 U10378 ( .ip1(n11609), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [8]), 
        .op(n8562) );
  nand2_1 U10379 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [8]), .ip2(n11787), 
        .op(n8561) );
  nand2_1 U10380 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [8]), .ip2(n10265), 
        .op(n8560) );
  nand2_1 U10381 ( .ip1(n11610), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [8]), 
        .op(n8559) );
  nand4_1 U10382 ( .ip1(n8562), .ip2(n8561), .ip3(n8560), .ip4(n8559), .op(
        n3977) );
  inv_1 U10383 ( .ip(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .op(n12402) );
  nor2_1 U10384 ( .ip1(n9813), .ip2(n12402), .op(n12679) );
  inv_1 U10385 ( .ip(n11009), .op(n11464) );
  and2_1 U10386 ( .ip1(n8564), .ip2(n9813), .op(
        \CORTEXM0DS_INST/u_logic/Oq42z4 ) );
  nand2_1 U10387 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Oq42z4 ), .op(n9862) );
  nor2_1 U10388 ( .ip1(n11269), .ip2(n9862), .op(n8566) );
  nor3_1 U10389 ( .ip1(n8564), .ip2(n8563), .ip3(n12402), .op(n9863) );
  nand2_1 U10390 ( .ip1(n9863), .ip2(n12671), .op(n5996) );
  inv_1 U10391 ( .ip(n5996), .op(n8565) );
  not_ab_or_c_or_d U10392 ( .ip1(n12679), .ip2(n11464), .ip3(n8566), .ip4(
        n8565), .op(\CORTEXM0DS_INST/u_logic/Sx3wx4 ) );
  mux2_1 U10393 ( .ip1(n8598), .ip2(n11308), .s(n12679), .op(
        \CORTEXM0DS_INST/u_logic/O24wx4 ) );
  nand4_1 U10394 ( .ip1(n3227), .ip2(n3226), .ip3(n3229), .ip4(n3228), .op(
        n3230) );
  nand2_1 U10395 ( .ip1(\CORTEXM0DS_INST/u_logic/H3evx4 ), .ip2(n2120), .op(
        n8569) );
  nand2_1 U10396 ( .ip1(\CORTEXM0DS_INST/vis_pc [28]), .ip2(n12321), .op(n8568) );
  nand2_1 U10397 ( .ip1(\CORTEXM0DS_INST/vis_apsr [1]), .ip2(n12320), .op(
        n8567) );
  nand4_1 U10398 ( .ip1(n1813), .ip2(n8569), .ip3(n8568), .ip4(n8567), .op(
        n6078) );
  nand2_1 U10399 ( .ip1(\CORTEXM0DS_INST/u_logic/S4evx4 ), .ip2(n2120), .op(
        n8572) );
  nand2_1 U10400 ( .ip1(\CORTEXM0DS_INST/vis_pc [29]), .ip2(n12321), .op(n8571) );
  nand2_1 U10401 ( .ip1(\CORTEXM0DS_INST/vis_apsr [2]), .ip2(n12320), .op(
        n8570) );
  nand4_1 U10402 ( .ip1(n1870), .ip2(n8572), .ip3(n8571), .ip4(n8570), .op(
        n6084) );
  nand2_1 U10403 ( .ip1(\CORTEXM0DS_INST/u_logic/D6evx4 ), .ip2(n2120), .op(
        n8575) );
  nand2_1 U10404 ( .ip1(\CORTEXM0DS_INST/vis_pc [30]), .ip2(n12321), .op(n8574) );
  nand2_1 U10405 ( .ip1(\CORTEXM0DS_INST/vis_apsr [3]), .ip2(n12320), .op(
        n8573) );
  nand4_1 U10406 ( .ip1(n2122), .ip2(n8575), .ip3(n8574), .ip4(n8573), .op(
        n6108) );
  not_ab_or_c_or_d U10407 ( .ip1(\CORTEXM0DS_INST/u_logic/Uth2z4 [0]), .ip2(
        n11851), .ip3(n8577), .ip4(n8576), .op(n8580) );
  nor2_1 U10408 ( .ip1(n8578), .ip2(n9910), .op(n8579) );
  not_ab_or_c_or_d U10409 ( .ip1(n9910), .ip2(n8581), .ip3(n8580), .ip4(n8579), 
        .op(n8591) );
  inv_1 U10410 ( .ip(n8582), .op(n8584) );
  mux2_1 U10411 ( .ip1(n8584), .ip2(n8583), .s(n9910), .op(n8590) );
  inv_1 U10412 ( .ip(n8585), .op(n8587) );
  nor2_1 U10413 ( .ip1(n8590), .ip2(n8591), .op(n8586) );
  nor2_1 U10414 ( .ip1(n8587), .ip2(n8586), .op(n8589) );
  ab_or_c_or_d U10415 ( .ip1(n8591), .ip2(n8590), .ip3(n8589), .ip4(n8588), 
        .op(n8592) );
  nand3_1 U10416 ( .ip1(n9879), .ip2(n8592), .ip3(n12646), .op(n8597) );
  or2_1 U10417 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [0]), .ip2(n12646), .op(n8594)
         );
  or2_1 U10418 ( .ip1(\CORTEXM0DS_INST/u_logic/Eqgvx4 ), .ip2(n12646), .op(
        n8593) );
  nand2_1 U10419 ( .ip1(n8594), .ip2(n8593), .op(n8595) );
  or2_1 U10420 ( .ip1(n8596), .ip2(n8595), .op(n8635) );
  nand2_1 U10421 ( .ip1(n8597), .ip2(n8635), .op(n5664) );
  nand4_1 U10422 ( .ip1(\CORTEXM0DS_INST/u_logic/I4gvx4 ), .ip2(n12090), .ip3(
        n11038), .ip4(n12528), .op(n10989) );
  nand3_1 U10423 ( .ip1(n10915), .ip2(n10713), .ip3(
        \CORTEXM0DS_INST/u_logic/Fs8vx4 ), .op(n8603) );
  inv_1 U10424 ( .ip(n8598), .op(n11472) );
  nor2_1 U10425 ( .ip1(n10588), .ip2(n10646), .op(n8599) );
  or2_1 U10426 ( .ip1(n12034), .ip2(n8599), .op(n8601) );
  or2_1 U10427 ( .ip1(n11207), .ip2(n8599), .op(n8600) );
  nand2_1 U10428 ( .ip1(n8601), .ip2(n8600), .op(n8629) );
  inv_1 U10429 ( .ip(n8629), .op(n11768) );
  nand2_1 U10430 ( .ip1(n11472), .ip2(n11768), .op(n8602) );
  nand2_1 U10431 ( .ip1(n8603), .ip2(n8602), .op(n8633) );
  nand2_1 U10432 ( .ip1(n11730), .ip2(n10949), .op(n8825) );
  inv_1 U10433 ( .ip(n8825), .op(n12094) );
  nand2_1 U10434 ( .ip1(n12094), .ip2(n9597), .op(n9531) );
  inv_1 U10435 ( .ip(n9531), .op(n8608) );
  nor3_1 U10436 ( .ip1(n12095), .ip2(n10865), .ip3(n9934), .op(n8607) );
  nor2_1 U10437 ( .ip1(n12613), .ip2(n8831), .op(n11659) );
  nor2_1 U10438 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n12618), .op(
        n12605) );
  not_ab_or_c_or_d U10439 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(
        n12651), .ip3(n11182), .ip4(n11715), .op(n8604) );
  nor2_1 U10440 ( .ip1(n12605), .ip2(n8604), .op(n8605) );
  nor2_1 U10441 ( .ip1(n11038), .ip2(n8605), .op(n8606) );
  nor4_1 U10442 ( .ip1(n8608), .ip2(n8607), .ip3(n11659), .ip4(n8606), .op(
        n11238) );
  nor2_1 U10443 ( .ip1(n11238), .ip2(n12365), .op(n8627) );
  or2_1 U10444 ( .ip1(n8831), .ip2(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .op(
        n8613) );
  or2_1 U10445 ( .ip1(n8609), .ip2(n12095), .op(n8610) );
  nand2_1 U10446 ( .ip1(n10547), .ip2(n8610), .op(n8611) );
  or2_1 U10447 ( .ip1(n8611), .ip2(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .op(
        n8612) );
  nand2_1 U10448 ( .ip1(n8613), .ip2(n8612), .op(n8620) );
  nor4_1 U10449 ( .ip1(n9753), .ip2(n8614), .ip3(n10972), .ip4(n10865), .op(
        n8619) );
  nor3_1 U10450 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n10949), .ip3(
        n8823), .op(n8618) );
  inv_1 U10451 ( .ip(n10587), .op(n9612) );
  inv_1 U10452 ( .ip(n8986), .op(n10939) );
  nand2_1 U10453 ( .ip1(n9612), .ip2(n10939), .op(n8615) );
  nand4_1 U10454 ( .ip1(n8616), .ip2(n11191), .ip3(n8615), .ip4(n11213), .op(
        n8617) );
  nor4_1 U10455 ( .ip1(n8620), .ip2(n8619), .ip3(n8618), .ip4(n8617), .op(
        n11237) );
  nor2_1 U10456 ( .ip1(n11237), .ip2(n8745), .op(n8626) );
  nor2_1 U10457 ( .ip1(n12095), .ip2(n12352), .op(n12626) );
  nor4_1 U10458 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip3(n11164), .ip4(n12608), .op(
        n8621) );
  not_ab_or_c_or_d U10459 ( .ip1(n8622), .ip2(n10899), .ip3(n12626), .ip4(
        n8621), .op(n11239) );
  nor2_1 U10460 ( .ip1(n11239), .ip2(n8666), .op(n8625) );
  nand3_1 U10461 ( .ip1(n11038), .ip2(n9869), .ip3(
        \CORTEXM0DS_INST/u_logic/Efgvx4 ), .op(n8624) );
  nand2_1 U10462 ( .ip1(n8624), .ip2(n8623), .op(n11236) );
  nor4_1 U10463 ( .ip1(n8627), .ip2(n8626), .ip3(n8625), .ip4(n11236), .op(
        n11556) );
  inv_1 U10464 ( .ip(n10881), .op(n8628) );
  nor4_1 U10465 ( .ip1(n11556), .ip2(n10865), .ip3(n12095), .ip4(n8628), .op(
        n8631) );
  nor2_1 U10466 ( .ip1(n8629), .ip2(n11479), .op(n8630) );
  nor2_1 U10467 ( .ip1(n8631), .ip2(n8630), .op(n8632) );
  mux2_1 U10468 ( .ip1(n8633), .ip2(\CORTEXM0DS_INST/cm0_primask[0] ), .s(
        n8632), .op(n12429) );
  inv_1 U10469 ( .ip(n5664), .op(n8634) );
  or2_1 U10470 ( .ip1(n12429), .ip2(n8634), .op(n8636) );
  nand2_1 U10471 ( .ip1(n8636), .ip2(n8635), .op(n12472) );
  inv_1 U10472 ( .ip(n12472), .op(n12026) );
  inv_1 U10473 ( .ip(\CORTEXM0DS_INST/u_logic/Xlevx4 ), .op(n12446) );
  nand2_1 U10474 ( .ip1(n12026), .ip2(n12446), .op(n8760) );
  or2_1 U10475 ( .ip1(n10989), .ip2(n8760), .op(n8639) );
  nand3_1 U10476 ( .ip1(n12090), .ip2(\CORTEXM0DS_INST/u_logic/V8evx4 ), .ip3(
        n12574), .op(n8637) );
  or2_1 U10477 ( .ip1(n8637), .ip2(n8760), .op(n8638) );
  nand2_1 U10478 ( .ip1(n8639), .ip2(n8638), .op(n6048) );
  inv_1 U10479 ( .ip(n10828), .op(n11028) );
  nor2_1 U10480 ( .ip1(n12570), .ip2(n11028), .op(n8664) );
  or2_1 U10481 ( .ip1(n10880), .ip2(n11736), .op(n8640) );
  nand2_1 U10482 ( .ip1(n8640), .ip2(n8738), .op(n12059) );
  inv_1 U10483 ( .ip(n12059), .op(n8641) );
  not_ab_or_c_or_d U10484 ( .ip1(n11052), .ip2(n8664), .ip3(n1770), .ip4(n8641), .op(n12384) );
  nand2_1 U10485 ( .ip1(\CORTEXM0DS_INST/u_logic/R89vx4 ), .ip2(n12381), .op(
        n8651) );
  inv_1 U10486 ( .ip(n5100), .op(n8642) );
  inv_1 U10487 ( .ip(n10830), .op(n10488) );
  nor2_1 U10488 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n10488), .op(
        n10807) );
  or2_1 U10489 ( .ip1(n8642), .ip2(n10807), .op(n8643) );
  nand2_1 U10490 ( .ip1(n8643), .ip2(n12338), .op(n12378) );
  inv_1 U10491 ( .ip(n8809), .op(n10457) );
  inv_1 U10492 ( .ip(n10749), .op(n12328) );
  inv_1 U10493 ( .ip(n10652), .op(n11032) );
  nand3_1 U10494 ( .ip1(n10457), .ip2(n12328), .ip3(n11032), .op(n8645) );
  nor2_1 U10495 ( .ip1(n10652), .ip2(n10605), .op(n9679) );
  nor2_1 U10496 ( .ip1(n12588), .ip2(n12327), .op(n9559) );
  inv_1 U10497 ( .ip(n9559), .op(n10917) );
  nand2_1 U10498 ( .ip1(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip2(n10917), .op(
        n8644) );
  nand2_1 U10499 ( .ip1(n9679), .ip2(n8644), .op(n12377) );
  nor2_1 U10500 ( .ip1(n12330), .ip2(n9695), .op(n11135) );
  nand2_1 U10501 ( .ip1(n9657), .ip2(n11135), .op(n12324) );
  nand4_1 U10502 ( .ip1(n12378), .ip2(n8645), .ip3(n12377), .ip4(n12324), .op(
        n12366) );
  nand2_1 U10503 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n12366), .op(
        n8650) );
  nor2_1 U10504 ( .ip1(n10757), .ip2(n12592), .op(n9629) );
  nor2_1 U10505 ( .ip1(n12580), .ip2(n12588), .op(n9535) );
  inv_1 U10506 ( .ip(n9535), .op(n9540) );
  and3_1 U10507 ( .ip1(n9679), .ip2(n9629), .ip3(n9540), .op(n8646) );
  or2_1 U10508 ( .ip1(n11135), .ip2(n8646), .op(n8648) );
  or2_1 U10509 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(n8646), .op(
        n8647) );
  nand2_1 U10510 ( .ip1(n8648), .ip2(n8647), .op(n12382) );
  inv_1 U10511 ( .ip(n9679), .op(n10033) );
  nand2_1 U10512 ( .ip1(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip2(n12584), .op(
        n10750) );
  or2_1 U10513 ( .ip1(n10033), .ip2(n10750), .op(n10926) );
  or2_1 U10514 ( .ip1(n10652), .ip2(n9695), .op(n11069) );
  inv_1 U10515 ( .ip(n9566), .op(n12337) );
  nand4_1 U10516 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n9657), .ip3(
        n12338), .ip4(n12337), .op(n9669) );
  nand4_1 U10517 ( .ip1(n12382), .ip2(n10926), .ip3(n11069), .ip4(n9669), .op(
        n12367) );
  nand2_1 U10518 ( .ip1(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), .ip2(n12367), .op(
        n8649) );
  and4_1 U10519 ( .ip1(n12384), .ip2(n8651), .ip3(n8650), .ip4(n8649), .op(
        n8652) );
  or2_1 U10520 ( .ip1(n1770), .ip2(n8652), .op(n8654) );
  or2_1 U10521 ( .ip1(n11159), .ip2(n8652), .op(n8653) );
  nand2_1 U10522 ( .ip1(n8654), .ip2(n8653), .op(n6073) );
  inv_1 U10523 ( .ip(n9826), .op(n1521) );
  inv_1 U10524 ( .ip(n11222), .op(n12033) );
  nor4_1 U10525 ( .ip1(n12033), .ip2(n10790), .ip3(n10810), .ip4(n3348), .op(
        n8680) );
  nand2_1 U10526 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n11068), .op(
        n8655) );
  nand2_1 U10527 ( .ip1(n10506), .ip2(n8655), .op(n8699) );
  nand2_1 U10528 ( .ip1(\CORTEXM0DS_INST/u_logic/W49vx4 ), .ip2(n8699), .op(
        n8662) );
  nand2_1 U10529 ( .ip1(n12376), .ip2(n12356), .op(n8657) );
  nand2_1 U10530 ( .ip1(n8657), .ip2(n8656), .op(n8658) );
  nand2_1 U10531 ( .ip1(n8658), .ip2(n10040), .op(n8659) );
  nand2_1 U10532 ( .ip1(n8659), .ip2(n10727), .op(n8661) );
  nor2_1 U10533 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n10605), .op(
        n10526) );
  nand2_1 U10534 ( .ip1(\CORTEXM0DS_INST/u_logic/B19vx4 ), .ip2(n10526), .op(
        n8660) );
  nand4_1 U10535 ( .ip1(n8680), .ip2(n8662), .ip3(n8661), .ip4(n8660), .op(
        n8663) );
  not_ab_or_c_or_d U10536 ( .ip1(n11650), .ip2(
        \CORTEXM0DS_INST/u_logic/Su9vx4 ), .ip3(n8664), .ip4(n8663), .op(n8665) );
  or2_1 U10537 ( .ip1(n3348), .ip2(n8665), .op(n8668) );
  or2_1 U10538 ( .ip1(n8666), .ip2(n8665), .op(n8667) );
  nand2_1 U10539 ( .ip1(n8668), .ip2(n8667), .op(
        \CORTEXM0DS_INST/u_logic/G2mvx4 ) );
  nor2_1 U10540 ( .ip1(n12564), .ip2(n11028), .op(n8685) );
  nor2_1 U10541 ( .ip1(n11159), .ip2(n12649), .op(n8683) );
  or2_1 U10542 ( .ip1(\CORTEXM0DS_INST/u_logic/Bx9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Su9vx4 ), .op(n8670) );
  or2_1 U10543 ( .ip1(n12356), .ip2(\CORTEXM0DS_INST/u_logic/Su9vx4 ), .op(
        n8669) );
  nand2_1 U10544 ( .ip1(n8670), .ip2(n8669), .op(n8671) );
  nor2_1 U10545 ( .ip1(\CORTEXM0DS_INST/u_logic/Ot9vx4 ), .ip2(n8671), .op(
        n8677) );
  or2_1 U10546 ( .ip1(\CORTEXM0DS_INST/u_logic/Ks9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Cq9vx4 ), .op(n8673) );
  or2_1 U10547 ( .ip1(n10038), .ip2(\CORTEXM0DS_INST/u_logic/Cq9vx4 ), .op(
        n8672) );
  nand2_1 U10548 ( .ip1(n8673), .ip2(n8672), .op(n8674) );
  nor2_1 U10549 ( .ip1(n8675), .ip2(n8674), .op(n8676) );
  nor2_1 U10550 ( .ip1(n8677), .ip2(n8676), .op(n8679) );
  nor2_1 U10551 ( .ip1(n8679), .ip2(n8678), .op(n8682) );
  inv_1 U10552 ( .ip(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), .op(n12535) );
  inv_1 U10553 ( .ip(n10526), .op(n9681) );
  nor2_1 U10554 ( .ip1(n12535), .ip2(n9681), .op(n8681) );
  nand2_1 U10555 ( .ip1(n8680), .ip2(n10488), .op(n8705) );
  or4_1 U10556 ( .ip1(n8683), .ip2(n8682), .ip3(n8681), .ip4(n8705), .op(n8684) );
  not_ab_or_c_or_d U10557 ( .ip1(\CORTEXM0DS_INST/u_logic/P39vx4 ), .ip2(n8699), .ip3(n8685), .ip4(n8684), .op(n8686) );
  or2_1 U10558 ( .ip1(n3348), .ip2(n8686), .op(n8688) );
  or2_1 U10559 ( .ip1(n11160), .ip2(n8686), .op(n8687) );
  nand2_1 U10560 ( .ip1(n8688), .ip2(n8687), .op(
        \CORTEXM0DS_INST/u_logic/Kuhvx4 ) );
  inv_1 U10561 ( .ip(\CORTEXM0DS_INST/u_logic/I29vx4 ), .op(n12544) );
  nor2_1 U10562 ( .ip1(n12544), .ip2(n9681), .op(n8689) );
  not_ab_or_c_or_d U10563 ( .ip1(\CORTEXM0DS_INST/u_logic/D69vx4 ), .ip2(n8699), .ip3(n8689), .ip4(n8705), .op(n8693) );
  nand2_1 U10564 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n10828), .op(
        n8692) );
  nand2_1 U10565 ( .ip1(n8698), .ip2(n10727), .op(n8691) );
  nand2_1 U10566 ( .ip1(\CORTEXM0DS_INST/u_logic/Wv9vx4 ), .ip2(n11650), .op(
        n8690) );
  and4_1 U10567 ( .ip1(n8693), .ip2(n8692), .ip3(n8691), .ip4(n8690), .op(
        n8694) );
  or2_1 U10568 ( .ip1(n3348), .ip2(n8694), .op(n8697) );
  or2_1 U10569 ( .ip1(n8695), .ip2(n8694), .op(n8696) );
  nand2_1 U10570 ( .ip1(n8697), .ip2(n8696), .op(
        \CORTEXM0DS_INST/u_logic/Pfhvx4 ) );
  nor2_1 U10571 ( .ip1(\CORTEXM0DS_INST/u_logic/Ks9vx4 ), .ip2(n10030), .op(
        n10898) );
  nand4_1 U10572 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip3(n8698), .ip4(n10727), .op(
        n8703) );
  nand3_1 U10573 ( .ip1(\CORTEXM0DS_INST/u_logic/K79vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip3(n8699), .op(n8702) );
  nand2_1 U10574 ( .ip1(\CORTEXM0DS_INST/u_logic/P39vx4 ), .ip2(n10526), .op(
        n8701) );
  nand2_1 U10575 ( .ip1(\CORTEXM0DS_INST/u_logic/Bx9vx4 ), .ip2(n11650), .op(
        n8700) );
  nand4_1 U10576 ( .ip1(n8703), .ip2(n8702), .ip3(n8701), .ip4(n8700), .op(
        n8704) );
  not_ab_or_c_or_d U10577 ( .ip1(n10727), .ip2(n10898), .ip3(n8705), .ip4(
        n8704), .op(n8706) );
  or2_1 U10578 ( .ip1(n3348), .ip2(n8706), .op(n8709) );
  or2_1 U10579 ( .ip1(n8707), .ip2(n8706), .op(n8708) );
  nand2_1 U10580 ( .ip1(n8709), .ip2(n8708), .op(
        \CORTEXM0DS_INST/u_logic/Ifhvx4 ) );
  nand3_1 U10581 ( .ip1(n9566), .ip2(n11725), .ip3(n11039), .op(n8730) );
  nor2_1 U10582 ( .ip1(n12584), .ip2(n8730), .op(n8710) );
  nor2_1 U10583 ( .ip1(n12034), .ip2(n8710), .op(n8711) );
  nor2_1 U10584 ( .ip1(n8711), .ip2(n12570), .op(n8718) );
  nor3_1 U10585 ( .ip1(n12075), .ip2(n8809), .ip3(n8738), .op(n8715) );
  nor2_1 U10586 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n10767), .op(
        n9552) );
  nor3_1 U10587 ( .ip1(n8712), .ip2(n9552), .ip3(n8730), .op(n8714) );
  inv_1 U10588 ( .ip(n12034), .op(n12333) );
  nor4_1 U10589 ( .ip1(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/B19vx4 ), .ip3(n12550), .ip4(n12333), .op(
        n8713) );
  nor4_1 U10590 ( .ip1(n3392), .ip2(n8715), .ip3(n8714), .ip4(n8713), .op(
        n8740) );
  nand2_1 U10591 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Kg9vx4 ), .op(n8716) );
  nand2_1 U10592 ( .ip1(n10457), .ip2(n8716), .op(n8727) );
  nand2_1 U10593 ( .ip1(n12034), .ip2(n12550), .op(n8729) );
  nand2_1 U10594 ( .ip1(n8738), .ip2(n8729), .op(n8717) );
  nand2_1 U10595 ( .ip1(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip2(n11033), .op(
        n8737) );
  nand4_1 U10596 ( .ip1(n8740), .ip2(n8727), .ip3(n8717), .ip4(n8737), .op(
        n8753) );
  nor2_1 U10597 ( .ip1(n8718), .ip2(n8753), .op(n8719) );
  or2_1 U10598 ( .ip1(n3392), .ip2(n8719), .op(n8722) );
  or2_1 U10599 ( .ip1(n8720), .ip2(n8719), .op(n8721) );
  nand2_1 U10600 ( .ip1(n8722), .ip2(n8721), .op(
        \CORTEXM0DS_INST/u_logic/Jxhvx4 ) );
  nand2_1 U10601 ( .ip1(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip2(n12329), .op(
        n10607) );
  not_ab_or_c_or_d U10602 ( .ip1(n12075), .ip2(n10607), .ip3(n11039), .ip4(
        n8738), .op(n8754) );
  nand2_1 U10603 ( .ip1(n12530), .ip2(n12075), .op(n8724) );
  nand2_1 U10604 ( .ip1(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip2(n10607), .op(
        n8723) );
  nand2_1 U10605 ( .ip1(n8724), .ip2(n8723), .op(n8725) );
  or2_1 U10606 ( .ip1(n8725), .ip2(n10617), .op(n8726) );
  nand2_1 U10607 ( .ip1(n8727), .ip2(n8726), .op(n8728) );
  nor2_1 U10608 ( .ip1(n8728), .ip2(n8738), .op(n8748) );
  nand2_1 U10609 ( .ip1(\CORTEXM0DS_INST/u_logic/P39vx4 ), .ip2(n8748), .op(
        n8732) );
  nand2_1 U10610 ( .ip1(n8730), .ip2(n8729), .op(n8749) );
  nand2_1 U10611 ( .ip1(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), .ip2(n8749), .op(
        n8731) );
  nand2_1 U10612 ( .ip1(n8732), .ip2(n8731), .op(n8733) );
  not_ab_or_c_or_d U10613 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n8754), .ip3(n8753), .ip4(n8733), .op(n8734) );
  or2_1 U10614 ( .ip1(n3392), .ip2(n8734), .op(n8736) );
  or2_1 U10615 ( .ip1(n11158), .ip2(n8734), .op(n8735) );
  nand2_1 U10616 ( .ip1(n8736), .ip2(n8735), .op(
        \CORTEXM0DS_INST/u_logic/Awhvx4 ) );
  nor3_1 U10617 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n8738), .ip3(
        n8737), .op(n8743) );
  nand2_1 U10618 ( .ip1(n8748), .ip2(\CORTEXM0DS_INST/u_logic/W49vx4 ), .op(
        n8741) );
  nand2_1 U10619 ( .ip1(\CORTEXM0DS_INST/u_logic/B19vx4 ), .ip2(n8749), .op(
        n8739) );
  nand3_1 U10620 ( .ip1(n8741), .ip2(n8740), .ip3(n8739), .op(n8742) );
  not_ab_or_c_or_d U10621 ( .ip1(n8754), .ip2(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip3(n8743), .ip4(n8742), .op(n8744) );
  or2_1 U10622 ( .ip1(n3392), .ip2(n8744), .op(n8747) );
  or2_1 U10623 ( .ip1(n8745), .ip2(n8744), .op(n8746) );
  nand2_1 U10624 ( .ip1(n8747), .ip2(n8746), .op(
        \CORTEXM0DS_INST/u_logic/Pthvx4 ) );
  nand2_1 U10625 ( .ip1(\CORTEXM0DS_INST/u_logic/D69vx4 ), .ip2(n8748), .op(
        n8751) );
  nand2_1 U10626 ( .ip1(\CORTEXM0DS_INST/u_logic/I29vx4 ), .ip2(n8749), .op(
        n8750) );
  nand2_1 U10627 ( .ip1(n8751), .ip2(n8750), .op(n8752) );
  not_ab_or_c_or_d U10628 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n8754), .ip3(n8753), .ip4(n8752), .op(n8755) );
  or2_1 U10629 ( .ip1(n3392), .ip2(n8755), .op(n8758) );
  or2_1 U10630 ( .ip1(n8756), .ip2(n8755), .op(n8757) );
  nand2_1 U10631 ( .ip1(n8758), .ip2(n8757), .op(
        \CORTEXM0DS_INST/u_logic/Rghvx4 ) );
  inv_1 U10632 ( .ip(n8760), .op(n12024) );
  nand2_1 U10633 ( .ip1(n12024), .ip2(n10989), .op(n4814) );
  nor2_1 U10634 ( .ip1(\CORTEXM0DS_INST/u_logic/R9fvx4 ), .ip2(n4814), .op(
        n8761) );
  or2_1 U10635 ( .ip1(n8759), .ip2(n8761), .op(n8763) );
  nor2_1 U10636 ( .ip1(n10989), .ip2(n8760), .op(n12430) );
  or2_1 U10637 ( .ip1(n12430), .ip2(n8761), .op(n8762) );
  nand2_1 U10638 ( .ip1(n8763), .ip2(n8762), .op(
        \CORTEXM0DS_INST/u_logic/Slnvx4 ) );
  nand2_1 U10639 ( .ip1(\CORTEXM0DS_INST/u_logic/N6hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Xahvx4 ), .op(n8764) );
  nand2_1 U10640 ( .ip1(n11867), .ip2(\CORTEXM0DS_INST/u_logic/Mf8vx4 ), .op(
        n12684) );
  nor2_1 U10641 ( .ip1(n8764), .ip2(n12684), .op(n12688) );
  nand2_1 U10642 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(n12681), .op(
        n6167) );
  inv_1 U10643 ( .ip(n12688), .op(n8766) );
  nor2_1 U10644 ( .ip1(n6167), .ip2(n11666), .op(n8765) );
  not_ab_or_c_or_d U10645 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [7]), .ip2(
        n8766), .ip3(n12751), .ip4(n8765), .op(n8767) );
  or2_1 U10646 ( .ip1(n12687), .ip2(n8767), .op(n8770) );
  or2_1 U10647 ( .ip1(n8768), .ip2(n8767), .op(n8769) );
  nand2_1 U10648 ( .ip1(n8770), .ip2(n8769), .op(
        \CORTEXM0DS_INST/u_logic/W0ivx4 ) );
  nand2_1 U10649 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(n12667), .op(
        n6172) );
  nor2_1 U10650 ( .ip1(n11666), .ip2(n6172), .op(n8771) );
  or2_1 U10651 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [2]), .ip2(n8771), .op(
        n8772) );
  nand2_1 U10652 ( .ip1(n2620), .ip2(n8772), .op(n8773) );
  or2_1 U10653 ( .ip1(n12687), .ip2(n8773), .op(n8776) );
  or2_1 U10654 ( .ip1(n8774), .ip2(n8773), .op(n8775) );
  nand2_1 U10655 ( .ip1(n8776), .ip2(n8775), .op(
        \CORTEXM0DS_INST/u_logic/F2ivx4 ) );
  nand2_1 U10656 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(n12671), .op(
        n6176) );
  nor2_1 U10657 ( .ip1(n11666), .ip2(n6176), .op(n8777) );
  or2_1 U10658 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [4]), .ip2(n8777), .op(
        n8778) );
  nand2_1 U10659 ( .ip1(n8778), .ip2(n2641), .op(n8779) );
  or2_1 U10660 ( .ip1(n12687), .ip2(n8779), .op(n8782) );
  or2_1 U10661 ( .ip1(n8780), .ip2(n8779), .op(n8781) );
  nand2_1 U10662 ( .ip1(n8782), .ip2(n8781), .op(
        \CORTEXM0DS_INST/u_logic/R1ivx4 ) );
  inv_1 U10663 ( .ip(n12677), .op(n9864) );
  mux2_1 U10664 ( .ip1(n11295), .ip2(n9864), .s(n9863), .op(
        \CORTEXM0DS_INST/u_logic/Bq5wx4 ) );
  nor2_1 U10665 ( .ip1(\CORTEXM0DS_INST/u_logic/Bq5wx4 ), .ip2(n11666), .op(
        n8783) );
  or2_1 U10666 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [14]), .ip2(n8783), .op(
        n8784) );
  nand2_1 U10667 ( .ip1(n8784), .ip2(n2754), .op(n8785) );
  or2_1 U10668 ( .ip1(n12687), .ip2(n8785), .op(n8788) );
  or2_1 U10669 ( .ip1(n8786), .ip2(n8785), .op(n8787) );
  nand2_1 U10670 ( .ip1(n8788), .ip2(n8787), .op(
        \CORTEXM0DS_INST/u_logic/Zyhvx4 ) );
  inv_1 U10671 ( .ip(n8789), .op(n12669) );
  nand2_1 U10672 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(n12669), .op(
        n6190) );
  nor2_1 U10673 ( .ip1(n11666), .ip2(n6190), .op(n8790) );
  or2_1 U10674 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [1]), .ip2(n8790), .op(
        n8791) );
  nand2_1 U10675 ( .ip1(n8791), .ip2(n2776), .op(n8792) );
  or2_1 U10676 ( .ip1(n12687), .ip2(n8792), .op(n8795) );
  or2_1 U10677 ( .ip1(n8793), .ip2(n8792), .op(n8794) );
  nand2_1 U10678 ( .ip1(n8795), .ip2(n8794), .op(
        \CORTEXM0DS_INST/u_logic/M2ivx4 ) );
  or2_1 U10679 ( .ip1(n12305), .ip2(n9826), .op(n8797) );
  nand2_1 U10680 ( .ip1(n8797), .ip2(n8796), .op(
        \CORTEXM0DS_INST/u_logic/N4421 ) );
  nor3_1 U10681 ( .ip1(\interconnect_ip_inst/i_ahb_U_mux_hsel_prev [1]), .ip2(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [2]), .ip3(
        \interconnect_ip_inst/i_ahb_U_dfltslv_current_state ), .op(n8799) );
  not_ab_or_c_or_d U10682 ( .ip1(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [2]), .ip2(
        \interconnect_ip_inst/i_apb_hready_resp ), .ip3(n8799), .ip4(n8798), 
        .op(\interconnect_ip_inst/n6491 ) );
  or2_1 U10683 ( .ip1(\interconnect_ip_inst/n6491 ), .ip2(n5926), .op(n8802)
         );
  or2_1 U10684 ( .ip1(n8800), .ip2(n5926), .op(n8801) );
  nand2_1 U10685 ( .ip1(n8802), .ip2(n8801), .op(\interconnect_ip_inst/n4861 )
         );
  nor2_1 U10686 ( .ip1(n8803), .ip2(n12635), .op(n12690) );
  and2_1 U10687 ( .ip1(n12430), .ip2(n4815), .op(n12692) );
  nor2_1 U10688 ( .ip1(n1186), .ip2(n12527), .op(n12693) );
  nand2_1 U10690 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(n12686), .op(
        n10927) );
  mux2_1 U10691 ( .ip1(n12564), .ip2(\CORTEXM0DS_INST/u_logic/K79vx4 ), .s(
        \CORTEXM0DS_INST/u_logic/D69vx4 ), .op(n11045) );
  nand4_1 U10692 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/R89vx4 ), .ip4(n11045), .op(n10616) );
  nor4_1 U10693 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n10707), .ip3(
        n10927), .ip4(n10616), .op(n8808) );
  nor4_1 U10694 ( .ip1(n9723), .ip2(n12095), .ip3(n12096), .ip4(n12613), .op(
        n8807) );
  or2_1 U10695 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n10874), .op(
        n8805) );
  or2_1 U10696 ( .ip1(n11184), .ip2(n10874), .op(n8804) );
  nand2_1 U10697 ( .ip1(n8805), .ip2(n8804), .op(n10471) );
  nor2_1 U10698 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Ki8vx4 ), .op(n9727) );
  nor3_1 U10699 ( .ip1(n10471), .ip2(n9727), .ip3(n12614), .op(n8806) );
  nand3_1 U10700 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n11184), .ip3(
        n11754), .op(n12631) );
  inv_1 U10701 ( .ip(n5938), .op(n12642) );
  nand3_1 U10702 ( .ip1(n12631), .ip2(n12642), .ip3(n10719), .op(n9665) );
  nor4_1 U10703 ( .ip1(n8808), .ip2(n8807), .ip3(n8806), .ip4(n9665), .op(
        n9580) );
  nor2_1 U10704 ( .ip1(n12075), .ip2(n8809), .op(n9659) );
  not_ab_or_c_or_d U10705 ( .ip1(n9659), .ip2(n8810), .ip3(n10970), .ip4(
        n11756), .op(n9579) );
  nand2_1 U10706 ( .ip1(n10975), .ip2(n9634), .op(n8815) );
  nand3_1 U10707 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip3(n9566), .op(n10685) );
  nor3_1 U10708 ( .ip1(\CORTEXM0DS_INST/u_logic/Ho8vx4 ), .ip2(n12075), .ip3(
        n10685), .op(n8812) );
  not_ab_or_c_or_d U10709 ( .ip1(n11661), .ip2(n11697), .ip3(n8812), .ip4(
        n8811), .op(n8814) );
  nand3_1 U10710 ( .ip1(n8815), .ip2(n8814), .ip3(n8813), .op(n9577) );
  nand3_1 U10711 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n12570), .ip3(
        n12564), .op(n8817) );
  nor2_1 U10712 ( .ip1(n9754), .ip2(\CORTEXM0DS_INST/u_logic/K79vx4 ), .op(
        n9741) );
  nor2_1 U10713 ( .ip1(n12570), .ip2(n9741), .op(n10505) );
  inv_1 U10714 ( .ip(n10505), .op(n8816) );
  nand2_1 U10715 ( .ip1(n8817), .ip2(n8816), .op(n8818) );
  nand2_1 U10716 ( .ip1(n9692), .ip2(n8818), .op(n10951) );
  inv_1 U10717 ( .ip(n10705), .op(n8994) );
  nor3_1 U10718 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip3(n8994), .op(n11180) );
  or2_1 U10719 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n11180), .op(
        n8830) );
  nand2_1 U10720 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n8819), .op(
        n11166) );
  nand2_1 U10721 ( .ip1(n8996), .ip2(n11166), .op(n8822) );
  nand2_1 U10722 ( .ip1(n10949), .ip2(n10539), .op(n9521) );
  inv_1 U10723 ( .ip(n9521), .op(n8821) );
  not_ab_or_c_or_d U10724 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n8822), .ip3(n8821), .ip4(n8820), .op(n8827) );
  nand2_1 U10725 ( .ip1(n11654), .ip2(n8823), .op(n8824) );
  nand2_1 U10726 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n8824), .op(
        n9524) );
  nand4_1 U10727 ( .ip1(n8827), .ip2(n9524), .ip3(n8826), .ip4(n8825), .op(
        n8828) );
  or2_1 U10728 ( .ip1(n8828), .ip2(n11180), .op(n8829) );
  nand2_1 U10729 ( .ip1(n8830), .ip2(n8829), .op(n11629) );
  nor3_1 U10730 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n12095), .ip3(
        n8831), .op(n10601) );
  nand2_1 U10731 ( .ip1(\CORTEXM0DS_INST/u_logic/O8gvx4 ), .ip2(n10601), .op(
        n11478) );
  nor3_1 U10732 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip3(n11478), .op(n11450) );
  nand2_1 U10733 ( .ip1(\CORTEXM0DS_INST/vis_apsr [3]), .ip2(n11450), .op(
        n9014) );
  and2_1 U10734 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [31]), .ip2(n8966), .op(n8840)
         );
  inv_1 U10735 ( .ip(\CORTEXM0DS_INST/u_logic/S4evx4 ), .op(n8879) );
  nor2_1 U10736 ( .ip1(n12051), .ip2(n8879), .op(n8834) );
  nor2_1 U10737 ( .ip1(n8832), .ip2(n8887), .op(n8833) );
  not_ab_or_c_or_d U10738 ( .ip1(\CORTEXM0DS_INST/vis_msp [29]), .ip2(n8949), 
        .ip3(n8834), .ip4(n8833), .op(n8838) );
  nand2_1 U10739 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [31]), .ip2(n8957), .op(n8837) );
  nand2_1 U10740 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [31]), .ip2(n8956), .op(n8836) );
  nand2_1 U10741 ( .ip1(\CORTEXM0DS_INST/u_logic/D6evx4 ), .ip2(n8947), .op(
        n8835) );
  not_ab_or_c_or_d U10742 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [31]), .ip2(n8944), 
        .ip3(n8840), .ip4(n8839), .op(n8844) );
  nand2_1 U10743 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [31]), .ip2(n8945), .op(n8843) );
  nand2_1 U10744 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [31]), .ip2(n8958), .op(n8842) );
  nand2_1 U10745 ( .ip1(\CORTEXM0DS_INST/vis_psp [29]), .ip2(n8959), .op(n8841) );
  nand2_1 U10746 ( .ip1(n9776), .ip2(n8969), .op(n9545) );
  nand2_1 U10747 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [31]), .op(n8847) );
  nand2_1 U10748 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [31]), .op(n8846) );
  nand2_1 U10749 ( .ip1(n8902), .ip2(\CORTEXM0DS_INST/cm0_r08 [31]), .op(n8845) );
  nand3_1 U10750 ( .ip1(n8847), .ip2(n8846), .ip3(n8845), .op(n8865) );
  and2_1 U10751 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [29]), .op(n8849)
         );
  and2_1 U10752 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [31]), .op(n8848)
         );
  not_ab_or_c_or_d U10753 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [31]), 
        .ip3(n8849), .ip4(n8848), .op(n8863) );
  nand2_1 U10754 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [31]), .op(n8852) );
  nand2_1 U10755 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [31]), .op(n8851) );
  nand2_1 U10756 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [31]), .op(n8850) );
  nand3_1 U10757 ( .ip1(n8852), .ip2(n8851), .ip3(n8850), .op(n8859) );
  nand2_1 U10758 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [31]), .op(n8857) );
  nand2_1 U10759 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [31]), .op(n8856) );
  nand2_1 U10760 ( .ip1(n8853), .ip2(\CORTEXM0DS_INST/u_logic/D6evx4 ), .op(
        n8855) );
  nand2_1 U10761 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [31]), .op(n8854) );
  not_ab_or_c_or_d U10762 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [31]), 
        .ip3(n8859), .ip4(n8858), .op(n8862) );
  nand2_1 U10763 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [29]), .op(n8861) );
  nand2_1 U10764 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [31]), .op(n8860) );
  not_ab_or_c_or_d U10765 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [31]), 
        .ip3(n8865), .ip4(n8864), .op(n11624) );
  mux2_1 U10766 ( .ip1(n8943), .ip2(n8942), .s(n11624), .op(n9544) );
  nand2_1 U10767 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [28]), .op(n8869) );
  nand2_1 U10768 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [28]), .op(n8868) );
  nand2_1 U10769 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [30]), .op(n8867) );
  nand2_1 U10770 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [30]), .op(n8866) );
  nand2_1 U10771 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [30]), .ip2(n8902), .op(n8884) );
  nand2_1 U10772 ( .ip1(n8910), .ip2(\CORTEXM0DS_INST/cm0_r14 [30]), .op(n8873) );
  nand2_1 U10773 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [30]), .op(n8872) );
  nand2_1 U10774 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [30]), .op(n8871) );
  nand2_1 U10775 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [30]), .op(n8870) );
  nand2_1 U10776 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [30]), .ip2(n8914), .op(n8876) );
  nand2_1 U10777 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [30]), .op(n8875) );
  nand2_1 U10778 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [30]), .op(n8874) );
  nand3_1 U10779 ( .ip1(n8876), .ip2(n8875), .ip3(n8874), .op(n8877) );
  not_ab_or_c_or_d U10780 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [30]), 
        .ip3(n8878), .ip4(n8877), .op(n8883) );
  and2_1 U10781 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [30]), .op(n8881)
         );
  nor2_1 U10782 ( .ip1(n8909), .ip2(n8879), .op(n8880) );
  not_ab_or_c_or_d U10783 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [30]), .ip2(n8917), 
        .ip3(n8881), .ip4(n8880), .op(n8882) );
  nand3_1 U10784 ( .ip1(n8884), .ip2(n8883), .ip3(n8882), .op(n8885) );
  not_ab_or_c_or_d U10785 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [30]), 
        .ip3(n8886), .ip4(n8885), .op(n11632) );
  mux2_1 U10786 ( .ip1(n8943), .ip2(n8942), .s(n11632), .op(n9123) );
  and2_1 U10787 ( .ip1(n8956), .ip2(\CORTEXM0DS_INST/cm0_r09 [30]), .op(n8896)
         );
  nor2_1 U10788 ( .ip1(n8888), .ip2(n8887), .op(n8890) );
  inv_1 U10789 ( .ip(\CORTEXM0DS_INST/u_logic/H3evx4 ), .op(n8908) );
  nor2_1 U10790 ( .ip1(n12051), .ip2(n8908), .op(n8889) );
  not_ab_or_c_or_d U10791 ( .ip1(\CORTEXM0DS_INST/u_logic/S4evx4 ), .ip2(n8947), .ip3(n8890), .ip4(n8889), .op(n8894) );
  nand2_1 U10792 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [30]), .op(n8893) );
  nand2_1 U10793 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [30]), .op(n8892) );
  nand2_1 U10794 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [28]), .op(n8891) );
  not_ab_or_c_or_d U10795 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [30]), .ip2(n8944), 
        .ip3(n8896), .ip4(n8895), .op(n8900) );
  nand2_1 U10796 ( .ip1(n8966), .ip2(\CORTEXM0DS_INST/cm0_r12 [30]), .op(n8899) );
  nand2_1 U10797 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [30]), .op(n8898) );
  nand2_1 U10798 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [28]), .op(n8897) );
  inv_1 U10799 ( .ip(n9122), .op(n9816) );
  nor2_1 U10800 ( .ip1(n9123), .ip2(n9816), .op(n11457) );
  nand2_1 U10801 ( .ip1(n8969), .ip2(n11457), .op(n8979) );
  nand2_1 U10802 ( .ip1(n9122), .ip2(n8969), .op(n8901) );
  xor2_1 U10803 ( .ip1(n9123), .ip2(n8901), .op(n8981) );
  nand2_1 U10804 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [29]), .ip2(n8902), .op(n8907) );
  nand2_1 U10805 ( .ip1(n8903), .ip2(\CORTEXM0DS_INST/cm0_r05 [29]), .op(n8906) );
  nand2_1 U10806 ( .ip1(n8904), .ip2(\CORTEXM0DS_INST/cm0_r04 [29]), .op(n8905) );
  nand3_1 U10807 ( .ip1(n8907), .ip2(n8906), .ip3(n8905), .op(n8940) );
  nor2_1 U10808 ( .ip1(n8909), .ip2(n8908), .op(n8911) );
  or2_1 U10809 ( .ip1(n8910), .ip2(n8911), .op(n8913) );
  or2_1 U10810 ( .ip1(\CORTEXM0DS_INST/cm0_r14 [29]), .ip2(n8911), .op(n8912)
         );
  nand2_1 U10811 ( .ip1(n8913), .ip2(n8912), .op(n8938) );
  nand2_1 U10812 ( .ip1(n8914), .ip2(\CORTEXM0DS_INST/cm0_r11 [29]), .op(n8921) );
  nand2_1 U10813 ( .ip1(n8915), .ip2(\CORTEXM0DS_INST/cm0_r03 [29]), .op(n8920) );
  nand2_1 U10814 ( .ip1(n8916), .ip2(\CORTEXM0DS_INST/cm0_r10 [29]), .op(n8919) );
  nand2_1 U10815 ( .ip1(n8917), .ip2(\CORTEXM0DS_INST/cm0_r01 [29]), .op(n8918) );
  nand2_1 U10816 ( .ip1(n8922), .ip2(\CORTEXM0DS_INST/vis_msp [27]), .op(n8929) );
  nand2_1 U10817 ( .ip1(n8923), .ip2(\CORTEXM0DS_INST/vis_psp [27]), .op(n8928) );
  nand2_1 U10818 ( .ip1(n8924), .ip2(\CORTEXM0DS_INST/cm0_r12 [29]), .op(n8927) );
  nand2_1 U10819 ( .ip1(n8925), .ip2(\CORTEXM0DS_INST/cm0_r06 [29]), .op(n8926) );
  not_ab_or_c_or_d U10820 ( .ip1(n8932), .ip2(\CORTEXM0DS_INST/cm0_r00 [29]), 
        .ip3(n8931), .ip4(n8930), .op(n8937) );
  nand2_1 U10821 ( .ip1(n8933), .ip2(\CORTEXM0DS_INST/cm0_r09 [29]), .op(n8936) );
  nand2_1 U10822 ( .ip1(n8934), .ip2(\CORTEXM0DS_INST/cm0_r07 [29]), .op(n8935) );
  not_ab_or_c_or_d U10823 ( .ip1(n8941), .ip2(\CORTEXM0DS_INST/cm0_r02 [29]), 
        .ip3(n8940), .ip4(n8939), .op(n11777) );
  mux2_1 U10824 ( .ip1(n8943), .ip2(n8942), .s(n11777), .op(n9186) );
  and2_1 U10825 ( .ip1(n8944), .ip2(\CORTEXM0DS_INST/cm0_r10 [29]), .op(n8965)
         );
  and2_1 U10826 ( .ip1(n8945), .ip2(\CORTEXM0DS_INST/cm0_r08 [29]), .op(n8955)
         );
  nand2_1 U10827 ( .ip1(n8946), .ip2(n9304), .op(n8953) );
  nand2_1 U10828 ( .ip1(n8947), .ip2(\CORTEXM0DS_INST/u_logic/H3evx4 ), .op(
        n8952) );
  nand2_1 U10829 ( .ip1(\CORTEXM0DS_INST/u_logic/W1evx4 ), .ip2(n8948), .op(
        n8951) );
  nand2_1 U10830 ( .ip1(n8949), .ip2(\CORTEXM0DS_INST/vis_msp [27]), .op(n8950) );
  not_ab_or_c_or_d U10831 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [29]), .ip2(n8956), 
        .ip3(n8955), .ip4(n8954), .op(n8963) );
  nand2_1 U10832 ( .ip1(n8957), .ip2(\CORTEXM0DS_INST/cm0_r11 [29]), .op(n8962) );
  nand2_1 U10833 ( .ip1(n8958), .ip2(\CORTEXM0DS_INST/cm0_r14 [29]), .op(n8961) );
  nand2_1 U10834 ( .ip1(n8959), .ip2(\CORTEXM0DS_INST/vis_psp [27]), .op(n8960) );
  not_ab_or_c_or_d U10835 ( .ip1(\CORTEXM0DS_INST/cm0_r12 [29]), .ip2(n8966), 
        .ip3(n8965), .ip4(n8964), .op(n9825) );
  nor2_1 U10836 ( .ip1(n9186), .ip2(n9825), .op(n8967) );
  nand2_1 U10837 ( .ip1(n8967), .ip2(n8969), .op(n8977) );
  or2_1 U10838 ( .ip1(n9160), .ip2(n9159), .op(n8968) );
  nand2_1 U10839 ( .ip1(n8969), .ip2(n8968), .op(n8973) );
  nor2_1 U10840 ( .ip1(n8971), .ip2(n8970), .op(n8972) );
  nor2_1 U10841 ( .ip1(n8973), .ip2(n8972), .op(n8985) );
  or2_1 U10842 ( .ip1(n9825), .ip2(n8974), .op(n8975) );
  xor2_1 U10843 ( .ip1(n9186), .ip2(n8975), .op(n8984) );
  nand2_1 U10844 ( .ip1(n8985), .ip2(n8984), .op(n8976) );
  nand2_1 U10845 ( .ip1(n8977), .ip2(n8976), .op(n8980) );
  nand2_1 U10846 ( .ip1(n8981), .ip2(n8980), .op(n8978) );
  and2_1 U10847 ( .ip1(n8979), .ip2(n8978), .op(n9513) );
  xor2_1 U10848 ( .ip1(n8981), .ip2(n8980), .op(n9249) );
  nor2_1 U10849 ( .ip1(n8983), .ip2(n8982), .op(n9237) );
  xor2_1 U10850 ( .ip1(n8985), .ip2(n8984), .op(n9236) );
  and2_1 U10851 ( .ip1(n9237), .ip2(n9236), .op(n9248) );
  nand2_1 U10852 ( .ip1(n9249), .ip2(n9248), .op(n9511) );
  xor2_1 U10853 ( .ip1(n9512), .ip2(n9511), .op(n10421) );
  nand3_1 U10854 ( .ip1(n10587), .ip2(n8987), .ip3(n8986), .op(n8989) );
  nor3_1 U10855 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n10865), .ip3(
        n6210), .op(n8988) );
  not_ab_or_c_or_d U10856 ( .ip1(n10865), .ip2(n8989), .ip3(n8988), .ip4(n9597), .op(n8990) );
  or2_1 U10857 ( .ip1(n8990), .ip2(n9582), .op(n8991) );
  nand2_1 U10858 ( .ip1(n8992), .ip2(n8991), .op(n11534) );
  nor3_1 U10859 ( .ip1(n8994), .ip2(n9582), .ip3(n8993), .op(n11538) );
  inv_1 U10860 ( .ip(n11538), .op(n11511) );
  or2_1 U10861 ( .ip1(n9544), .ip2(n11511), .op(n8995) );
  inv_1 U10862 ( .ip(n9776), .op(n9006) );
  nand2_1 U10863 ( .ip1(n8995), .ip2(n9006), .op(n9004) );
  not_ab_or_c_or_d U10864 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(
        n11164), .ip3(n12338), .ip4(n10770), .op(n8999) );
  nor3_1 U10865 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip3(n8996), .op(n8998) );
  nor3_1 U10866 ( .ip1(n11730), .ip2(n6210), .ip3(n10488), .op(n8997) );
  or4_1 U10867 ( .ip1(n10779), .ip2(n8999), .ip3(n8998), .ip4(n8997), .op(
        n9000) );
  nand2_1 U10868 ( .ip1(\CORTEXM0DS_INST/u_logic/O8gvx4 ), .ip2(n9000), .op(
        n9001) );
  nand2_1 U10869 ( .ip1(n9002), .ip2(n9001), .op(n9024) );
  nor2_1 U10870 ( .ip1(n11538), .ip2(n9024), .op(n11545) );
  nand2_1 U10871 ( .ip1(n9544), .ip2(n11545), .op(n9003) );
  nand2_1 U10872 ( .ip1(n9004), .ip2(n9003), .op(n9008) );
  nor2_1 U10873 ( .ip1(n11170), .ip2(n11186), .op(n9005) );
  not_ab_or_c_or_d U10874 ( .ip1(n11754), .ip2(n6210), .ip3(
        \CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip4(n9005), .op(n9025) );
  nor2_1 U10875 ( .ip1(n9024), .ip2(n9025), .op(n11434) );
  inv_1 U10876 ( .ip(n11434), .op(n11537) );
  nor3_1 U10877 ( .ip1(n9006), .ip2(n11537), .ip3(n9544), .op(n9007) );
  nor2_1 U10878 ( .ip1(n9008), .ip2(n9007), .op(n9012) );
  nand2_1 U10879 ( .ip1(n9009), .ip2(n11231), .op(n9010) );
  nand2_1 U10880 ( .ip1(\CORTEXM0DS_INST/u_logic/O8gvx4 ), .ip2(n9010), .op(
        n11331) );
  nor2_1 U10881 ( .ip1(n11624), .ip2(n11331), .op(n9011) );
  not_ab_or_c_or_d U10882 ( .ip1(n10421), .ip2(n11534), .ip3(n9012), .ip4(
        n9011), .op(n9013) );
  nor2_1 U10883 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n11754), .op(
        n11199) );
  nand3_1 U10884 ( .ip1(\CORTEXM0DS_INST/u_logic/O8gvx4 ), .ip2(n11199), .ip3(
        n12625), .op(n11451) );
  nand3_1 U10885 ( .ip1(n9014), .ip2(n9013), .ip3(n11451), .op(n11461) );
  nor2_1 U10886 ( .ip1(\CORTEXM0DS_INST/u_logic/Dw8vx4 ), .ip2(n11461), .op(
        n9536) );
  inv_1 U10887 ( .ip(n11534), .op(n11530) );
  xor2_1 U10888 ( .ip1(n9016), .ip2(n9015), .op(n12271) );
  nor2_1 U10889 ( .ip1(n11530), .ip2(n12271), .op(n11441) );
  xor2_1 U10890 ( .ip1(n9018), .ip2(n9017), .op(n12250) );
  nor2_1 U10891 ( .ip1(n11530), .ip2(n12250), .op(n11421) );
  xor2_1 U10892 ( .ip1(n9020), .ip2(n9019), .op(n12126) );
  inv_1 U10893 ( .ip(n11451), .op(n11548) );
  or2_1 U10894 ( .ip1(n12126), .ip2(n11548), .op(n9022) );
  or2_1 U10895 ( .ip1(n11534), .ip2(n11548), .op(n9021) );
  nand2_1 U10896 ( .ip1(n9022), .ip2(n9021), .op(n11259) );
  nor2_1 U10897 ( .ip1(n11530), .ip2(n10012), .op(n11155) );
  nor2_1 U10898 ( .ip1(n11511), .ip2(n9026), .op(n9023) );
  not_ab_or_c_or_d U10899 ( .ip1(n9025), .ip2(n9026), .ip3(n9024), .ip4(n9023), 
        .op(n9028) );
  nand2_1 U10900 ( .ip1(n11538), .ip2(n9026), .op(n9027) );
  mux2_1 U10901 ( .ip1(n9028), .ip2(n9027), .s(n12296), .op(n9033) );
  xor2_1 U10902 ( .ip1(n9030), .ip2(n9029), .op(n12299) );
  nand2_1 U10903 ( .ip1(n12299), .ip2(n11534), .op(n9032) );
  inv_1 U10904 ( .ip(n11331), .op(n11549) );
  nand2_1 U10905 ( .ip1(n11549), .ip2(n12681), .op(n9031) );
  nand4_1 U10906 ( .ip1(n9033), .ip2(n11451), .ip3(n9032), .ip4(n9031), .op(
        n11471) );
  nand2_1 U10907 ( .ip1(n11342), .ip2(n9141), .op(n9042) );
  nand2_1 U10908 ( .ip1(n12175), .ip2(n9132), .op(n11332) );
  nand2_1 U10909 ( .ip1(n12134), .ip2(n9145), .op(n11261) );
  nand2_1 U10910 ( .ip1(n9804), .ip2(n9137), .op(n11286) );
  nand3_1 U10911 ( .ip1(n11332), .ip2(n11261), .ip3(n11286), .op(n9039) );
  and2_1 U10912 ( .ip1(n9147), .ip2(n9810), .op(n11298) );
  nor2_1 U10913 ( .ip1(n11427), .ip2(n11431), .op(n9034) );
  not_ab_or_c_or_d U10914 ( .ip1(n12114), .ip2(n9136), .ip3(n11298), .ip4(
        n9034), .op(n9037) );
  and2_1 U10915 ( .ip1(n9139), .ip2(n9102), .op(n11379) );
  and2_1 U10916 ( .ip1(n9144), .ip2(n9097), .op(n11353) );
  not_ab_or_c_or_d U10917 ( .ip1(n11319), .ip2(n9140), .ip3(n11379), .ip4(
        n11353), .op(n9036) );
  nand2_1 U10918 ( .ip1(n12240), .ip2(n11406), .op(n11404) );
  nand2_1 U10919 ( .ip1(n10964), .ip2(n11540), .op(n9035) );
  nand4_1 U10920 ( .ip1(n9037), .ip2(n9036), .ip3(n11404), .ip4(n9035), .op(
        n9038) );
  not_ab_or_c_or_d U10921 ( .ip1(n12141), .ip2(n9143), .ip3(n9039), .ip4(n9038), .op(n9041) );
  and2_1 U10922 ( .ip1(n9100), .ip2(n9099), .op(n11422) );
  and2_1 U10923 ( .ip1(n9134), .ip2(n12159), .op(n11305) );
  not_ab_or_c_or_d U10924 ( .ip1(n11366), .ip2(n9142), .ip3(n11422), .ip4(
        n11305), .op(n9040) );
  nand3_1 U10925 ( .ip1(n9042), .ip2(n9041), .ip3(n9040), .op(n9088) );
  nand2_1 U10926 ( .ip1(n9047), .ip2(n11538), .op(n9043) );
  nand2_1 U10927 ( .ip1(n9043), .ip2(n9046), .op(n9045) );
  inv_1 U10928 ( .ip(n11545), .op(n11513) );
  or2_1 U10929 ( .ip1(n11513), .ip2(n9047), .op(n9044) );
  nand2_1 U10930 ( .ip1(n9045), .ip2(n9044), .op(n9049) );
  inv_1 U10931 ( .ip(n9046), .op(n12313) );
  and3_1 U10932 ( .ip1(n11434), .ip2(n12313), .ip3(n9047), .op(n9048) );
  nor2_1 U10933 ( .ip1(n9049), .ip2(n9048), .op(n11415) );
  nand2_1 U10934 ( .ip1(n11538), .ip2(n9050), .op(n9054) );
  nor2_1 U10935 ( .ip1(n11513), .ip2(n9050), .op(n9053) );
  nand2_1 U10936 ( .ip1(n11434), .ip2(n9050), .op(n9051) );
  nor2_1 U10937 ( .ip1(n9051), .ip2(n9055), .op(n9052) );
  not_ab_or_c_or_d U10938 ( .ip1(n9055), .ip2(n9054), .ip3(n9053), .ip4(n9052), 
        .op(n11154) );
  nand2_1 U10939 ( .ip1(n11538), .ip2(n9056), .op(n9060) );
  nor2_1 U10940 ( .ip1(n11513), .ip2(n9056), .op(n9059) );
  nand2_1 U10941 ( .ip1(n11434), .ip2(n9056), .op(n9057) );
  nor2_1 U10942 ( .ip1(n9057), .ip2(n12099), .op(n9058) );
  not_ab_or_c_or_d U10943 ( .ip1(n12099), .ip2(n9060), .ip3(n9059), .ip4(n9058), .op(n11529) );
  nand2_1 U10944 ( .ip1(n11538), .ip2(n9061), .op(n9065) );
  nor2_1 U10945 ( .ip1(n11513), .ip2(n9061), .op(n9064) );
  nand2_1 U10946 ( .ip1(n11434), .ip2(n9061), .op(n9062) );
  nor2_1 U10947 ( .ip1(n9062), .ip2(n12123), .op(n9063) );
  not_ab_or_c_or_d U10948 ( .ip1(n12123), .ip2(n9065), .ip3(n9064), .ip4(n9063), .op(n11257) );
  nand2_1 U10949 ( .ip1(n9066), .ip2(n11538), .op(n9067) );
  nand2_1 U10950 ( .ip1(n9067), .ip2(n9070), .op(n9069) );
  nand2_1 U10951 ( .ip1(n11545), .ip2(n9071), .op(n9068) );
  nand2_1 U10952 ( .ip1(n9069), .ip2(n9068), .op(n9073) );
  nor3_1 U10953 ( .ip1(n9071), .ip2(n11537), .ip3(n9070), .op(n9072) );
  nor2_1 U10954 ( .ip1(n9073), .ip2(n9072), .op(n11389) );
  nor4_1 U10955 ( .ip1(n11154), .ip2(n11529), .ip3(n11257), .ip4(n11389), .op(
        n9086) );
  nor2_1 U10956 ( .ip1(n9077), .ip2(n11511), .op(n9076) );
  or2_1 U10957 ( .ip1(n9077), .ip2(n11537), .op(n9075) );
  mux2_1 U10958 ( .ip1(n9076), .ip2(n9075), .s(n9074), .op(n9079) );
  nand2_1 U10959 ( .ip1(n11545), .ip2(n9077), .op(n9078) );
  nand2_1 U10960 ( .ip1(n9079), .ip2(n9078), .op(n11487) );
  inv_1 U10961 ( .ip(n9080), .op(n9083) );
  nor2_1 U10962 ( .ip1(n9083), .ip2(n11511), .op(n9082) );
  nand2_1 U10963 ( .ip1(n11434), .ip2(n9080), .op(n9081) );
  mux2_1 U10964 ( .ip1(n9082), .ip2(n9081), .s(n12233), .op(n9085) );
  nand2_1 U10965 ( .ip1(n11545), .ip2(n9083), .op(n9084) );
  nand2_1 U10966 ( .ip1(n9085), .ip2(n9084), .op(n11401) );
  nand3_1 U10967 ( .ip1(n9086), .ip2(n11487), .ip3(n11401), .op(n9087) );
  not_ab_or_c_or_d U10968 ( .ip1(n11538), .ip2(n9088), .ip3(n11415), .ip4(
        n9087), .op(n9129) );
  nor3_1 U10969 ( .ip1(n11545), .ip2(n12159), .ip3(n9134), .op(n11311) );
  nor3_1 U10970 ( .ip1(n11545), .ip2(n12134), .ip3(n9145), .op(n11263) );
  nor3_1 U10971 ( .ip1(n11545), .ip2(n9810), .ip3(n9147), .op(n11297) );
  nor3_1 U10972 ( .ip1(n11545), .ip2(n9804), .ip3(n9137), .op(n11288) );
  nor4_1 U10973 ( .ip1(n11311), .ip2(n11263), .ip3(n11297), .ip4(n11288), .op(
        n9128) );
  nor2_1 U10974 ( .ip1(n10964), .ip2(n11540), .op(n9092) );
  nor2_1 U10975 ( .ip1(n12114), .ip2(n9136), .op(n9091) );
  nor2_1 U10976 ( .ip1(n11342), .ip2(n9141), .op(n9090) );
  nor2_1 U10977 ( .ip1(n11366), .ip2(n9142), .op(n9089) );
  nor4_1 U10978 ( .ip1(n9092), .ip2(n9091), .ip3(n9090), .ip4(n9089), .op(
        n9096) );
  nor2_1 U10979 ( .ip1(n11319), .ip2(n9140), .op(n9094) );
  nor2_1 U10980 ( .ip1(n12141), .ip2(n9143), .op(n9093) );
  not_ab_or_c_or_d U10981 ( .ip1(n11427), .ip2(n11431), .ip3(n9094), .ip4(
        n9093), .op(n9095) );
  nand2_1 U10982 ( .ip1(n9096), .ip2(n9095), .op(n9101) );
  nor3_1 U10983 ( .ip1(n11545), .ip2(n9097), .ip3(n9144), .op(n11359) );
  nor2_1 U10984 ( .ip1(n11513), .ip2(n9100), .op(n9098) );
  not_ab_or_c_or_d U10985 ( .ip1(n11434), .ip2(n9100), .ip3(n9099), .ip4(n9098), .op(n11420) );
  not_ab_or_c_or_d U10986 ( .ip1(n11513), .ip2(n9101), .ip3(n11359), .ip4(
        n11420), .op(n9127) );
  nor3_1 U10987 ( .ip1(n11545), .ip2(n9102), .ip3(n9139), .op(n11384) );
  nor3_1 U10988 ( .ip1(n11545), .ip2(n12175), .ip3(n9132), .op(n11336) );
  nand2_1 U10989 ( .ip1(n11548), .ip2(\CORTEXM0DS_INST/cm0_control[1] ), .op(
        n9106) );
  nor2_1 U10990 ( .ip1(n12096), .ip2(n12625), .op(n10029) );
  nand4_1 U10991 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/O8gvx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Oy8vx4 ), .ip4(n10029), .op(n9105) );
  nor3_1 U10992 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(n11145), .ip3(
        n11478), .op(n11481) );
  nand2_1 U10993 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [2]), .ip2(n11481), .op(
        n9104) );
  nand2_1 U10994 ( .ip1(n10392), .ip2(n11534), .op(n9103) );
  nand4_1 U10995 ( .ip1(n9106), .ip2(n9105), .ip3(n9104), .ip4(n9103), .op(
        n11251) );
  and2_1 U10996 ( .ip1(n11481), .ip2(\CORTEXM0DS_INST/vis_ipsr [4]), .op(n9107) );
  not_ab_or_c_or_d U10997 ( .ip1(n11549), .ip2(n12671), .ip3(n11548), .ip4(
        n9107), .op(n11399) );
  inv_1 U10998 ( .ip(n11777), .op(n11447) );
  inv_1 U10999 ( .ip(n11632), .op(n11456) );
  nor4_1 U11000 ( .ip1(n11447), .ip2(n11456), .ip3(n11413), .ip4(n11423), .op(
        n9118) );
  inv_1 U11001 ( .ip(n9108), .op(n12672) );
  inv_1 U11002 ( .ip(n9109), .op(n12674) );
  nor4_1 U11003 ( .ip1(n12676), .ip2(n12672), .ip3(n12674), .ip4(n12673), .op(
        n9117) );
  nor4_1 U11004 ( .ip1(n11472), .ip2(n12669), .ip3(n12677), .ip4(n12678), .op(
        n9116) );
  nand4_1 U11005 ( .ip1(n11285), .ip2(n9858), .ip3(n11269), .ip4(n11260), .op(
        n9114) );
  inv_1 U11006 ( .ip(n12667), .op(n9110) );
  nand4_1 U11007 ( .ip1(n12666), .ip2(n11316), .ip3(n11356), .ip4(n9110), .op(
        n9113) );
  nand4_1 U11008 ( .ip1(n11009), .ip2(n9850), .ip3(n11308), .ip4(n11295), .op(
        n9112) );
  inv_1 U11009 ( .ip(n12658), .op(n9844) );
  inv_1 U11010 ( .ip(n12659), .op(n9847) );
  nand4_1 U11011 ( .ip1(n9853), .ip2(n9844), .ip3(n9847), .ip4(n11255), .op(
        n9111) );
  nor4_1 U11012 ( .ip1(n9114), .ip2(n9113), .ip3(n9112), .ip4(n9111), .op(
        n9115) );
  nand4_1 U11013 ( .ip1(n9118), .ip2(n9117), .ip3(n9116), .ip4(n9115), .op(
        n9121) );
  nor3_1 U11014 ( .ip1(n9123), .ip2(n11511), .ip3(n9122), .op(n11455) );
  nand2_1 U11015 ( .ip1(n11481), .ip2(\CORTEXM0DS_INST/vis_ipsr [5]), .op(
        n9120) );
  nand2_1 U11016 ( .ip1(n11549), .ip2(n12675), .op(n9119) );
  nand2_1 U11017 ( .ip1(n9120), .ip2(n9119), .op(n11400) );
  not_ab_or_c_or_d U11018 ( .ip1(n11549), .ip2(n9121), .ip3(n11455), .ip4(
        n11400), .op(n9124) );
  nand3_1 U11019 ( .ip1(n9123), .ip2(n11513), .ip3(n9122), .op(n11452) );
  nand3_1 U11020 ( .ip1(n11399), .ip2(n9124), .ip3(n11452), .op(n9125) );
  nor4_1 U11021 ( .ip1(n11384), .ip2(n11336), .ip3(n11251), .ip4(n9125), .op(
        n9126) );
  nand4_1 U11022 ( .ip1(n9129), .ip2(n9128), .ip3(n9127), .ip4(n9126), .op(
        n9204) );
  or2_1 U11023 ( .ip1(n11545), .ip2(n12240), .op(n9131) );
  inv_1 U11024 ( .ip(n11406), .op(n9199) );
  or2_1 U11025 ( .ip1(n9199), .ip2(n12240), .op(n9130) );
  nand2_1 U11026 ( .ip1(n9131), .ip2(n9130), .op(n11408) );
  inv_1 U11027 ( .ip(n12175), .op(n9133) );
  nand2_1 U11028 ( .ip1(n9133), .ip2(n9132), .op(n11330) );
  nand2_1 U11029 ( .ip1(n9135), .ip2(n9134), .op(n11309) );
  inv_1 U11030 ( .ip(n9136), .op(n11510) );
  or2_1 U11031 ( .ip1(n12114), .ip2(n11510), .op(n11518) );
  inv_1 U11032 ( .ip(n9804), .op(n9138) );
  nand2_1 U11033 ( .ip1(n9138), .ip2(n9137), .op(n11289) );
  nand4_1 U11034 ( .ip1(n11330), .ip2(n11309), .ip3(n11518), .ip4(n11289), 
        .op(n9152) );
  nand2_1 U11035 ( .ip1(n12222), .ip2(n9139), .op(n11382) );
  inv_1 U11036 ( .ip(n9140), .op(n11317) );
  or2_1 U11037 ( .ip1(n11319), .ip2(n11317), .op(n11323) );
  inv_1 U11038 ( .ip(n9141), .op(n11340) );
  or2_1 U11039 ( .ip1(n11342), .ip2(n11340), .op(n11346) );
  inv_1 U11040 ( .ip(n10964), .op(n11539) );
  nand2_1 U11041 ( .ip1(n11539), .ip2(n11540), .op(n11536) );
  nand4_1 U11042 ( .ip1(n11382), .ip2(n11323), .ip3(n11346), .ip4(n11536), 
        .op(n9151) );
  inv_1 U11043 ( .ip(n9142), .op(n11363) );
  nor2_1 U11044 ( .ip1(n11366), .ip2(n11363), .op(n11370) );
  inv_1 U11045 ( .ip(n9143), .op(n11270) );
  nor2_1 U11046 ( .ip1(n12141), .ip2(n11270), .op(n11277) );
  nor4_1 U11047 ( .ip1(n11435), .ip2(n11457), .ip3(n11370), .ip4(n11277), .op(
        n9149) );
  nand2_1 U11048 ( .ip1(n12201), .ip2(n9144), .op(n11357) );
  inv_1 U11049 ( .ip(n12134), .op(n9146) );
  nand2_1 U11050 ( .ip1(n9146), .ip2(n9145), .op(n11264) );
  nand2_1 U11051 ( .ip1(n9148), .ip2(n9147), .op(n11299) );
  nand4_1 U11052 ( .ip1(n9149), .ip2(n11357), .ip3(n11264), .ip4(n11299), .op(
        n9150) );
  or4_1 U11053 ( .ip1(n11408), .ip2(n9152), .ip3(n9151), .ip4(n9150), .op(
        n9168) );
  nor2_1 U11054 ( .ip1(n11530), .ip2(n10856), .op(n9158) );
  nand3_1 U11055 ( .ip1(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip3(
        \CORTEXM0DS_INST/cm0_control[1] ), .op(n9153) );
  or2_1 U11056 ( .ip1(n9153), .ip2(n11478), .op(n9156) );
  nand3_1 U11057 ( .ip1(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip2(
        \CORTEXM0DS_INST/vis_ipsr [1]), .ip3(n12065), .op(n9154) );
  or2_1 U11058 ( .ip1(n9154), .ip2(n11478), .op(n9155) );
  nand2_1 U11059 ( .ip1(n9156), .ip2(n9155), .op(n9157) );
  or2_1 U11060 ( .ip1(n9158), .ip2(n9157), .op(n11486) );
  nand2_1 U11061 ( .ip1(\CORTEXM0DS_INST/vis_apsr [0]), .ip2(n11450), .op(
        n9167) );
  nor2_1 U11062 ( .ip1(n9163), .ip2(n11511), .op(n9162) );
  nand2_1 U11063 ( .ip1(n9159), .ip2(n11434), .op(n9161) );
  mux2_1 U11064 ( .ip1(n9162), .ip2(n9161), .s(n9160), .op(n9165) );
  nand2_1 U11065 ( .ip1(n11545), .ip2(n9163), .op(n9164) );
  nand2_1 U11066 ( .ip1(n9165), .ip2(n9164), .op(n9166) );
  nand3_1 U11067 ( .ip1(n9167), .ip2(n9166), .ip3(n11451), .op(n11463) );
  not_ab_or_c_or_d U11068 ( .ip1(n11537), .ip2(n9168), .ip3(n11486), .ip4(
        n11463), .op(n9202) );
  nand2_1 U11069 ( .ip1(n11538), .ip2(n9169), .op(n9173) );
  nor2_1 U11070 ( .ip1(n11513), .ip2(n9169), .op(n9172) );
  nand2_1 U11071 ( .ip1(n11434), .ip2(n9169), .op(n9170) );
  nor2_1 U11072 ( .ip1(n9170), .ip2(n9174), .op(n9171) );
  not_ab_or_c_or_d U11073 ( .ip1(n9174), .ip2(n9173), .ip3(n9172), .ip4(n9171), 
        .op(n11396) );
  nand2_1 U11074 ( .ip1(n11538), .ip2(n9175), .op(n9179) );
  nor2_1 U11075 ( .ip1(n11513), .ip2(n9175), .op(n9178) );
  nand2_1 U11076 ( .ip1(n11434), .ip2(n9175), .op(n9176) );
  nor2_1 U11077 ( .ip1(n9176), .ip2(n9180), .op(n9177) );
  not_ab_or_c_or_d U11078 ( .ip1(n9180), .ip2(n9179), .ip3(n9178), .ip4(n9177), 
        .op(n11252) );
  inv_1 U11079 ( .ip(n9181), .op(n9182) );
  mux2_1 U11080 ( .ip1(n11537), .ip2(n11513), .s(n9182), .op(n9185) );
  nor2_1 U11081 ( .ip1(n9182), .ip2(n11511), .op(n9184) );
  mux2_1 U11082 ( .ip1(n9185), .ip2(n9184), .s(n9183), .op(n11475) );
  nand2_1 U11083 ( .ip1(n9186), .ip2(n11545), .op(n9190) );
  or2_1 U11084 ( .ip1(n9186), .ip2(n11537), .op(n9188) );
  nor2_1 U11085 ( .ip1(n9186), .ip2(n11511), .op(n9187) );
  mux2_1 U11086 ( .ip1(n9188), .ip2(n9187), .s(n9825), .op(n9189) );
  nand2_1 U11087 ( .ip1(n9190), .ip2(n9189), .op(n9192) );
  nand2_1 U11088 ( .ip1(\CORTEXM0DS_INST/vis_apsr [1]), .ip2(n11450), .op(
        n9191) );
  nand2_1 U11089 ( .ip1(n9192), .ip2(n9191), .op(n11446) );
  nor4_1 U11090 ( .ip1(n11396), .ip2(n11252), .ip3(n11475), .ip4(n11446), .op(
        n9201) );
  nor2_1 U11091 ( .ip1(n9196), .ip2(n11511), .op(n9195) );
  nand2_1 U11092 ( .ip1(n9193), .ip2(n11434), .op(n9194) );
  mux2_1 U11093 ( .ip1(n9195), .ip2(n9194), .s(n12274), .op(n9198) );
  nand2_1 U11094 ( .ip1(n11545), .ip2(n9196), .op(n9197) );
  nand2_1 U11095 ( .ip1(n9198), .ip2(n9197), .op(n11443) );
  nand2_1 U11096 ( .ip1(n9199), .ip2(n11408), .op(n9200) );
  nand4_1 U11097 ( .ip1(n9202), .ip2(n9201), .ip3(n11443), .ip4(n9200), .op(
        n9203) );
  nor4_1 U11098 ( .ip1(n11155), .ip2(n11471), .ip3(n9204), .ip4(n9203), .op(
        n9239) );
  xor2_1 U11099 ( .ip1(n9206), .ip2(n9205), .op(n12103) );
  xor2_1 U11100 ( .ip1(n9208), .ip2(n9207), .op(n12162) );
  xor2_1 U11101 ( .ip1(n9210), .ip2(n9209), .op(n12182) );
  xor2_1 U11102 ( .ip1(n9212), .ip2(n9211), .op(n11302) );
  xor2_1 U11103 ( .ip1(n9214), .ip2(n9213), .op(n12243) );
  xor2_1 U11104 ( .ip1(n9216), .ip2(n9215), .op(n12230) );
  or4_1 U11105 ( .ip1(n12243), .ip2(n12230), .ip3(n11476), .ip4(n11390), .op(
        n9224) );
  xor2_1 U11106 ( .ip1(n9218), .ip2(n9217), .op(n12137) );
  xor2_1 U11107 ( .ip1(n9220), .ip2(n9219), .op(n12117) );
  xor2_1 U11108 ( .ip1(n9222), .ip2(n9221), .op(n12147) );
  or3_1 U11109 ( .ip1(n12137), .ip2(n12117), .ip3(n12147), .op(n9223) );
  nor4_1 U11110 ( .ip1(n11302), .ip2(n11397), .ip3(n9224), .ip4(n9223), .op(
        n9230) );
  xor2_1 U11111 ( .ip1(n9226), .ip2(n9225), .op(n12168) );
  xor2_1 U11112 ( .ip1(n9228), .ip2(n9227), .op(n9943) );
  nand4_1 U11113 ( .ip1(n9230), .ip2(n12168), .ip3(n9943), .ip4(n9229), .op(
        n9231) );
  nor3_1 U11114 ( .ip1(n12162), .ip2(n12182), .ip3(n9231), .op(n9234) );
  xor2_1 U11115 ( .ip1(n9233), .ip2(n9232), .op(n12209) );
  nand3_1 U11116 ( .ip1(n12103), .ip2(n9234), .ip3(n12209), .op(n9235) );
  nand2_1 U11117 ( .ip1(n9235), .ip2(n11534), .op(n9238) );
  xor2_1 U11118 ( .ip1(n9237), .ip2(n9236), .op(n10063) );
  nand2_1 U11119 ( .ip1(n10063), .ip2(n11534), .op(n11448) );
  nand4_1 U11120 ( .ip1(n11259), .ip2(n9239), .ip3(n9238), .ip4(n11448), .op(
        n9254) );
  xnor2_1 U11121 ( .ip1(n9241), .ip2(n9240), .op(n12310) );
  nor2_1 U11122 ( .ip1(n11530), .ip2(n12310), .op(n11416) );
  xnor2_1 U11123 ( .ip1(n9243), .ip2(n9242), .op(n12219) );
  nor2_1 U11124 ( .ip1(n11530), .ip2(n12219), .op(n11381) );
  xnor2_1 U11125 ( .ip1(n9245), .ip2(n9244), .op(n12198) );
  nor2_1 U11126 ( .ip1(n11530), .ip2(n12198), .op(n11355) );
  xor2_1 U11127 ( .ip1(n9247), .ip2(n9246), .op(n12189) );
  nor2_1 U11128 ( .ip1(n11530), .ip2(n12189), .op(n11350) );
  nor4_1 U11129 ( .ip1(n11416), .ip2(n11381), .ip3(n11355), .ip4(n11350), .op(
        n9252) );
  xor2_1 U11130 ( .ip1(n9249), .ip2(n9248), .op(n10571) );
  nand2_1 U11131 ( .ip1(n10571), .ip2(n11534), .op(n11459) );
  nand2_1 U11132 ( .ip1(n10071), .ip2(n11534), .op(n11466) );
  xor2_1 U11133 ( .ip1(n9251), .ip2(n9250), .op(n12262) );
  nand2_1 U11134 ( .ip1(n12262), .ip2(n11534), .op(n11438) );
  nand4_1 U11135 ( .ip1(n9252), .ip2(n11459), .ip3(n11466), .ip4(n11438), .op(
        n9253) );
  nor4_1 U11136 ( .ip1(n11441), .ip2(n11421), .ip3(n9254), .ip4(n9253), .op(
        n9458) );
  nor2_1 U11137 ( .ip1(n10055), .ip2(n9476), .op(n9255) );
  not_ab_or_c_or_d U11138 ( .ip1(n9476), .ip2(n9256), .ip3(n9361), .ip4(n9255), 
        .op(n9456) );
  nor2_1 U11139 ( .ip1(n9296), .ip2(n9416), .op(n9262) );
  nor2_1 U11140 ( .ip1(n9293), .ip2(n9420), .op(n9261) );
  nor2_1 U11141 ( .ip1(n9257), .ip2(n9418), .op(n9260) );
  nor2_1 U11142 ( .ip1(n9258), .ip2(n9392), .op(n9259) );
  nor4_1 U11143 ( .ip1(n9262), .ip2(n9261), .ip3(n9260), .ip4(n9259), .op(
        n9343) );
  nand2_1 U11144 ( .ip1(n9429), .ip2(n9263), .op(n9268) );
  nand2_1 U11145 ( .ip1(n9431), .ip2(n9264), .op(n9267) );
  nand2_1 U11146 ( .ip1(n9433), .ip2(n9282), .op(n9266) );
  nand2_1 U11147 ( .ip1(n9435), .ip2(n9281), .op(n9265) );
  nand4_1 U11148 ( .ip1(n9268), .ip2(n9267), .ip3(n9266), .ip4(n9265), .op(
        n9301) );
  nor2_1 U11149 ( .ip1(n9443), .ip2(n9301), .op(n9921) );
  nand4_1 U11150 ( .ip1(n9339), .ip2(n9987), .ip3(n9343), .ip4(n9921), .op(
        n9290) );
  nand2_1 U11151 ( .ip1(n9429), .ip2(n9276), .op(n9274) );
  nand2_1 U11152 ( .ip1(n9433), .ip2(n9269), .op(n9273) );
  nand2_1 U11153 ( .ip1(n9431), .ip2(n9275), .op(n9272) );
  nand2_1 U11154 ( .ip1(n9435), .ip2(n9270), .op(n9271) );
  nand4_1 U11155 ( .ip1(n9274), .ip2(n9273), .ip3(n9272), .ip4(n9271), .op(
        n10183) );
  nor2_1 U11156 ( .ip1(n9982), .ip2(n10183), .op(n9427) );
  nand2_1 U11157 ( .ip1(n9429), .ip2(n9284), .op(n9280) );
  nand2_1 U11158 ( .ip1(n9431), .ip2(n9283), .op(n9279) );
  nand2_1 U11159 ( .ip1(n9433), .ip2(n9275), .op(n9278) );
  nand2_1 U11160 ( .ip1(n9435), .ip2(n9276), .op(n9277) );
  nand4_1 U11161 ( .ip1(n9280), .ip2(n9279), .ip3(n9278), .ip4(n9277), .op(
        n9442) );
  nor2_1 U11162 ( .ip1(n9338), .ip2(n9442), .op(n9920) );
  nand3_1 U11163 ( .ip1(n9292), .ip2(n9427), .ip3(n9920), .op(n9289) );
  nand2_1 U11164 ( .ip1(n9429), .ip2(n9281), .op(n9288) );
  nand2_1 U11165 ( .ip1(n9431), .ip2(n9282), .op(n9287) );
  nand2_1 U11166 ( .ip1(n9433), .ip2(n9283), .op(n9286) );
  nand2_1 U11167 ( .ip1(n9435), .ip2(n9284), .op(n9285) );
  nand4_1 U11168 ( .ip1(n9288), .ip2(n9287), .ip3(n9286), .ip4(n9285), .op(
        n10185) );
  not_ab_or_c_or_d U11169 ( .ip1(n9290), .ip2(n9289), .ip3(n9994), .ip4(n10185), .op(n9302) );
  mux2_1 U11170 ( .ip1(n9292), .ip2(n9291), .s(n9443), .op(n9467) );
  nor2_1 U11171 ( .ip1(n9293), .ip2(n9418), .op(n9300) );
  nor2_1 U11172 ( .ip1(n9294), .ip2(n9420), .op(n9299) );
  nor2_1 U11173 ( .ip1(n9295), .ip2(n9416), .op(n9298) );
  nor2_1 U11174 ( .ip1(n9296), .ip2(n9392), .op(n9297) );
  or4_1 U11175 ( .ip1(n9300), .ip2(n9299), .ip3(n9298), .ip4(n9297), .op(n9309) );
  mux2_1 U11176 ( .ip1(n9309), .ip2(n9301), .s(n9443), .op(n9475) );
  inv_1 U11177 ( .ip(n9475), .op(n10258) );
  nand3_1 U11178 ( .ip1(n9302), .ip2(n9467), .ip3(n10258), .op(n9455) );
  nand2_1 U11179 ( .ip1(n9431), .ip2(n9303), .op(n9308) );
  nand2_1 U11180 ( .ip1(n9433), .ip2(n9330), .op(n9307) );
  nand2_1 U11181 ( .ip1(n9429), .ip2(n9304), .op(n9306) );
  nand2_1 U11182 ( .ip1(n9435), .ip2(n9329), .op(n9305) );
  nand4_1 U11183 ( .ip1(n9308), .ip2(n9307), .ip3(n9306), .ip4(n9305), .op(
        n9356) );
  mux2_1 U11184 ( .ip1(n9356), .ip2(n9309), .s(n9443), .op(n9310) );
  mux2_1 U11185 ( .ip1(n9362), .ip2(n9310), .s(n9346), .op(n9930) );
  nor2_1 U11186 ( .ip1(n9311), .ip2(n9338), .op(n9313) );
  mux2_1 U11187 ( .ip1(n9357), .ip2(n9312), .s(n9435), .op(n10005) );
  not_ab_or_c_or_d U11188 ( .ip1(n9338), .ip2(n9383), .ip3(n9313), .ip4(n10005), .op(n10006) );
  nor4_1 U11189 ( .ip1(n9315), .ip2(n9930), .ip3(n10006), .ip4(n9314), .op(
        n9316) );
  or2_1 U11190 ( .ip1(n9316), .ip2(n9361), .op(n9360) );
  nor2_1 U11191 ( .ip1(n9317), .ip2(n9418), .op(n9324) );
  nor2_1 U11192 ( .ip1(n9318), .ip2(n9420), .op(n9323) );
  nor2_1 U11193 ( .ip1(n9319), .ip2(n9416), .op(n9322) );
  nor2_1 U11194 ( .ip1(n9320), .ip2(n9392), .op(n9321) );
  nor4_1 U11195 ( .ip1(n9324), .ip2(n9323), .ip3(n9322), .ip4(n9321), .op(
        n10216) );
  inv_1 U11196 ( .ip(n9325), .op(n9328) );
  nor2_1 U11197 ( .ip1(n9338), .ip2(n9345), .op(n9327) );
  nor2_1 U11198 ( .ip1(n9328), .ip2(n9327), .op(n9326) );
  not_ab_or_c_or_d U11199 ( .ip1(n9328), .ip2(n9327), .ip3(n11730), .ip4(n9326), .op(n10108) );
  nand2_1 U11200 ( .ip1(n9429), .ip2(n9329), .op(n9336) );
  nand2_1 U11201 ( .ip1(n9431), .ip2(n9330), .op(n9335) );
  nand2_1 U11202 ( .ip1(n9433), .ip2(n9331), .op(n9334) );
  nand2_1 U11203 ( .ip1(n9435), .ip2(n9332), .op(n9333) );
  nand4_1 U11204 ( .ip1(n9336), .ip2(n9335), .ip3(n9334), .ip4(n9333), .op(
        n9344) );
  nor2_1 U11205 ( .ip1(n9344), .ip2(n9338), .op(n9337) );
  not_ab_or_c_or_d U11206 ( .ip1(n9338), .ip2(n10216), .ip3(n10108), .ip4(
        n9337), .op(n10104) );
  mux2_1 U11207 ( .ip1(n9340), .ip2(n9339), .s(n9443), .op(n9341) );
  inv_1 U11208 ( .ip(n9341), .op(n9473) );
  mux2_1 U11209 ( .ip1(n9346), .ip2(n9347), .s(n9420), .op(n9342) );
  mux2_1 U11210 ( .ip1(n9362), .ip2(n9473), .s(n9342), .op(n11822) );
  inv_1 U11211 ( .ip(n9343), .op(n10094) );
  mux2_1 U11212 ( .ip1(n9344), .ip2(n10094), .s(n9443), .op(n9349) );
  mux2_1 U11213 ( .ip1(n9347), .ip2(n9346), .s(n9345), .op(n9348) );
  mux2_1 U11214 ( .ip1(n9362), .ip2(n9349), .s(n9348), .op(n10182) );
  inv_1 U11215 ( .ip(n9350), .op(n9404) );
  nand2_1 U11216 ( .ip1(n9429), .ip2(n9404), .op(n9355) );
  nand2_1 U11217 ( .ip1(n9433), .ip2(n9377), .op(n9354) );
  nand2_1 U11218 ( .ip1(n9431), .ip2(n9402), .op(n9353) );
  nand2_1 U11219 ( .ip1(n9435), .ip2(n9351), .op(n9352) );
  nand4_1 U11220 ( .ip1(n9355), .ip2(n9354), .ip3(n9353), .ip4(n9352), .op(
        n9382) );
  mux2_1 U11221 ( .ip1(n9382), .ip2(n9356), .s(n9443), .op(n9486) );
  mux2_1 U11222 ( .ip1(n9486), .ip2(n9362), .s(n9357), .op(n10255) );
  nor4_1 U11223 ( .ip1(n10104), .ip2(n11822), .ip3(n10182), .ip4(n10255), .op(
        n9358) );
  or2_1 U11224 ( .ip1(n9358), .ip2(n9361), .op(n9359) );
  nand2_1 U11225 ( .ip1(n9360), .ip2(n9359), .op(n9454) );
  nor2_1 U11226 ( .ip1(n9361), .ip2(n10048), .op(n9495) );
  nor2_1 U11227 ( .ip1(n9361), .ip2(n9874), .op(n9490) );
  nor2_1 U11228 ( .ip1(n9495), .ip2(n9490), .op(n10044) );
  nand2_1 U11229 ( .ip1(n9362), .ip2(n10044), .op(n9489) );
  or2_1 U11230 ( .ip1(n10055), .ip2(n9387), .op(n9413) );
  nand2_1 U11231 ( .ip1(n9429), .ip2(n9370), .op(n9366) );
  nand2_1 U11232 ( .ip1(n9431), .ip2(n9367), .op(n9365) );
  nand2_1 U11233 ( .ip1(n9433), .ip2(n9401), .op(n9364) );
  nand2_1 U11234 ( .ip1(n9435), .ip2(n9403), .op(n9363) );
  nand4_1 U11235 ( .ip1(n9366), .ip2(n9365), .ip3(n9364), .ip4(n9363), .op(
        n11608) );
  nand2_1 U11236 ( .ip1(n9433), .ip2(n9367), .op(n9374) );
  nand2_1 U11237 ( .ip1(n9431), .ip2(n9368), .op(n9373) );
  nand2_1 U11238 ( .ip1(n9429), .ip2(n9369), .op(n9372) );
  nand2_1 U11239 ( .ip1(n9435), .ip2(n9370), .op(n9371) );
  nand4_1 U11240 ( .ip1(n9374), .ip2(n9373), .ip3(n9372), .ip4(n9371), .op(
        n10110) );
  nor2_1 U11241 ( .ip1(n9998), .ip2(n10110), .op(n9415) );
  inv_1 U11242 ( .ip(n9415), .op(n9375) );
  nor3_1 U11243 ( .ip1(n11608), .ip2(n9376), .ip3(n9375), .op(n9385) );
  nand2_1 U11244 ( .ip1(n9433), .ip2(n9404), .op(n9381) );
  nand2_1 U11245 ( .ip1(n9431), .ip2(n9403), .op(n9380) );
  nand2_1 U11246 ( .ip1(n9429), .ip2(n9402), .op(n9379) );
  nand2_1 U11247 ( .ip1(n9435), .ip2(n9377), .op(n9378) );
  nand4_1 U11248 ( .ip1(n9381), .ip2(n9380), .ip3(n9379), .ip4(n9378), .op(
        n9400) );
  inv_1 U11249 ( .ip(n9400), .op(n11599) );
  inv_1 U11250 ( .ip(n9382), .op(n11615) );
  and4_1 U11251 ( .ip1(n11599), .ip2(n11615), .ip3(n9383), .ip4(n10216), .op(
        n9384) );
  mux2_1 U11252 ( .ip1(n9385), .ip2(n9384), .s(n9443), .op(n9388) );
  nor2_1 U11253 ( .ip1(n9387), .ip2(n9386), .op(n9409) );
  or2_1 U11254 ( .ip1(n9388), .ip2(n9409), .op(n9412) );
  nor2_1 U11255 ( .ip1(n9389), .ip2(n9416), .op(n9397) );
  nor2_1 U11256 ( .ip1(n9390), .ip2(n9420), .op(n9396) );
  nor2_1 U11257 ( .ip1(n9391), .ip2(n9418), .op(n9395) );
  nor2_1 U11258 ( .ip1(n9393), .ip2(n9392), .op(n9394) );
  nor4_1 U11259 ( .ip1(n9397), .ip2(n9396), .ip3(n9395), .ip4(n9394), .op(
        n9914) );
  inv_1 U11260 ( .ip(n9914), .op(n9398) );
  mux2_1 U11261 ( .ip1(n9398), .ip2(n11608), .s(n9443), .op(n10271) );
  mux2_1 U11262 ( .ip1(n9400), .ip2(n9399), .s(n9443), .op(n9468) );
  nand2_1 U11263 ( .ip1(n9431), .ip2(n9401), .op(n9408) );
  nand2_1 U11264 ( .ip1(n9433), .ip2(n9402), .op(n9407) );
  nand2_1 U11265 ( .ip1(n9429), .ip2(n9403), .op(n9406) );
  nand2_1 U11266 ( .ip1(n9435), .ip2(n9404), .op(n9405) );
  nand4_1 U11267 ( .ip1(n9408), .ip2(n9407), .ip3(n9406), .ip4(n9405), .op(
        n10219) );
  nor4_1 U11268 ( .ip1(n10271), .ip2(n9468), .ip3(n9999), .ip4(n10219), .op(
        n9410) );
  or2_1 U11269 ( .ip1(n9410), .ip2(n9409), .op(n9411) );
  nand2_1 U11270 ( .ip1(n9412), .ip2(n9411), .op(n9446) );
  or2_1 U11271 ( .ip1(n9413), .ip2(n9446), .op(n9449) );
  nand3_1 U11272 ( .ip1(n9914), .ip2(n9415), .ip3(n9414), .op(n9441) );
  nor2_1 U11273 ( .ip1(n9417), .ip2(n9416), .op(n9425) );
  nor2_1 U11274 ( .ip1(n9419), .ip2(n9418), .op(n9424) );
  nor2_1 U11275 ( .ip1(n9421), .ip2(n9420), .op(n9423) );
  and2_1 U11276 ( .ip1(n9428), .ip2(n9435), .op(n9422) );
  nor4_1 U11277 ( .ip1(n9425), .ip2(n9424), .ip3(n9423), .ip4(n9422), .op(
        n9913) );
  nand3_1 U11278 ( .ip1(n9427), .ip2(n9913), .ip3(n9426), .op(n9440) );
  nand2_1 U11279 ( .ip1(n9429), .ip2(n9428), .op(n9439) );
  nand2_1 U11280 ( .ip1(n9431), .ip2(n9430), .op(n9438) );
  nand2_1 U11281 ( .ip1(n9433), .ip2(n9432), .op(n9437) );
  nand2_1 U11282 ( .ip1(n9435), .ip2(n9434), .op(n9436) );
  nand4_1 U11283 ( .ip1(n9439), .ip2(n9438), .ip3(n9437), .ip4(n9436), .op(
        n10095) );
  not_ab_or_c_or_d U11284 ( .ip1(n9441), .ip2(n9440), .ip3(n9978), .ip4(n10095), .op(n9445) );
  inv_1 U11285 ( .ip(n9442), .op(n9444) );
  mux2_1 U11286 ( .ip1(n9444), .ip2(n9913), .s(n9443), .op(n11623) );
  nand3_1 U11287 ( .ip1(n9445), .ip2(n11623), .ip3(n9470), .op(n9447) );
  or2_1 U11288 ( .ip1(n9447), .ip2(n9446), .op(n9448) );
  nand2_1 U11289 ( .ip1(n9449), .ip2(n9448), .op(n9450) );
  or2_1 U11290 ( .ip1(n9451), .ip2(n9450), .op(n9452) );
  nand3_1 U11291 ( .ip1(n9489), .ip2(\CORTEXM0DS_INST/u_logic/Dw8vx4 ), .ip3(
        n9452), .op(n9453) );
  not_ab_or_c_or_d U11292 ( .ip1(n9456), .ip2(n9455), .ip3(n9454), .ip4(n9453), 
        .op(n9457) );
  not_ab_or_c_or_d U11293 ( .ip1(n9536), .ip2(n9458), .ip3(n11629), .ip4(n9457), .op(n11634) );
  or2_1 U11294 ( .ip1(n11629), .ip2(n11634), .op(n9461) );
  inv_1 U11295 ( .ip(\CORTEXM0DS_INST/vis_apsr [2]), .op(n9459) );
  or2_1 U11296 ( .ip1(n9459), .ip2(n11634), .op(n9460) );
  nand2_1 U11297 ( .ip1(n9461), .ip2(n9460), .op(n9462) );
  mux2_1 U11298 ( .ip1(n9463), .ip2(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .s(
        n9462), .op(n9557) );
  and2_1 U11299 ( .ip1(n9505), .ip2(n9464), .op(n9510) );
  nor2_1 U11300 ( .ip1(n9466), .ip2(n9465), .op(n9477) );
  inv_1 U11301 ( .ip(n9467), .op(n11788) );
  inv_1 U11302 ( .ip(n9468), .op(n11812) );
  nor2_1 U11303 ( .ip1(n9469), .ip2(n11812), .op(n9472) );
  nor2_1 U11304 ( .ip1(n9479), .ip2(n9470), .op(n9471) );
  not_ab_or_c_or_d U11305 ( .ip1(n9477), .ip2(n11788), .ip3(n9472), .ip4(n9471), .op(n9492) );
  nand2_1 U11306 ( .ip1(n9476), .ip2(n9473), .op(n9474) );
  nand2_1 U11307 ( .ip1(n9492), .ip2(n9474), .op(n9496) );
  inv_1 U11308 ( .ip(n9496), .op(n9488) );
  nand2_1 U11309 ( .ip1(n9476), .ip2(n9475), .op(n9483) );
  inv_1 U11310 ( .ip(n11623), .op(n9478) );
  nand2_1 U11311 ( .ip1(n9478), .ip2(n9477), .op(n9482) );
  inv_1 U11312 ( .ip(n9479), .op(n9480) );
  nand2_1 U11313 ( .ip1(n9480), .ip2(n10271), .op(n9481) );
  nand3_1 U11314 ( .ip1(n9483), .ip2(n9482), .ip3(n9481), .op(n9484) );
  not_ab_or_c_or_d U11315 ( .ip1(n9486), .ip2(n9485), .ip3(n11754), .ip4(n9484), .op(n9487) );
  not_ab_or_c_or_d U11316 ( .ip1(n9488), .ip2(n11754), .ip3(n9487), .ip4(n9510), .op(n9508) );
  inv_1 U11317 ( .ip(n9489), .op(n9494) );
  inv_1 U11318 ( .ip(n9490), .op(n9491) );
  nor2_1 U11319 ( .ip1(n9492), .ip2(n9491), .op(n9493) );
  not_ab_or_c_or_d U11320 ( .ip1(n11822), .ip2(n9495), .ip3(n9494), .ip4(n9493), .op(n9537) );
  nand2_1 U11321 ( .ip1(n11730), .ip2(n9496), .op(n9497) );
  nand2_1 U11322 ( .ip1(n9537), .ip2(n9497), .op(n9507) );
  or2_1 U11323 ( .ip1(n9499), .ip2(n9498), .op(n9501) );
  or2_1 U11324 ( .ip1(n9501), .ip2(n9500), .op(n9502) );
  nand2_1 U11325 ( .ip1(n9503), .ip2(n9502), .op(n9504) );
  nor2_1 U11326 ( .ip1(n9505), .ip2(n9504), .op(n9506) );
  mux2_1 U11327 ( .ip1(n9508), .ip2(n9507), .s(n9506), .op(n9509) );
  not_ab_or_c_or_d U11328 ( .ip1(n9510), .ip2(\CORTEXM0DS_INST/vis_apsr [1]), 
        .ip3(n9514), .ip4(n9509), .op(n9518) );
  or2_1 U11329 ( .ip1(n9512), .ip2(n9511), .op(n9516) );
  fulladder U11330 ( .a(n9545), .b(n9544), .ci(n9513), .co(n9515), .s(n9512)
         );
  and3_1 U11331 ( .ip1(n9516), .ip2(n9515), .ip3(n9514), .op(n9517) );
  nor2_1 U11332 ( .ip1(n9518), .ip2(n9517), .op(n11782) );
  inv_1 U11333 ( .ip(n9519), .op(n10657) );
  or4_1 U11334 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n9520), .ip3(
        n10899), .ip4(n10657), .op(n9533) );
  or2_1 U11335 ( .ip1(n9521), .ip2(n11038), .op(n9523) );
  inv_1 U11336 ( .ip(n12334), .op(n12652) );
  or2_1 U11337 ( .ip1(n12652), .ip2(n11038), .op(n9522) );
  nand2_1 U11338 ( .ip1(n9523), .ip2(n9522), .op(n9532) );
  inv_1 U11339 ( .ip(n9524), .op(n9525) );
  or2_1 U11340 ( .ip1(n11651), .ip2(n9525), .op(n9527) );
  or2_1 U11341 ( .ip1(n10915), .ip2(n9525), .op(n9526) );
  nand2_1 U11342 ( .ip1(n9527), .ip2(n9526), .op(n9528) );
  or2_1 U11343 ( .ip1(n11038), .ip2(n9528), .op(n9529) );
  nand3_1 U11344 ( .ip1(n9531), .ip2(n9530), .ip3(n9529), .op(n9548) );
  not_ab_or_c_or_d U11345 ( .ip1(n10705), .ip2(n9533), .ip3(n9532), .ip4(n9548), .op(n11784) );
  mux2_1 U11346 ( .ip1(n11782), .ip2(\CORTEXM0DS_INST/vis_apsr [1]), .s(n11784), .op(n9534) );
  not_ab_or_c_or_d U11347 ( .ip1(n10742), .ip2(n10758), .ip3(n9535), .ip4(
        n9534), .op(n9556) );
  or2_1 U11348 ( .ip1(\CORTEXM0DS_INST/u_logic/Dw8vx4 ), .ip2(n9536), .op(
        n9539) );
  or2_1 U11349 ( .ip1(n9537), .ip2(n9536), .op(n9538) );
  nand2_1 U11350 ( .ip1(n9539), .ip2(n9538), .op(n11628) );
  mux2_1 U11351 ( .ip1(n11628), .ip2(\CORTEXM0DS_INST/vis_apsr [3]), .s(n11629), .op(n9541) );
  or2_1 U11352 ( .ip1(n9540), .ip2(n9541), .op(n9543) );
  or2_1 U11353 ( .ip1(n10751), .ip2(n9541), .op(n9542) );
  nand2_1 U11354 ( .ip1(n9543), .ip2(n9542), .op(n9554) );
  nand3_1 U11355 ( .ip1(n10421), .ip2(n9545), .ip3(n9544), .op(n9547) );
  or3_1 U11356 ( .ip1(n10421), .ip2(n9545), .ip3(n9544), .op(n9546) );
  nand2_1 U11357 ( .ip1(n9547), .ip2(n9546), .op(n11012) );
  inv_1 U11358 ( .ip(n11715), .op(n10439) );
  nand2_1 U11359 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Vdgvx4 ), .op(n12653) );
  nor3_1 U11360 ( .ip1(n10892), .ip2(n10439), .ip3(n12653), .op(n9549) );
  not_ab_or_c_or_d U11361 ( .ip1(n12607), .ip2(n9550), .ip3(n9549), .ip4(n9548), .op(n11013) );
  mux2_1 U11362 ( .ip1(n11012), .ip2(\CORTEXM0DS_INST/vis_apsr [0]), .s(n11013), .op(n9551) );
  nor3_1 U11363 ( .ip1(n9692), .ip2(n9552), .ip3(n9551), .op(n9553) );
  xor2_1 U11364 ( .ip1(n9554), .ip2(n9553), .op(n9555) );
  not_ab_or_c_or_d U11365 ( .ip1(n9557), .ip2(n12580), .ip3(n9556), .ip4(n9555), .op(n9558) );
  mux2_1 U11366 ( .ip1(n9754), .ip2(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .s(
        n9558), .op(n10916) );
  nor3_1 U11367 ( .ip1(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip2(n9559), .ip3(
        n10916), .op(n9564) );
  nand2_1 U11368 ( .ip1(n12584), .ip2(n10869), .op(n9561) );
  inv_1 U11369 ( .ip(\CORTEXM0DS_INST/u_logic/W49vx4 ), .op(n12554) );
  nand4_1 U11370 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n12570), .ip3(
        n12554), .ip4(n12564), .op(n10759) );
  nor4_1 U11371 ( .ip1(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/P39vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/I29vx4 ), .ip4(n11046), .op(n9678) );
  nand4_1 U11372 ( .ip1(n9678), .ip2(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip3(
        n12564), .ip4(n12558), .op(n10459) );
  nor3_1 U11373 ( .ip1(n12584), .ip2(n10759), .ip3(n10459), .op(n9560) );
  not_ab_or_c_or_d U11374 ( .ip1(n12580), .ip2(n9561), .ip3(n9560), .ip4(
        n12530), .op(n9562) );
  nor2_1 U11375 ( .ip1(n9562), .ip2(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .op(
        n9563) );
  nor2_1 U11376 ( .ip1(n9564), .ip2(n9563), .op(n9565) );
  nor2_1 U11377 ( .ip1(n9565), .ip2(n12329), .op(n9568) );
  nor2_1 U11378 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n10612), .op(
        n10615) );
  nor3_1 U11379 ( .ip1(n9566), .ip2(n10615), .ip3(n10782), .op(n9567) );
  not_ab_or_c_or_d U11380 ( .ip1(n10462), .ip2(n10951), .ip3(n9568), .ip4(
        n9567), .op(n9569) );
  nor2_1 U11381 ( .ip1(n9569), .ip2(n12615), .op(n9576) );
  nor2_1 U11382 ( .ip1(n12075), .ip2(n12588), .op(n12074) );
  nor3_1 U11383 ( .ip1(n12074), .ip2(n10506), .ip3(n10927), .op(n10473) );
  nor3_1 U11384 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n12616), .ip3(
        n11212), .op(n11710) );
  not_ab_or_c_or_d U11385 ( .ip1(n9570), .ip2(n12079), .ip3(n10473), .ip4(
        n11710), .op(n9574) );
  nand2_1 U11386 ( .ip1(n11033), .ip2(n9571), .op(n10649) );
  nor4_1 U11387 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(n10665), .ip3(
        n12651), .ip4(n10649), .op(n9662) );
  nand2_1 U11388 ( .ip1(n9662), .ip2(n12075), .op(n9573) );
  nand4_1 U11389 ( .ip1(n9574), .ip2(n11758), .ip3(n9573), .ip4(n9572), .op(
        n9575) );
  not_ab_or_c_or_d U11390 ( .ip1(n12686), .ip2(n9577), .ip3(n9576), .ip4(n9575), .op(n9578) );
  and4_1 U11391 ( .ip1(n9841), .ip2(n9580), .ip3(n9579), .ip4(n9578), .op(
        n9581) );
  not_ab_or_c_or_d U11392 ( .ip1(n5938), .ip2(n9582), .ip3(1'b0), .ip4(n9581), 
        .op(\CORTEXM0DS_INST/u_logic/Eyhvx4 ) );
  nor4_1 U11393 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip3(n12625), .ip4(n10588), .op(
        n9583) );
  or2_1 U11394 ( .ip1(n11697), .ip2(n9583), .op(n9586) );
  or2_1 U11395 ( .ip1(n9584), .ip2(n9583), .op(n9585) );
  nand2_1 U11396 ( .ip1(n9586), .ip2(n9585), .op(n9587) );
  nor2_1 U11397 ( .ip1(n9587), .ip2(n10908), .op(n9648) );
  nor2_1 U11398 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(n11726), .op(
        n10595) );
  inv_1 U11399 ( .ip(n10595), .op(n9590) );
  nand2_1 U11400 ( .ip1(n6210), .ip2(n12618), .op(n9588) );
  nand4_1 U11401 ( .ip1(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip3(n10908), .ip4(n9588), .op(
        n9589) );
  not_ab_or_c_or_d U11402 ( .ip1(n9590), .ip2(n9589), .ip3(
        \CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip4(n10770), .op(n9647) );
  or2_1 U11403 ( .ip1(n10685), .ip2(n12329), .op(n9593) );
  nand2_1 U11404 ( .ip1(n10455), .ip2(n12279), .op(n9591) );
  or2_1 U11405 ( .ip1(n9591), .ip2(n12329), .op(n9592) );
  nand2_1 U11406 ( .ip1(n9593), .ip2(n9592), .op(n9596) );
  nor2_1 U11407 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n9594), .op(
        n9595) );
  not_ab_or_c_or_d U11408 ( .ip1(n9639), .ip2(n11186), .ip3(n9596), .ip4(n9595), .op(n9619) );
  not_ab_or_c_or_d U11409 ( .ip1(n9598), .ip2(n11726), .ip3(n9597), .ip4(
        n11231), .op(n9611) );
  nor2_1 U11410 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n12592), .op(
        n10806) );
  nand2_1 U11411 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n12564), .op(
        n9599) );
  nand3_1 U11412 ( .ip1(n9599), .ip2(n10882), .ip3(n9754), .op(n9600) );
  nand2_1 U11413 ( .ip1(n10806), .ip2(n9600), .op(n9601) );
  or2_1 U11414 ( .ip1(n9601), .ip2(n10605), .op(n9604) );
  nand2_1 U11415 ( .ip1(n10457), .ip2(n10742), .op(n9602) );
  or2_1 U11416 ( .ip1(n9602), .ip2(n10605), .op(n9603) );
  nand2_1 U11417 ( .ip1(n9604), .ip2(n9603), .op(n9610) );
  or2_1 U11418 ( .ip1(n10512), .ip2(n10827), .op(n9607) );
  nand2_1 U11419 ( .ip1(n12554), .ip2(n12564), .op(n9728) );
  nand4_1 U11420 ( .ip1(\CORTEXM0DS_INST/u_logic/R89vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/D69vx4 ), .ip3(n12584), .ip4(n9728), .op(
        n9605) );
  or2_1 U11421 ( .ip1(n9605), .ip2(n10827), .op(n9606) );
  nand2_1 U11422 ( .ip1(n9607), .ip2(n9606), .op(n9608) );
  inv_1 U11423 ( .ip(n10617), .op(n10510) );
  nor2_1 U11424 ( .ip1(n9608), .ip2(n10510), .op(n9609) );
  not_ab_or_c_or_d U11425 ( .ip1(n9611), .ip2(n10587), .ip3(n9610), .ip4(n9609), .op(n9618) );
  nand2_1 U11426 ( .ip1(n11660), .ip2(n10586), .op(n9617) );
  or2_1 U11427 ( .ip1(n10734), .ip2(n10657), .op(n9614) );
  or2_1 U11428 ( .ip1(n9612), .ip2(n10657), .op(n9613) );
  nand2_1 U11429 ( .ip1(n9614), .ip2(n9613), .op(n9615) );
  or2_1 U11430 ( .ip1(n9615), .ip2(n12649), .op(n9616) );
  nand4_1 U11431 ( .ip1(n9619), .ip2(n9618), .ip3(n9617), .ip4(n9616), .op(
        n9646) );
  nand2_1 U11432 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Cf9vx4 ), .op(n10441) );
  nor3_1 U11433 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n12073), .ip3(
        n10441), .op(n9622) );
  nor4_1 U11434 ( .ip1(n9727), .ip2(n9620), .ip3(n12095), .ip4(n10665), .op(
        n9621) );
  not_ab_or_c_or_d U11435 ( .ip1(n9623), .ip2(n12074), .ip3(n9622), .ip4(n9621), .op(n9644) );
  inv_1 U11436 ( .ip(n9653), .op(n9640) );
  inv_1 U11437 ( .ip(n10827), .op(n9628) );
  nor2_1 U11438 ( .ip1(n9754), .ip2(n12570), .op(n10613) );
  nor3_1 U11439 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/K79vx4 ), .ip3(n9754), .op(n10501) );
  or2_1 U11440 ( .ip1(\CORTEXM0DS_INST/u_logic/K79vx4 ), .ip2(n10501), .op(
        n9625) );
  nand2_1 U11441 ( .ip1(n12580), .ip2(n12570), .op(n10783) );
  or2_1 U11442 ( .ip1(n10783), .ip2(n10501), .op(n9624) );
  nand2_1 U11443 ( .ip1(n9625), .ip2(n9624), .op(n9626) );
  nor2_1 U11444 ( .ip1(n10613), .ip2(n9626), .op(n9627) );
  nor2_1 U11445 ( .ip1(n9628), .ip2(n9627), .op(n9632) );
  nor3_1 U11446 ( .ip1(n9629), .ip2(n12588), .ip3(
        \CORTEXM0DS_INST/u_logic/Kg9vx4 ), .op(n9630) );
  nor2_1 U11447 ( .ip1(n9630), .ip2(n10701), .op(n9631) );
  not_ab_or_c_or_d U11448 ( .ip1(n12280), .ip2(
        \CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip3(n9632), .ip4(n9631), .op(n9633) );
  nor2_1 U11449 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(n9633), .op(
        n9638) );
  nor2_1 U11450 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n12631), .op(
        n9636) );
  nor3_1 U11451 ( .ip1(n10751), .ip2(n10749), .ip3(n10441), .op(n9635) );
  inv_1 U11452 ( .ip(n9634), .op(n10597) );
  nor2_1 U11453 ( .ip1(n12388), .ip2(n10597), .op(n11762) );
  or4_1 U11454 ( .ip1(n9636), .ip2(n9635), .ip3(n11762), .ip4(n5428), .op(
        n9637) );
  not_ab_or_c_or_d U11455 ( .ip1(n9640), .ip2(n9639), .ip3(n9638), .ip4(n9637), 
        .op(n9643) );
  inv_1 U11456 ( .ip(n10898), .op(n10592) );
  nand3_1 U11457 ( .ip1(n11744), .ip2(n12606), .ip3(n10592), .op(n9642) );
  nand3_1 U11458 ( .ip1(n9869), .ip2(n11038), .ip3(n10949), .op(n9641) );
  nand4_1 U11459 ( .ip1(n9644), .ip2(n9643), .ip3(n9642), .ip4(n9641), .op(
        n9645) );
  nor4_1 U11460 ( .ip1(n9648), .ip2(n9647), .ip3(n9646), .ip4(n9645), .op(
        n9649) );
  not_ab_or_c_or_d U11461 ( .ip1(n5938), .ip2(n12625), .ip3(1'b0), .ip4(n9649), 
        .op(\CORTEXM0DS_INST/u_logic/Fvhvx4 ) );
  or2_1 U11462 ( .ip1(n11130), .ip2(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .op(
        n12326) );
  nor3_1 U11463 ( .ip1(n10903), .ip2(n10592), .ip3(n12326), .op(n9651) );
  nand2_1 U11464 ( .ip1(n10975), .ip2(n10959), .op(n10909) );
  nor2_1 U11465 ( .ip1(n12095), .ip2(n10909), .op(n9650) );
  not_ab_or_c_or_d U11466 ( .ip1(n9652), .ip2(n10547), .ip3(n9651), .ip4(n9650), .op(n9654) );
  nor2_1 U11467 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n9653), .op(
        n11197) );
  nand2_1 U11468 ( .ip1(n11197), .ip2(n11038), .op(n12341) );
  nand2_1 U11469 ( .ip1(n9654), .ip2(n12341), .op(n9708) );
  nor2_1 U11470 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n12570), .op(
        n9656) );
  nand2_1 U11471 ( .ip1(n9754), .ip2(n12564), .op(n9730) );
  nand4_1 U11472 ( .ip1(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/I29vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/R89vx4 ), .ip4(
        \CORTEXM0DS_INST/u_logic/B19vx4 ), .op(n10745) );
  nor2_1 U11473 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n10745), .op(
        n10879) );
  nor3_1 U11474 ( .ip1(\CORTEXM0DS_INST/u_logic/R89vx4 ), .ip2(n9754), .ip3(
        n12327), .op(n10456) );
  nor2_1 U11475 ( .ip1(n10879), .ip2(n10456), .op(n9655) );
  nor2_1 U11476 ( .ip1(n10756), .ip2(n9655), .op(n10670) );
  not_ab_or_c_or_d U11477 ( .ip1(n9656), .ip2(n9730), .ip3(n9692), .ip4(n10670), .op(n9658) );
  nand2_1 U11478 ( .ip1(n9657), .ip2(n10728), .op(n10706) );
  nor3_1 U11479 ( .ip1(n10612), .ip2(n10506), .ip3(n10706), .op(n10883) );
  inv_1 U11480 ( .ip(n10883), .op(n10950) );
  nor3_1 U11481 ( .ip1(n9658), .ip2(n10950), .ip3(n12075), .op(n9661) );
  nand2_1 U11482 ( .ip1(n9659), .ip2(n10807), .op(n10666) );
  nor3_1 U11483 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n11213), .ip3(
        n10666), .op(n9660) );
  not_ab_or_c_or_d U11484 ( .ip1(n11032), .ip2(n9662), .ip3(n9661), .ip4(n9660), .op(n9677) );
  nor4_1 U11485 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip3(n10865), .ip4(n11729), .op(
        n9830) );
  nor2_1 U11486 ( .ip1(n10676), .ip2(n11130), .op(n9667) );
  nand2_1 U11487 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n10776), .op(
        n9663) );
  not_ab_or_c_or_d U11488 ( .ip1(n9664), .ip2(n9663), .ip3(n11730), .ip4(
        n10900), .op(n9666) );
  nor4_1 U11489 ( .ip1(n9830), .ip2(n9667), .ip3(n9666), .ip4(n9665), .op(
        n9676) );
  nor2_1 U11490 ( .ip1(n9669), .ip2(n9668), .op(n9670) );
  or2_1 U11491 ( .ip1(n11052), .ip2(n9670), .op(n9673) );
  not_ab_or_c_or_d U11492 ( .ip1(n10767), .ip2(n9754), .ip3(n10749), .ip4(
        n12592), .op(n9671) );
  or2_1 U11493 ( .ip1(n9671), .ip2(n9670), .op(n9672) );
  nand2_1 U11494 ( .ip1(n9673), .ip2(n9672), .op(n9674) );
  or2_1 U11495 ( .ip1(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip2(n9674), .op(
        n9675) );
  nand3_1 U11496 ( .ip1(n9677), .ip2(n9676), .ip3(n9675), .op(n9707) );
  inv_1 U11497 ( .ip(n9678), .op(n10760) );
  inv_1 U11498 ( .ip(n10927), .op(n10919) );
  nand2_1 U11499 ( .ip1(n10919), .ip2(n9679), .op(n10868) );
  or4_1 U11500 ( .ip1(n9754), .ip2(n10760), .ip3(n10917), .ip4(n10868), .op(
        n10875) );
  not_ab_or_c_or_d U11501 ( .ip1(\CORTEXM0DS_INST/u_logic/W49vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/K79vx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/R89vx4 ), .ip4(n10875), .op(n9690) );
  or2_1 U11502 ( .ip1(n9680), .ip2(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .op(
        n9685) );
  nand2_1 U11503 ( .ip1(n11068), .ip2(n12592), .op(n10831) );
  nand2_1 U11504 ( .ip1(n10831), .ip2(n9681), .op(n9682) );
  nand4_1 U11505 ( .ip1(n10919), .ip2(n12588), .ip3(n11139), .ip4(n9682), .op(
        n9683) );
  or2_1 U11506 ( .ip1(n9683), .ip2(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .op(
        n9684) );
  nand2_1 U11507 ( .ip1(n9685), .ip2(n9684), .op(n9689) );
  nand2_1 U11508 ( .ip1(n9749), .ip2(n10949), .op(n10474) );
  or2_1 U11509 ( .ip1(n10474), .ip2(n12095), .op(n9687) );
  nand2_1 U11510 ( .ip1(n11697), .ip2(n6210), .op(n10821) );
  or2_1 U11511 ( .ip1(n12608), .ip2(n10821), .op(n9833) );
  or2_1 U11512 ( .ip1(n9833), .ip2(n12095), .op(n9686) );
  nand2_1 U11513 ( .ip1(n9687), .ip2(n9686), .op(n9688) );
  not_ab_or_c_or_d U11514 ( .ip1(n9690), .ip2(n12558), .ip3(n9689), .ip4(n9688), .op(n9705) );
  nand3_1 U11515 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n10726), .ip3(
        n12096), .op(n12325) );
  nand2_1 U11516 ( .ip1(n10972), .ip2(n12032), .op(n9691) );
  nand2_1 U11517 ( .ip1(n12325), .ip2(n9691), .op(n9697) );
  inv_1 U11518 ( .ip(n9692), .op(n10606) );
  nor2_1 U11519 ( .ip1(n10606), .ip2(n11028), .op(n9745) );
  inv_1 U11520 ( .ip(n9745), .op(n9694) );
  nor2_1 U11521 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n10706), .op(
        n10933) );
  inv_1 U11522 ( .ip(n10933), .op(n9693) );
  not_ab_or_c_or_d U11523 ( .ip1(n9695), .ip2(n9694), .ip3(n12588), .ip4(n9693), .op(n9696) );
  not_ab_or_c_or_d U11524 ( .ip1(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip2(
        n10693), .ip3(n10927), .ip4(n10033), .op(n10888) );
  not_ab_or_c_or_d U11525 ( .ip1(n6210), .ip2(n9697), .ip3(n9696), .ip4(n10888), .op(n9704) );
  nand2_1 U11526 ( .ip1(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip2(n9698), .op(
        n9699) );
  nand2_1 U11527 ( .ip1(n10728), .ip2(n12588), .op(n10712) );
  not_ab_or_c_or_d U11528 ( .ip1(n10441), .ip2(n9699), .ip3(n12073), .ip4(
        n10712), .op(n9701) );
  nand3_1 U11529 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n11170), .ip3(
        n11730), .op(n11748) );
  inv_1 U11530 ( .ip(n11035), .op(n10537) );
  nand3_1 U11531 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n10537), .ip3(
        n9700), .op(n9829) );
  nand2_1 U11532 ( .ip1(n11748), .ip2(n9829), .op(n10930) );
  not_ab_or_c_or_d U11533 ( .ip1(n9702), .ip2(n11746), .ip3(n9701), .ip4(
        n10930), .op(n9703) );
  nand3_1 U11534 ( .ip1(n9705), .ip2(n9704), .ip3(n9703), .op(n9706) );
  not_ab_or_c_or_d U11535 ( .ip1(n10820), .ip2(n9708), .ip3(n9707), .ip4(n9706), .op(n9709) );
  not_ab_or_c_or_d U11536 ( .ip1(n5938), .ip2(n10865), .ip3(1'b0), .ip4(n9709), 
        .op(\CORTEXM0DS_INST/u_logic/Ruhvx4 ) );
  nor2_1 U11537 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [10]), .ip2(n9716), 
        .op(n9710) );
  or2_1 U11538 ( .ip1(n12742), .ip2(n9710), .op(n2543) );
  nor2_1 U11539 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [15]), .ip2(n9716), 
        .op(n9711) );
  or2_1 U11540 ( .ip1(n12744), .ip2(n9711), .op(n2463) );
  nor2_1 U11541 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [8]), .ip2(n9716), .op(
        n9712) );
  or2_1 U11542 ( .ip1(n12745), .ip2(n9712), .op(n2511) );
  nor2_1 U11543 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [12]), .ip2(n9716), 
        .op(n9713) );
  or2_1 U11544 ( .ip1(n12746), .ip2(n9713), .op(n2647) );
  nor2_1 U11545 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [0]), .ip2(n9716), .op(
        n9714) );
  or2_1 U11546 ( .ip1(n12747), .ip2(n9714), .op(n2790) );
  nor2_1 U11547 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [3]), .ip2(n9716), .op(
        n9715) );
  or2_1 U11548 ( .ip1(n12748), .ip2(n9715), .op(n2626) );
  nor2_1 U11549 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [6]), .ip2(n9716), .op(
        n9717) );
  or2_1 U11550 ( .ip1(n12749), .ip2(n9717), .op(n2713) );
  nor2_1 U11551 ( .ip1(n11825), .ip2(n12635), .op(n3224) );
  nor2_1 U11552 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [1]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [2]), .op(n11890) );
  nor2_1 U11553 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [16]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [17]), .op(n11974) );
  inv_1 U11554 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [4]), .op(n11896) );
  nand4_1 U11555 ( .ip1(n11890), .ip2(n11974), .ip3(n11896), .ip4(n11894), 
        .op(n9721) );
  nor3_1 U11556 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [12]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [13]), .ip3(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [7]), .op(n11949) );
  nor4_1 U11557 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [9]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [10]), .ip3(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [11]), .ip4(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [8]), .op(n11939) );
  nor4_1 U11558 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [23]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [22]), .ip3(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [21]), .ip4(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [20]), .op(n9719) );
  nor4_1 U11559 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [15]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [14]), .ip3(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [18]), .ip4(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [19]), .op(n9718) );
  nand4_1 U11560 ( .ip1(n11949), .ip2(n11939), .ip3(n9719), .ip4(n9718), .op(
        n9720) );
  nor4_1 U11561 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [6]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [5]), .ip3(n9721), .ip4(n9720), .op(
        n11871) );
  and4_1 U11562 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [0]), .ip2(
        \CORTEXM0DS_INST/u_logic/F2hvx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/S0hvx4 ), .ip4(n11871), .op(n2326) );
  inv_1 U11563 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [7]), .op(n3223) );
  nor3_1 U11564 ( .ip1(n9723), .ip2(n9722), .ip3(n12096), .op(n9724) );
  not_ab_or_c_or_d U11565 ( .ip1(n12079), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip3(n9725), .ip4(n9724), .op(n9726) );
  nor2_1 U11566 ( .ip1(n9726), .ip2(n10949), .op(n9774) );
  nor4_1 U11567 ( .ip1(n10820), .ip2(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip3(
        n9727), .ip4(n11729), .op(n9771) );
  nor2_1 U11568 ( .ip1(n10770), .ip2(n10489), .op(n9770) );
  nor2_1 U11569 ( .ip1(n10760), .ip2(n9728), .op(n9729) );
  nor2_1 U11570 ( .ip1(n9729), .ip2(n12588), .op(n9732) );
  nand4_1 U11571 ( .ip1(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/D69vx4 ), .ip3(n12075), .ip4(n9730), .op(
        n9731) );
  nor4_1 U11572 ( .ip1(\CORTEXM0DS_INST/u_logic/R89vx4 ), .ip2(n9732), .ip3(
        n12327), .ip4(n9731), .op(n9733) );
  nor2_1 U11573 ( .ip1(n9733), .ip2(n12073), .op(n9769) );
  nor2_1 U11574 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(n12570), .op(
        n10743) );
  nand3_1 U11575 ( .ip1(n12584), .ip2(n9754), .ip3(n12564), .op(n10451) );
  nor2_1 U11576 ( .ip1(n10783), .ip2(n10451), .op(n9740) );
  or2_1 U11577 ( .ip1(n9754), .ip2(n12584), .op(n9735) );
  or2_1 U11578 ( .ip1(n10745), .ip2(n12584), .op(n9734) );
  nand2_1 U11579 ( .ip1(n9735), .ip2(n9734), .op(n9736) );
  or2_1 U11580 ( .ip1(n10756), .ip2(n9736), .op(n9738) );
  or2_1 U11581 ( .ip1(\CORTEXM0DS_INST/u_logic/R89vx4 ), .ip2(n9736), .op(
        n9737) );
  nand2_1 U11582 ( .ip1(n9738), .ip2(n9737), .op(n10452) );
  nand3_1 U11583 ( .ip1(n10455), .ip2(n10452), .ip3(n10669), .op(n9739) );
  not_ab_or_c_or_d U11584 ( .ip1(n10743), .ip2(n9741), .ip3(n9740), .ip4(n9739), .op(n9742) );
  nor2_1 U11585 ( .ip1(n12075), .ip2(n9742), .op(n9743) );
  nor2_1 U11586 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(n9743), .op(
        n9744) );
  nor2_1 U11587 ( .ip1(n9744), .ip2(n10506), .op(n9767) );
  nor2_1 U11588 ( .ip1(n11038), .ip2(n12588), .op(n11040) );
  nor2_1 U11589 ( .ip1(n12327), .ip2(n10749), .op(n9746) );
  not_ab_or_c_or_d U11590 ( .ip1(n11040), .ip2(n12584), .ip3(n9746), .ip4(
        n9745), .op(n9747) );
  nor2_1 U11591 ( .ip1(n9747), .ip2(n12075), .op(n9766) );
  or2_1 U11592 ( .ip1(n9748), .ip2(n9749), .op(n9751) );
  or2_1 U11593 ( .ip1(n11038), .ip2(n9749), .op(n9750) );
  nand2_1 U11594 ( .ip1(n9751), .ip2(n9750), .op(n9752) );
  nor2_1 U11595 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n9752), .op(
        n9765) );
  not_ab_or_c_or_d U11596 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(
        n11168), .ip3(n9753), .ip4(n10770), .op(n9756) );
  nor2_1 U11597 ( .ip1(n9754), .ip2(n11029), .op(n9755) );
  not_ab_or_c_or_d U11598 ( .ip1(n9757), .ip2(n11184), .ip3(n9756), .ip4(n9755), .op(n9763) );
  nor2_1 U11599 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n10770), .op(
        n9759) );
  nor3_1 U11600 ( .ip1(n12075), .ip2(n12588), .ip3(n10605), .op(n9758) );
  nor4_1 U11601 ( .ip1(n10029), .ip2(n9759), .ip3(n5428), .ip4(n9758), .op(
        n9762) );
  inv_1 U11602 ( .ip(n10677), .op(n10444) );
  nor2_1 U11603 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n11729), .op(
        n9760) );
  not_ab_or_c_or_d U11604 ( .ip1(n10708), .ip2(n9827), .ip3(n10444), .ip4(
        n9760), .op(n9761) );
  nand4_1 U11605 ( .ip1(n9763), .ip2(n9762), .ip3(n9761), .ip4(n10474), .op(
        n9764) );
  or4_1 U11606 ( .ip1(n9767), .ip2(n9766), .ip3(n9765), .ip4(n9764), .op(n9768) );
  nor4_1 U11607 ( .ip1(n9771), .ip2(n9770), .ip3(n9769), .ip4(n9768), .op(
        n9772) );
  not_ab_or_c_or_d U11608 ( .ip1(n5938), .ip2(n10949), .ip3(1'b0), .ip4(n9772), 
        .op(n9773) );
  or2_1 U11609 ( .ip1(n9774), .ip2(n9773), .op(
        \CORTEXM0DS_INST/u_logic/Qxhvx4 ) );
  inv_1 U11610 ( .ip(\CORTEXM0DS_INST/vis_pc [30]), .op(n9775) );
  nor2_1 U11611 ( .ip1(n10417), .ip2(n9821), .op(n9815) );
  mux2_1 U11612 ( .ip1(n9775), .ip2(\CORTEXM0DS_INST/vis_pc [30]), .s(n9815), 
        .op(n5889) );
  nor2_1 U11613 ( .ip1(n12305), .ip2(n5889), .op(n9779) );
  nand2_1 U11614 ( .ip1(n12300), .ip2(n10421), .op(n9778) );
  nand2_1 U11615 ( .ip1(n12314), .ip2(n9776), .op(n9777) );
  nand2_1 U11616 ( .ip1(n9778), .ip2(n9777), .op(n9824) );
  nor2_1 U11617 ( .ip1(n9779), .ip2(n9824), .op(
        \CORTEXM0DS_INST/u_logic/N4518 ) );
  nor2_1 U11618 ( .ip1(n3227), .ip2(n11825), .op(n9780) );
  nor2_1 U11619 ( .ip1(\CORTEXM0DS_INST/u_logic/Eqgvx4 ), .ip2(n9780), .op(
        n9784) );
  nor3_1 U11620 ( .ip1(n11862), .ip2(n9782), .ip3(n9781), .op(n9783) );
  nor2_1 U11621 ( .ip1(n9784), .ip2(n9783), .op(
        \CORTEXM0DS_INST/u_logic/Owgvx4 ) );
  nand2_1 U11622 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(n12675), .op(
        n6181) );
  nor2_1 U11623 ( .ip1(n11666), .ip2(n6181), .op(n9785) );
  or2_1 U11624 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [5]), .ip2(n9785), .op(
        n9786) );
  nand2_1 U11625 ( .ip1(n9786), .ip2(n2683), .op(n9789) );
  nor2_1 U11626 ( .ip1(n11862), .ip2(n9787), .op(n9788) );
  nor2_1 U11627 ( .ip1(n9789), .ip2(n9788), .op(
        \CORTEXM0DS_INST/u_logic/K1ivx4 ) );
  inv_1 U11628 ( .ip(\interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state [2]), 
        .op(n9791) );
  inv_1 U11629 ( .ip(\interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state [0]), 
        .op(n9800) );
  nand2_1 U11630 ( .ip1(n5939), .ip2(n9800), .op(n9790) );
  nand2_1 U11631 ( .ip1(n9791), .ip2(n9790), .op(
        \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_nextstate [2]) );
  or2_1 U11632 ( .ip1(\interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state [2]), 
        .ip2(n5940), .op(n9798) );
  nand3_1 U11633 ( .ip1(n9798), .ip2(
        \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state [0]), .ip3(
        \interconnect_ip_inst/i_apb_hready_resp ), .op(n9793) );
  or2_1 U11634 ( .ip1(\interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_state [0]), 
        .ip2(\interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_nextstate [2]), .op(
        n9792) );
  nand2_1 U11635 ( .ip1(n9793), .ip2(n9792), .op(\interconnect_ip_inst/n4829 )
         );
  and2_1 U11636 ( .ip1(n5938), .ip2(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [2]), .op(n9794) );
  or2_1 U11637 ( .ip1(n5937), .ip2(n9794), .op(\interconnect_ip_inst/n4862 )
         );
  nand2_1 U11638 ( .ip1(n5938), .ip2(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [3]), .op(n9795) );
  nand2_1 U11639 ( .ip1(n5935), .ip2(n9795), .op(\interconnect_ip_inst/n4863 )
         );
  nand2_1 U11640 ( .ip1(n5938), .ip2(
        \interconnect_ip_inst/i_ahb_U_mux_hsel_prev [4]), .op(n9796) );
  nand2_1 U11641 ( .ip1(n5931), .ip2(n9796), .op(\interconnect_ip_inst/n4864 )
         );
  inv_1 U11642 ( .ip(\interconnect_ip_inst/i_ahb_U_dfltslv_current_state ), 
        .op(n9797) );
  nand2_1 U11643 ( .ip1(n5928), .ip2(n9797), .op(
        \interconnect_ip_inst/i_ahb_U_dfltslv_N4 ) );
  or2_1 U11644 ( .ip1(n5924), .ip2(n9798), .op(n9799) );
  nand2_1 U11645 ( .ip1(n9800), .ip2(n9799), .op(
        \interconnect_ip_inst/i_apb_U_DW_apb_ahbsif_nextstate [0]) );
  nor2_1 U11646 ( .ip1(\interconnect_ip_inst/i_ahb_U_dfltslv_current_state ), 
        .ip2(n5928), .op(\interconnect_ip_inst/n10765 ) );
  nand2_1 U11647 ( .ip1(n9801), .ip2(n12286), .op(
        \CORTEXM0DS_INST/u_logic/N4816 ) );
  nor3_1 U11648 ( .ip1(n12292), .ip2(n12133), .ip3(n9802), .op(n12142) );
  nor2_1 U11649 ( .ip1(\CORTEXM0DS_INST/vis_pc [12]), .ip2(n12142), .op(n9803)
         );
  nor3_1 U11650 ( .ip1(n9803), .ip2(n9807), .ip3(n12305), .op(n9806) );
  nor2_1 U11651 ( .ip1(n9804), .ip2(n12295), .op(n9805) );
  not_ab_or_c_or_d U11652 ( .ip1(n12300), .ip2(n11292), .ip3(n9806), .ip4(
        n9805), .op(\CORTEXM0DS_INST/u_logic/N4767 ) );
  inv_1 U11653 ( .ip(n9807), .op(n9809) );
  inv_1 U11654 ( .ip(\CORTEXM0DS_INST/vis_pc [13]), .op(n10288) );
  inv_1 U11655 ( .ip(n10966), .op(n9808) );
  not_ab_or_c_or_d U11656 ( .ip1(n9809), .ip2(n10288), .ip3(n9808), .ip4(
        n12305), .op(n9812) );
  nor2_1 U11657 ( .ip1(n9810), .ip2(n12295), .op(n9811) );
  not_ab_or_c_or_d U11658 ( .ip1(n12300), .ip2(n11302), .ip3(n9812), .ip4(
        n9811), .op(\CORTEXM0DS_INST/u_logic/N4751 ) );
  nand3_1 U11659 ( .ip1(n9813), .ip2(n1521), .ip3(n11153), .op(
        \CORTEXM0DS_INST/u_logic/N4674 ) );
  inv_1 U11660 ( .ip(\CORTEXM0DS_INST/vis_pc [29]), .op(n10568) );
  nand2_1 U11661 ( .ip1(\CORTEXM0DS_INST/vis_pc [28]), .ip2(n9814), .op(n9819)
         );
  not_ab_or_c_or_d U11662 ( .ip1(n10568), .ip2(n9819), .ip3(n9815), .ip4(
        n12305), .op(n9818) );
  nor2_1 U11663 ( .ip1(n9816), .ip2(n12295), .op(n9817) );
  not_ab_or_c_or_d U11664 ( .ip1(n12300), .ip2(n10571), .ip3(n9818), .ip4(
        n9817), .op(\CORTEXM0DS_INST/u_logic/N4439 ) );
  and2_1 U11665 ( .ip1(n10063), .ip2(n12300), .op(n5888) );
  inv_1 U11666 ( .ip(\CORTEXM0DS_INST/vis_pc [28]), .op(n9822) );
  inv_1 U11667 ( .ip(n9819), .op(n9820) );
  not_ab_or_c_or_d U11668 ( .ip1(n9822), .ip2(n9821), .ip3(n9820), .ip4(n12305), .op(n9823) );
  or2_1 U11669 ( .ip1(n5888), .ip2(n9823), .op(
        \CORTEXM0DS_INST/u_logic/E562z4 ) );
  or2_1 U11670 ( .ip1(n5893), .ip2(n9824), .op(n5894) );
  nor2_1 U11671 ( .ip1(n9825), .ip2(n12295), .op(
        \CORTEXM0DS_INST/u_logic/Q462z4 ) );
  nor2_1 U11672 ( .ip1(n12599), .ip2(n9826), .op(
        \CORTEXM0DS_INST/u_logic/A362z4 ) );
  nor2_1 U11673 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Q5gvx4 ), .op(n10575) );
  nand2_1 U11674 ( .ip1(n9827), .ip2(n10575), .op(n9828) );
  nand2_1 U11675 ( .ip1(n9829), .ip2(n9828), .op(n9843) );
  nor2_1 U11676 ( .ip1(n9831), .ip2(n9830), .op(n9840) );
  nand2_1 U11677 ( .ip1(n12338), .ip2(n11089), .op(n10935) );
  inv_1 U11678 ( .ip(n10935), .op(n9838) );
  or2_1 U11679 ( .ip1(n9832), .ip2(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .op(
        n9835) );
  or2_1 U11680 ( .ip1(n9833), .ip2(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .op(
        n9834) );
  nand2_1 U11681 ( .ip1(n9835), .ip2(n9834), .op(n9837) );
  not_ab_or_c_or_d U11682 ( .ip1(n9838), .ip2(n12626), .ip3(n9837), .ip4(n9836), .op(n9839) );
  nand2_1 U11683 ( .ip1(n10880), .ip2(n10726), .op(n10731) );
  not_ab_or_c_or_d U11684 ( .ip1(n10734), .ip2(n10906), .ip3(n9843), .ip4(
        n9842), .op(\CORTEXM0DS_INST/u_logic/N4396 ) );
  nand2_1 U11685 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(n11472), .op(
        \CORTEXM0DS_INST/u_logic/N4359 ) );
  nand2_1 U11686 ( .ip1(n9863), .ip2(n11472), .op(n6004) );
  nor2_1 U11687 ( .ip1(n9844), .ip2(n9862), .op(n9846) );
  inv_1 U11688 ( .ip(n6004), .op(n9845) );
  not_ab_or_c_or_d U11689 ( .ip1(n12679), .ip2(n11413), .ip3(n9846), .ip4(
        n9845), .op(\CORTEXM0DS_INST/u_logic/N4282 ) );
  nand2_1 U11690 ( .ip1(n9863), .ip2(n12669), .op(n6002) );
  nor2_1 U11691 ( .ip1(n9847), .ip2(n9862), .op(n9849) );
  inv_1 U11692 ( .ip(n6002), .op(n9848) );
  not_ab_or_c_or_d U11693 ( .ip1(n12679), .ip2(n11423), .ip3(n9849), .ip4(
        n9848), .op(\CORTEXM0DS_INST/u_logic/N4227 ) );
  nand2_1 U11694 ( .ip1(n9863), .ip2(n12667), .op(n6000) );
  inv_1 U11695 ( .ip(n9850), .op(n11437) );
  nor2_1 U11696 ( .ip1(n11255), .ip2(n9862), .op(n9852) );
  inv_1 U11697 ( .ip(n6000), .op(n9851) );
  not_ab_or_c_or_d U11698 ( .ip1(n12679), .ip2(n11437), .ip3(n9852), .ip4(
        n9851), .op(\CORTEXM0DS_INST/u_logic/N4170 ) );
  nand2_1 U11699 ( .ip1(n9863), .ip2(n12673), .op(n5998) );
  inv_1 U11700 ( .ip(n9853), .op(n11442) );
  nor2_1 U11701 ( .ip1(n11260), .ip2(n9862), .op(n9855) );
  inv_1 U11702 ( .ip(n5998), .op(n9854) );
  not_ab_or_c_or_d U11703 ( .ip1(n12679), .ip2(n11442), .ip3(n9855), .ip4(
        n9854), .op(\CORTEXM0DS_INST/u_logic/N4116 ) );
  nand2_1 U11704 ( .ip1(n9863), .ip2(n12675), .op(n5994) );
  nor2_1 U11705 ( .ip1(n11285), .ip2(n9862), .op(n9857) );
  inv_1 U11706 ( .ip(n5994), .op(n9856) );
  not_ab_or_c_or_d U11707 ( .ip1(n12679), .ip2(n11447), .ip3(n9857), .ip4(
        n9856), .op(\CORTEXM0DS_INST/u_logic/N4005 ) );
  nand2_1 U11708 ( .ip1(n9863), .ip2(n12681), .op(n5992) );
  inv_1 U11709 ( .ip(n9862), .op(n9861) );
  inv_1 U11710 ( .ip(n9858), .op(n12665) );
  inv_1 U11711 ( .ip(n12679), .op(n12680) );
  nor2_1 U11712 ( .ip1(n11624), .ip2(n12680), .op(n9860) );
  inv_1 U11713 ( .ip(n5992), .op(n9859) );
  not_ab_or_c_or_d U11714 ( .ip1(n9861), .ip2(n12665), .ip3(n9860), .ip4(n9859), .op(\CORTEXM0DS_INST/u_logic/N3967 ) );
  nand2_1 U11715 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(n12673), .op(
        \CORTEXM0DS_INST/u_logic/N3966 ) );
  nand2_1 U11716 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(n12677), .op(
        \CORTEXM0DS_INST/u_logic/N3946 ) );
  nor2_1 U11717 ( .ip1(n11295), .ip2(n9862), .op(n9866) );
  inv_1 U11718 ( .ip(n9863), .op(n12664) );
  nor2_1 U11719 ( .ip1(n9864), .ip2(n12664), .op(n9865) );
  not_ab_or_c_or_d U11720 ( .ip1(n12679), .ip2(n11456), .ip3(n9866), .ip4(
        n9865), .op(\CORTEXM0DS_INST/u_logic/N3783 ) );
  inv_1 U11721 ( .ip(n10859), .op(n10562) );
  nor4_1 U11722 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip3(n11038), .ip4(n12095), .op(
        n9868) );
  not_ab_or_c_or_d U11723 ( .ip1(n9869), .ip2(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip3(n9868), .ip4(n9867), .op(n9870) );
  or2_1 U11724 ( .ip1(n9871), .ip2(n9870), .op(n10046) );
  nor4_1 U11725 ( .ip1(n10053), .ip2(n10052), .ip3(n9872), .ip4(n10046), .op(
        n9875) );
  nor2_1 U11726 ( .ip1(n9874), .ip2(n9873), .op(n10561) );
  inv_1 U11727 ( .ip(n10561), .op(n10426) );
  nand2_1 U11728 ( .ip1(n9875), .ip2(n10426), .op(n11306) );
  nor2_1 U11729 ( .ip1(n10562), .ip2(n11306), .op(n9876) );
  nor2_1 U11730 ( .ip1(n10858), .ip2(n9876), .op(n10240) );
  inv_1 U11731 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [12]), .op(n11668) );
  nor2_1 U11732 ( .ip1(n11668), .ip2(n11841), .op(n9878) );
  and2_1 U11733 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [12]), .ip2(n11787), 
        .op(n9877) );
  not_ab_or_c_or_d U11734 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [12]), .ip2(
        n11610), .ip3(n9878), .ip4(n9877), .op(n9919) );
  inv_1 U11735 ( .ip(n10146), .op(n9909) );
  inv_1 U11736 ( .ip(n9879), .op(n9908) );
  nor2_1 U11737 ( .ip1(n9880), .ip2(n9883), .op(n9881) );
  not_ab_or_c_or_d U11738 ( .ip1(n9883), .ip2(n9882), .ip3(n10138), .ip4(n9881), .op(n9885) );
  not_ab_or_c_or_d U11739 ( .ip1(n9887), .ip2(n9886), .ip3(n9885), .ip4(n9884), 
        .op(n9906) );
  nand3_1 U11740 ( .ip1(n9889), .ip2(n10138), .ip3(n9888), .op(n9905) );
  nand3_1 U11741 ( .ip1(n9891), .ip2(n9895), .ip3(n9890), .op(n9899) );
  inv_1 U11742 ( .ip(n9895), .op(n10136) );
  nand3_1 U11743 ( .ip1(n9893), .ip2(n9892), .ip3(n10136), .op(n9898) );
  nand3_1 U11744 ( .ip1(n9896), .ip2(n9895), .ip3(n9894), .op(n9897) );
  nand3_1 U11745 ( .ip1(n9899), .ip2(n9898), .ip3(n9897), .op(n9900) );
  not_ab_or_c_or_d U11746 ( .ip1(n9902), .ip2(n9901), .ip3(n10140), .ip4(n9900), .op(n9904) );
  inv_1 U11747 ( .ip(n9903), .op(n12439) );
  not_ab_or_c_or_d U11748 ( .ip1(n9906), .ip2(n9905), .ip3(n9904), .ip4(n12439), .op(n9907) );
  not_ab_or_c_or_d U11749 ( .ip1(n9910), .ip2(n9909), .ip3(n9908), .ip4(n9907), 
        .op(n9911) );
  nor2_1 U11750 ( .ip1(\CORTEXM0DS_INST/u_logic/Krgvx4 ), .ip2(n9911), .op(
        n9912) );
  nor2_1 U11751 ( .ip1(\CORTEXM0DS_INST/u_logic/Eqgvx4 ), .ip2(n9912), .op(
        n12457) );
  nor2_1 U11752 ( .ip1(n9913), .ip2(n10148), .op(n9916) );
  nor2_1 U11753 ( .ip1(n9914), .ip2(n11614), .op(n9915) );
  not_ab_or_c_or_d U11754 ( .ip1(n10152), .ip2(n12457), .ip3(n9916), .ip4(
        n9915), .op(n9918) );
  nand2_1 U11755 ( .ip1(n11609), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [12]), 
        .op(n9917) );
  nand4_1 U11756 ( .ip1(n4087), .ip2(n9919), .ip3(n9918), .ip4(n9917), .op(
        n10366) );
  nor2_1 U11757 ( .ip1(n10052), .ip2(n10054), .op(n10397) );
  inv_1 U11758 ( .ip(n10397), .op(n10257) );
  inv_1 U11759 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [4]), .op(n11642) );
  nor2_1 U11760 ( .ip1(n11642), .ip2(n11841), .op(n9927) );
  nand2_1 U11761 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [4]), .ip2(n11610), 
        .op(n9925) );
  nor2_1 U11762 ( .ip1(n12685), .ip2(n9976), .op(n10088) );
  nor3_1 U11763 ( .ip1(n9921), .ip2(n9920), .ip3(n11811), .op(n9923) );
  nor2_1 U11764 ( .ip1(n11810), .ip2(n11896), .op(n9922) );
  not_ab_or_c_or_d U11765 ( .ip1(n10088), .ip2(
        \CORTEXM0DS_INST/u_logic/Vogvx4 ), .ip3(n9923), .ip4(n9922), .op(n9924) );
  nand3_1 U11766 ( .ip1(n9925), .ip2(n9924), .ip3(n4097), .op(n9926) );
  not_ab_or_c_or_d U11767 ( .ip1(n11787), .ip2(
        \CORTEXM0DS_INST/u_logic/L0i2z4 [4]), .ip3(n9927), .ip4(n9926), .op(
        n10367) );
  nor2_1 U11768 ( .ip1(n10367), .ip2(n10426), .op(n9929) );
  nor2_1 U11769 ( .ip1(n4348), .ip2(n10395), .op(n9928) );
  not_ab_or_c_or_d U11770 ( .ip1(n10366), .ip2(n10257), .ip3(n9929), .ip4(
        n9928), .op(n9936) );
  nand2_1 U11771 ( .ip1(\CORTEXM0DS_INST/u_logic/Qsgvx4 ), .ip2(n10152), .op(
        n9932) );
  nand2_1 U11772 ( .ip1(n9930), .ip2(n11821), .op(n9931) );
  nand4_1 U11773 ( .ip1(n4092), .ip2(n10267), .ip3(n9932), .ip4(n9931), .op(
        n10370) );
  nor3_1 U11774 ( .ip1(n9934), .ip2(n9933), .ip3(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .op(n10051) );
  nor2_1 U11775 ( .ip1(n10051), .ip2(n10053), .op(n10400) );
  inv_1 U11776 ( .ip(n10400), .op(n10256) );
  nand2_1 U11777 ( .ip1(n10370), .ip2(n10256), .op(n9935) );
  nand2_1 U11778 ( .ip1(n9936), .ip2(n9935), .op(n11354) );
  nor2_1 U11779 ( .ip1(n9937), .ip2(n10335), .op(n10285) );
  nand2_1 U11780 ( .ip1(\CORTEXM0DS_INST/vis_pc [13]), .ip2(n10285), .op(n9947) );
  nor2_1 U11781 ( .ip1(n10965), .ip2(n9947), .op(n10250) );
  nand2_1 U11782 ( .ip1(\CORTEXM0DS_INST/vis_pc [15]), .ip2(n10250), .op(
        n10251) );
  nor3_1 U11783 ( .ip1(n5822), .ip2(n12166), .ip3(n10251), .op(n10245) );
  nand3_1 U11784 ( .ip1(\CORTEXM0DS_INST/vis_pc [17]), .ip2(
        \CORTEXM0DS_INST/vis_pc [18]), .ip3(n10245), .op(n9939) );
  inv_1 U11785 ( .ip(n9939), .op(n10406) );
  nand2_1 U11786 ( .ip1(\CORTEXM0DS_INST/vis_pc [19]), .ip2(n10406), .op(n9964) );
  inv_1 U11787 ( .ip(n9964), .op(n9938) );
  inv_1 U11788 ( .ip(n12091), .op(n10565) );
  not_ab_or_c_or_d U11789 ( .ip1(n12196), .ip2(n9939), .ip3(n9938), .ip4(
        n10565), .op(n9941) );
  inv_1 U11790 ( .ip(n10572), .op(n10855) );
  nor2_1 U11791 ( .ip1(n12198), .ip2(n10855), .op(n9940) );
  not_ab_or_c_or_d U11792 ( .ip1(n10859), .ip2(n11354), .ip3(n9941), .ip4(
        n9940), .op(n9942) );
  nand2_1 U11793 ( .ip1(n10240), .ip2(n9942), .op(
        \CORTEXM0DS_INST/u_logic/Ldhvx4 ) );
  inv_1 U11794 ( .ip(n9943), .op(n11535) );
  inv_1 U11795 ( .ip(n10310), .op(n10331) );
  inv_1 U11796 ( .ip(n10322), .op(n10311) );
  nor2_1 U11797 ( .ip1(n4130), .ip2(n10311), .op(n9945) );
  nor2_1 U11798 ( .ip1(n4150), .ip2(n10296), .op(n9944) );
  ab_or_c_or_d U11799 ( .ip1(n10416), .ip2(n10331), .ip3(n9945), .ip4(n9944), 
        .op(n9946) );
  not_ab_or_c_or_d U11800 ( .ip1(n10414), .ip2(n10323), .ip3(n10330), .ip4(
        n9946), .op(n11550) );
  nor2_1 U11801 ( .ip1(n11550), .ip2(n10562), .op(n9950) );
  nor2_1 U11802 ( .ip1(n5822), .ip2(n9947), .op(n10286) );
  nor2_1 U11803 ( .ip1(\CORTEXM0DS_INST/vis_pc [14]), .ip2(n10286), .op(n9948)
         );
  not_ab_or_c_or_d U11804 ( .ip1(n10250), .ip2(n10860), .ip3(n9948), .ip4(
        n10565), .op(n9949) );
  not_ab_or_c_or_d U11805 ( .ip1(n10572), .ip2(n11535), .ip3(n9950), .ip4(
        n9949), .op(n9951) );
  nand2_1 U11806 ( .ip1(n9951), .ip2(n10573), .op(
        \CORTEXM0DS_INST/u_logic/Sdhvx4 ) );
  nor2_1 U11807 ( .ip1(n4130), .ip2(n10400), .op(n9956) );
  nor2_1 U11808 ( .ip1(n9952), .ip2(n10395), .op(n9955) );
  nor2_1 U11809 ( .ip1(n4150), .ip2(n10426), .op(n9954) );
  and2_1 U11810 ( .ip1(n10414), .ip2(n10257), .op(n9953) );
  nor4_1 U11811 ( .ip1(n9956), .ip2(n9955), .ip3(n9954), .ip4(n9953), .op(
        n11532) );
  nor2_1 U11812 ( .ip1(n11532), .ip2(n10562), .op(n9959) );
  inv_1 U11813 ( .ip(\CORTEXM0DS_INST/vis_pc [22]), .op(n12101) );
  inv_1 U11814 ( .ip(\CORTEXM0DS_INST/vis_pc [20]), .op(n12207) );
  nor2_1 U11815 ( .ip1(n12207), .ip2(n9964), .op(n10223) );
  nand2_1 U11816 ( .ip1(\CORTEXM0DS_INST/vis_pc [21]), .ip2(n10223), .op(
        n10224) );
  nor2_1 U11817 ( .ip1(n12101), .ip2(n10224), .op(n10432) );
  not_ab_or_c_or_d U11818 ( .ip1(n12101), .ip2(n10224), .ip3(n10432), .ip4(
        n10565), .op(n9958) );
  nor2_1 U11819 ( .ip1(n12103), .ip2(n10855), .op(n9957) );
  inv_1 U11820 ( .ip(n10240), .op(n10408) );
  or4_1 U11821 ( .ip1(n9959), .ip2(n9958), .ip3(n9957), .ip4(n10408), .op(
        \CORTEXM0DS_INST/u_logic/Zdhvx4 ) );
  nor2_1 U11822 ( .ip1(n10357), .ip2(n10395), .op(n9961) );
  nor2_1 U11823 ( .ip1(n10356), .ip2(n10426), .op(n9960) );
  not_ab_or_c_or_d U11824 ( .ip1(n10362), .ip2(n10257), .ip3(n9961), .ip4(
        n9960), .op(n9963) );
  nand2_1 U11825 ( .ip1(n10360), .ip2(n10256), .op(n9962) );
  nand2_1 U11826 ( .ip1(n9963), .ip2(n9962), .op(n11374) );
  not_ab_or_c_or_d U11827 ( .ip1(n12207), .ip2(n9964), .ip3(n10223), .ip4(
        n10565), .op(n9966) );
  nor2_1 U11828 ( .ip1(n12209), .ip2(n10855), .op(n9965) );
  not_ab_or_c_or_d U11829 ( .ip1(n10859), .ip2(n11374), .ip3(n9966), .ip4(
        n9965), .op(n9967) );
  nand2_1 U11830 ( .ip1(n10240), .ip2(n9967), .op(
        \CORTEXM0DS_INST/u_logic/Gehvx4 ) );
  inv_1 U11831 ( .ip(n10396), .op(n10077) );
  nand2_1 U11832 ( .ip1(n10077), .ip2(n10323), .op(n9971) );
  nor2_1 U11833 ( .ip1(n10296), .ip2(n10398), .op(n9969) );
  nor2_1 U11834 ( .ip1(n10311), .ip2(n10399), .op(n9968) );
  not_ab_or_c_or_d U11835 ( .ip1(n10331), .ip2(n10079), .ip3(n9969), .ip4(
        n9968), .op(n9970) );
  nand3_1 U11836 ( .ip1(n9971), .ip2(n9970), .ip3(n10314), .op(n11265) );
  nand2_1 U11837 ( .ip1(n10859), .ip2(n11265), .op(n9975) );
  inv_1 U11838 ( .ip(\CORTEXM0DS_INST/vis_pc [9]), .op(n12122) );
  nor3_1 U11839 ( .ip1(n12113), .ip2(n10335), .ip3(n10861), .op(n10320) );
  nand2_1 U11840 ( .ip1(\CORTEXM0DS_INST/vis_pc [8]), .ip2(n10320), .op(n10308) );
  nor2_1 U11841 ( .ip1(n12122), .ip2(n10308), .op(n10307) );
  and2_1 U11842 ( .ip1(n12137), .ip2(n10572), .op(n9973) );
  nor3_1 U11843 ( .ip1(n10307), .ip2(n10565), .ip3(n12133), .op(n9972) );
  not_ab_or_c_or_d U11844 ( .ip1(n10307), .ip2(n12133), .ip3(n9973), .ip4(
        n9972), .op(n9974) );
  nand3_1 U11845 ( .ip1(n9975), .ip2(n9974), .ip3(n10573), .op(
        \CORTEXM0DS_INST/u_logic/Uehvx4 ) );
  nor2_1 U11846 ( .ip1(n10207), .ip2(n9976), .op(n4241) );
  not_ab_or_c_or_d U11847 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [9]), .ip2(
        n10265), .ip3(n4241), .ip4(n9977), .op(n9986) );
  nand2_1 U11848 ( .ip1(n10184), .ip2(n9978), .op(n9981) );
  nand2_1 U11849 ( .ip1(n11609), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [9]), 
        .op(n9980) );
  nand2_1 U11850 ( .ip1(n11610), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [9]), 
        .op(n9979) );
  and4_1 U11851 ( .ip1(n3197), .ip2(n9981), .ip3(n9980), .ip4(n9979), .op(
        n9985) );
  nand2_1 U11852 ( .ip1(n11607), .ip2(n9982), .op(n9984) );
  nand2_1 U11853 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [9]), .ip2(n11787), 
        .op(n9983) );
  nand4_1 U11854 ( .ip1(n9986), .ip2(n9985), .ip3(n9984), .ip4(n9983), .op(
        n10848) );
  nand2_1 U11855 ( .ip1(n10848), .ip2(n10323), .op(n10011) );
  inv_1 U11856 ( .ip(n10296), .op(n10325) );
  nor2_1 U11857 ( .ip1(n9987), .ip2(n10148), .op(n9993) );
  nand2_1 U11858 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [1]), .ip2(n11787), 
        .op(n9991) );
  nand2_1 U11859 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [1]), .ip2(n10265), 
        .op(n9990) );
  nand2_1 U11860 ( .ip1(n11610), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [1]), 
        .op(n9989) );
  nand3_1 U11861 ( .ip1(n12683), .ip2(n11807), .ip3(n11867), .op(n10091) );
  inv_1 U11862 ( .ip(n10091), .op(n10272) );
  nand2_1 U11863 ( .ip1(n10272), .ip2(\CORTEXM0DS_INST/u_logic/S0hvx4 ), .op(
        n9988) );
  nand4_1 U11864 ( .ip1(n9991), .ip2(n9990), .ip3(n9989), .ip4(n9988), .op(
        n9992) );
  not_ab_or_c_or_d U11865 ( .ip1(n10184), .ip2(n9994), .ip3(n9993), .ip4(n9992), .op(n9997) );
  nand2_1 U11866 ( .ip1(n11609), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [1]), 
        .op(n9996) );
  nand2_1 U11867 ( .ip1(\CORTEXM0DS_INST/u_logic/Eg8vx4 ), .ip2(n10088), .op(
        n9995) );
  nand4_1 U11868 ( .ip1(n3178), .ip2(n9997), .ip3(n9996), .ip4(n9995), .op(
        n10844) );
  and2_1 U11869 ( .ip1(n9998), .ip2(n11607), .op(n10003) );
  nand2_1 U11870 ( .ip1(n10184), .ip2(n9999), .op(n10001) );
  nand2_1 U11871 ( .ip1(n11609), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [17]), 
        .op(n10000) );
  nand3_1 U11872 ( .ip1(n10001), .ip2(n3204), .ip3(n10000), .op(n10002) );
  not_ab_or_c_or_d U11873 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [17]), .ip2(
        n11610), .ip3(n10003), .ip4(n10002), .op(n10845) );
  nor2_1 U11874 ( .ip1(n10310), .ip2(n10845), .op(n10004) );
  not_ab_or_c_or_d U11875 ( .ip1(n10325), .ip2(n10844), .ip3(n10330), .ip4(
        n10004), .op(n10010) );
  nand2_1 U11876 ( .ip1(n10109), .ip2(n10005), .op(n10008) );
  nand2_1 U11877 ( .ip1(n10006), .ip2(n11821), .op(n10007) );
  nand4_1 U11878 ( .ip1(n3164), .ip2(n10267), .ip3(n10008), .ip4(n10007), .op(
        n10850) );
  nand2_1 U11879 ( .ip1(n10322), .ip2(n10850), .op(n10009) );
  nand3_1 U11880 ( .ip1(n10011), .ip2(n10010), .ip3(n10009), .op(n11719) );
  nor2_1 U11881 ( .ip1(n10012), .ip2(n10855), .op(n10015) );
  nor2_1 U11882 ( .ip1(n10320), .ip2(n10565), .op(n10013) );
  mux2_1 U11883 ( .ip1(n10320), .ip2(n10013), .s(\CORTEXM0DS_INST/vis_pc [8]), 
        .op(n10014) );
  not_ab_or_c_or_d U11884 ( .ip1(n10859), .ip2(n11719), .ip3(n10015), .ip4(
        n10014), .op(n10016) );
  nand2_1 U11885 ( .ip1(n10016), .ip2(n10573), .op(
        \CORTEXM0DS_INST/u_logic/Bfhvx4 ) );
  nand2_1 U11886 ( .ip1(n12329), .ip2(n12588), .op(n10018) );
  nand2_1 U11887 ( .ip1(n12328), .ip2(n11032), .op(n12055) );
  mux2_1 U11888 ( .ip1(n10033), .ip2(n12055), .s(n10457), .op(n11044) );
  inv_1 U11889 ( .ip(n11044), .op(n10017) );
  not_ab_or_c_or_d U11890 ( .ip1(n11135), .ip2(n10018), .ip3(n10807), .ip4(
        n10017), .op(n10034) );
  or2_1 U11891 ( .ip1(n10034), .ip2(n12570), .op(n10021) );
  nand3_1 U11892 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n11032), .ip3(
        n11068), .op(n10019) );
  or2_1 U11893 ( .ip1(n10019), .ip2(n12570), .op(n10020) );
  nand2_1 U11894 ( .ip1(n10021), .ip2(n10020), .op(n10022) );
  or2_1 U11895 ( .ip1(\CORTEXM0DS_INST/u_logic/K79vx4 ), .ip2(n10022), .op(
        n10024) );
  nor2_1 U11896 ( .ip1(n12075), .ip2(n11070), .op(n10918) );
  nor2_1 U11897 ( .ip1(n10918), .ip2(n12381), .op(n12035) );
  inv_1 U11898 ( .ip(n12035), .op(n12064) );
  or2_1 U11899 ( .ip1(n12064), .ip2(n10022), .op(n10023) );
  nand2_1 U11900 ( .ip1(n10024), .ip2(n10023), .op(n10026) );
  inv_1 U11901 ( .ip(\CORTEXM0DS_INST/u_logic/Ks9vx4 ), .op(n10025) );
  mux2_1 U11902 ( .ip1(n10026), .ip2(n10025), .s(n5780), .op(n10032) );
  nand2_1 U11903 ( .ip1(n10027), .ip2(n6210), .op(n10549) );
  nand2_1 U11904 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10661), .op(
        n10028) );
  nand2_1 U11905 ( .ip1(n10549), .ip2(n10028), .op(n11075) );
  not_ab_or_c_or_d U11906 ( .ip1(n11725), .ip2(n10727), .ip3(n10029), .ip4(
        n11075), .op(n12043) );
  inv_1 U11907 ( .ip(n12043), .op(n12067) );
  nand3_1 U11908 ( .ip1(\CORTEXM0DS_INST/u_logic/Ks9vx4 ), .ip2(n10030), .ip3(
        n12067), .op(n10031) );
  nand2_1 U11909 ( .ip1(n10032), .ip2(n10031), .op(
        \CORTEXM0DS_INST/u_logic/Wfhvx4 ) );
  nor2_1 U11910 ( .ip1(n12035), .ip2(n12558), .op(n10035) );
  or2_1 U11911 ( .ip1(\CORTEXM0DS_INST/u_logic/K79vx4 ), .ip2(n10035), .op(
        n10037) );
  nand2_1 U11912 ( .ip1(n10034), .ip2(n10033), .op(n12052) );
  or2_1 U11913 ( .ip1(n12052), .ip2(n10035), .op(n10036) );
  nand2_1 U11914 ( .ip1(n10037), .ip2(n10036), .op(n10039) );
  mux2_1 U11915 ( .ip1(n10039), .ip2(n10038), .s(n5780), .op(n10042) );
  nand3_1 U11916 ( .ip1(\CORTEXM0DS_INST/u_logic/Gr9vx4 ), .ip2(n10040), .ip3(
        n12067), .op(n10041) );
  nand2_1 U11917 ( .ip1(n10042), .ip2(n10041), .op(
        \CORTEXM0DS_INST/u_logic/Dghvx4 ) );
  nor2_1 U11918 ( .ip1(n10044), .ip2(n10043), .op(n10045) );
  nor2_1 U11919 ( .ip1(n10046), .ip2(n10045), .op(n10559) );
  nor2_1 U11920 ( .ip1(n10048), .ip2(n10047), .op(n10049) );
  nor2_1 U11921 ( .ip1(n10050), .ip2(n10049), .op(n10553) );
  inv_1 U11922 ( .ip(n10553), .op(n10423) );
  nor2_1 U11923 ( .ip1(n10052), .ip2(n10051), .op(n10127) );
  nor2_1 U11924 ( .ip1(n10127), .ip2(n10357), .op(n10059) );
  or2_1 U11925 ( .ip1(n10053), .ip2(n10054), .op(n10057) );
  or2_1 U11926 ( .ip1(n10055), .ip2(n10054), .op(n10056) );
  nand2_1 U11927 ( .ip1(n10057), .ip2(n10056), .op(n10551) );
  nor2_1 U11928 ( .ip1(n10551), .ip2(n10356), .op(n10058) );
  ab_or_c_or_d U11929 ( .ip1(n10423), .ip2(n10360), .ip3(n10059), .ip4(n10058), 
        .op(n10060) );
  not_ab_or_c_or_d U11930 ( .ip1(n10561), .ip2(n10362), .ip3(n10559), .ip4(
        n10060), .op(n11779) );
  nor2_1 U11931 ( .ip1(n11779), .ip2(n10562), .op(n10062) );
  inv_1 U11932 ( .ip(\CORTEXM0DS_INST/vis_pc [24]), .op(n12248) );
  nand2_1 U11933 ( .ip1(\CORTEXM0DS_INST/vis_pc [23]), .ip2(n10432), .op(
        n10433) );
  nor3_1 U11934 ( .ip1(n12248), .ip2(n12257), .ip3(n10433), .op(n10120) );
  nand3_1 U11935 ( .ip1(\CORTEXM0DS_INST/vis_pc [27]), .ip2(
        \CORTEXM0DS_INST/vis_pc [26]), .ip3(n10120), .op(n10563) );
  nor3_1 U11936 ( .ip1(\CORTEXM0DS_INST/vis_pc [28]), .ip2(n10565), .ip3(
        n10563), .op(n10061) );
  not_ab_or_c_or_d U11937 ( .ip1(n10572), .ip2(n10063), .ip3(n10062), .ip4(
        n10061), .op(n10065) );
  nand3_1 U11938 ( .ip1(n12091), .ip2(\CORTEXM0DS_INST/vis_pc [28]), .ip3(
        n10563), .op(n10064) );
  nand3_1 U11939 ( .ip1(n10065), .ip2(n10573), .ip3(n10064), .op(
        \CORTEXM0DS_INST/u_logic/Mhhvx4 ) );
  nor2_1 U11940 ( .ip1(n10127), .ip2(n4348), .op(n10067) );
  nor2_1 U11941 ( .ip1(n10551), .ip2(n10367), .op(n10066) );
  ab_or_c_or_d U11942 ( .ip1(n10423), .ip2(n10370), .ip3(n10067), .ip4(n10066), 
        .op(n10068) );
  not_ab_or_c_or_d U11943 ( .ip1(n10561), .ip2(n10366), .ip3(n10559), .ip4(
        n10068), .op(n11467) );
  nor2_1 U11944 ( .ip1(n11467), .ip2(n10562), .op(n10070) );
  and3_1 U11945 ( .ip1(n12091), .ip2(\CORTEXM0DS_INST/vis_pc [27]), .ip3(
        n10563), .op(n10069) );
  not_ab_or_c_or_d U11946 ( .ip1(n10572), .ip2(n10071), .ip3(n10070), .ip4(
        n10069), .op(n10074) );
  nand4_1 U11947 ( .ip1(\CORTEXM0DS_INST/vis_pc [26]), .ip2(n12091), .ip3(
        n10120), .ip4(n10072), .op(n10073) );
  nand3_1 U11948 ( .ip1(n10074), .ip2(n10573), .ip3(n10073), .op(
        \CORTEXM0DS_INST/u_logic/Thhvx4 ) );
  inv_1 U11949 ( .ip(n10127), .op(n10557) );
  nor2_1 U11950 ( .ip1(n10553), .ip2(n10399), .op(n10076) );
  nor2_1 U11951 ( .ip1(n10551), .ip2(n10398), .op(n10075) );
  ab_or_c_or_d U11952 ( .ip1(n10561), .ip2(n10077), .ip3(n10076), .ip4(n10075), 
        .op(n10078) );
  not_ab_or_c_or_d U11953 ( .ip1(n10557), .ip2(n10079), .ip3(n10559), .ip4(
        n10078), .op(n11445) );
  nor2_1 U11954 ( .ip1(n11445), .ip2(n10562), .op(n10083) );
  nor2_1 U11955 ( .ip1(n12271), .ip2(n10855), .op(n10082) );
  nor2_1 U11956 ( .ip1(n10120), .ip2(\CORTEXM0DS_INST/vis_pc [26]), .op(n10080) );
  not_ab_or_c_or_d U11957 ( .ip1(n10120), .ip2(\CORTEXM0DS_INST/vis_pc [26]), 
        .ip3(n10080), .ip4(n10565), .op(n10081) );
  or4_1 U11958 ( .ip1(n10858), .ip2(n10083), .ip3(n10082), .ip4(n10081), .op(
        \CORTEXM0DS_INST/u_logic/Aihvx4 ) );
  inv_1 U11959 ( .ip(n10551), .op(n10126) );
  nand2_1 U11960 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [2]), .ip2(n11787), 
        .op(n10087) );
  nand2_1 U11961 ( .ip1(n11609), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [2]), 
        .op(n10086) );
  nand2_1 U11962 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [2]), .ip2(n10265), 
        .op(n10085) );
  nand2_1 U11963 ( .ip1(n11610), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [2]), 
        .op(n10084) );
  nand4_1 U11964 ( .ip1(n10087), .ip2(n10086), .ip3(n10085), .ip4(n10084), 
        .op(n10093) );
  nand2_1 U11965 ( .ip1(n10184), .ip2(n10185), .op(n10090) );
  nand2_1 U11966 ( .ip1(n10088), .ip2(\CORTEXM0DS_INST/u_logic/Nngvx4 ), .op(
        n10089) );
  nand4_1 U11967 ( .ip1(n4263), .ip2(n10091), .ip3(n10090), .ip4(n10089), .op(
        n10092) );
  not_ab_or_c_or_d U11968 ( .ip1(n11607), .ip2(n10094), .ip3(n10093), .ip4(
        n10092), .op(n10231) );
  inv_1 U11969 ( .ip(n10231), .op(n10389) );
  inv_1 U11970 ( .ip(n10095), .op(n10149) );
  nor2_1 U11971 ( .ip1(n10149), .ip2(n11614), .op(n10103) );
  inv_1 U11972 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [10]), .op(n11677) );
  nor2_1 U11973 ( .ip1(n11677), .ip2(n11841), .op(n10096) );
  or2_1 U11974 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [10]), .ip2(n10096), 
        .op(n10098) );
  or2_1 U11975 ( .ip1(n11610), .ip2(n10096), .op(n10097) );
  nand2_1 U11976 ( .ip1(n10098), .ip2(n10097), .op(n10101) );
  nand2_1 U11977 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [10]), .ip2(n11787), 
        .op(n10100) );
  nand2_1 U11978 ( .ip1(n11609), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [10]), 
        .op(n10099) );
  nand4_1 U11979 ( .ip1(n4237), .ip2(n10101), .ip3(n10100), .ip4(n10099), .op(
        n10102) );
  not_ab_or_c_or_d U11980 ( .ip1(n11607), .ip2(n10183), .ip3(n10103), .ip4(
        n10102), .op(n10230) );
  inv_1 U11981 ( .ip(n10230), .op(n10387) );
  nor2_1 U11982 ( .ip1(n11690), .ip2(n10266), .op(n10107) );
  nand2_1 U11983 ( .ip1(n10104), .ip2(n11821), .op(n10105) );
  nand2_1 U11984 ( .ip1(n4227), .ip2(n10105), .op(n10106) );
  not_ab_or_c_or_d U11985 ( .ip1(n10109), .ip2(n10108), .ip3(n10107), .ip4(
        n10106), .op(n10384) );
  nor2_1 U11986 ( .ip1(n10553), .ip2(n10384), .op(n10118) );
  inv_1 U11987 ( .ip(n10110), .op(n10147) );
  nor2_1 U11988 ( .ip1(n10147), .ip2(n10148), .op(n10111) );
  not_ab_or_c_or_d U11989 ( .ip1(n11610), .ip2(
        \CORTEXM0DS_INST/u_logic/Czh2z4 [18]), .ip3(n10111), .ip4(n4241), .op(
        n10113) );
  nand2_1 U11990 ( .ip1(n11609), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [18]), 
        .op(n10112) );
  nand4_1 U11991 ( .ip1(n4243), .ip2(n10113), .ip3(n10267), .ip4(n10112), .op(
        n10114) );
  or2_1 U11992 ( .ip1(n10184), .ip2(n10114), .op(n10116) );
  or2_1 U11993 ( .ip1(n10219), .ip2(n10114), .op(n10115) );
  nand2_1 U11994 ( .ip1(n10116), .ip2(n10115), .op(n10383) );
  nor2_1 U11995 ( .ip1(n10127), .ip2(n10383), .op(n10117) );
  ab_or_c_or_d U11996 ( .ip1(n10561), .ip2(n10387), .ip3(n10118), .ip4(n10117), 
        .op(n10119) );
  not_ab_or_c_or_d U11997 ( .ip1(n10126), .ip2(n10389), .ip3(n10559), .ip4(
        n10119), .op(n11440) );
  nor2_1 U11998 ( .ip1(n11440), .ip2(n10562), .op(n10123) );
  nor2_1 U11999 ( .ip1(n10565), .ip2(n10433), .op(n10125) );
  nand2_1 U12000 ( .ip1(\CORTEXM0DS_INST/vis_pc [24]), .ip2(n10125), .op(
        n10121) );
  not_ab_or_c_or_d U12001 ( .ip1(n12257), .ip2(n10121), .ip3(n10120), .ip4(
        n10565), .op(n10122) );
  not_ab_or_c_or_d U12002 ( .ip1(n10572), .ip2(n12262), .ip3(n10123), .ip4(
        n10122), .op(n10124) );
  nand2_1 U12003 ( .ip1(n10124), .ip2(n10573), .op(
        \CORTEXM0DS_INST/u_logic/Hihvx4 ) );
  nand2_1 U12004 ( .ip1(n10125), .ip2(n12248), .op(n10135) );
  nand2_1 U12005 ( .ip1(n10844), .ip2(n10126), .op(n10131) );
  nor2_1 U12006 ( .ip1(n10127), .ip2(n10845), .op(n10128) );
  not_ab_or_c_or_d U12007 ( .ip1(n10561), .ip2(n10848), .ip3(n10559), .ip4(
        n10128), .op(n10130) );
  nand2_1 U12008 ( .ip1(n10423), .ip2(n10850), .op(n10129) );
  nand3_1 U12009 ( .ip1(n10131), .ip2(n10130), .ip3(n10129), .op(n11419) );
  nor2_1 U12010 ( .ip1(n12250), .ip2(n10855), .op(n10132) );
  not_ab_or_c_or_d U12011 ( .ip1(n10859), .ip2(n11419), .ip3(n10858), .ip4(
        n10132), .op(n10134) );
  nand3_1 U12012 ( .ip1(n12091), .ip2(\CORTEXM0DS_INST/vis_pc [24]), .ip3(
        n10433), .op(n10133) );
  nand3_1 U12013 ( .ip1(n10135), .ip2(n10134), .ip3(n10133), .op(
        \CORTEXM0DS_INST/u_logic/Oihvx4 ) );
  nor2_1 U12014 ( .ip1(n10137), .ip2(n10136), .op(n10139) );
  or2_1 U12015 ( .ip1(n10138), .ip2(n10139), .op(n10142) );
  or2_1 U12016 ( .ip1(n10140), .ip2(n10139), .op(n10141) );
  nand2_1 U12017 ( .ip1(n10142), .ip2(n10141), .op(n10143) );
  nor2_1 U12018 ( .ip1(n10143), .ip2(n12439), .op(n10144) );
  not_ab_or_c_or_d U12019 ( .ip1(n10146), .ip2(n10145), .ip3(n10144), .ip4(
        n12440), .op(n12466) );
  nor2_1 U12020 ( .ip1(n10147), .ip2(n11614), .op(n10151) );
  nor2_1 U12021 ( .ip1(n10149), .ip2(n10148), .op(n10150) );
  not_ab_or_c_or_d U12022 ( .ip1(n10152), .ip2(n12466), .ip3(n10151), .ip4(
        n10150), .op(n10165) );
  inv_1 U12023 ( .ip(n4241), .op(n10164) );
  nand2_1 U12024 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [14]), .ip2(n11866), 
        .op(n10161) );
  and2_1 U12025 ( .ip1(n11827), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [18]), 
        .op(n10158) );
  nand2_1 U12026 ( .ip1(n11824), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [2]), 
        .op(n10156) );
  nand2_1 U12027 ( .ip1(n11833), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [10]), 
        .op(n10155) );
  nand2_1 U12028 ( .ip1(n11800), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [14]), 
        .op(n10154) );
  nand2_1 U12029 ( .ip1(n11823), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [26]), 
        .op(n10153) );
  nand4_1 U12030 ( .ip1(n10156), .ip2(n10155), .ip3(n10154), .ip4(n10153), 
        .op(n10157) );
  not_ab_or_c_or_d U12031 ( .ip1(n11799), .ip2(
        \CORTEXM0DS_INST/u_logic/Czh2z4 [14]), .ip3(n10158), .ip4(n10157), 
        .op(n10160) );
  nand2_1 U12032 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [14]), .ip2(n11801), 
        .op(n10159) );
  nand3_1 U12033 ( .ip1(n10161), .ip2(n10160), .ip3(n10159), .op(n10162) );
  nand2_1 U12034 ( .ip1(n11807), .ip2(n10162), .op(n10163) );
  nand4_1 U12035 ( .ip1(n3419), .ip2(n10165), .ip3(n10164), .ip4(n10163), .op(
        n10560) );
  nand2_1 U12036 ( .ip1(n10171), .ip2(n10166), .op(n12636) );
  nor2_1 U12037 ( .ip1(n10167), .ip2(n12636), .op(n10178) );
  nand2_1 U12038 ( .ip1(n11827), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [22]), 
        .op(n10176) );
  nand2_1 U12039 ( .ip1(\CORTEXM0DS_INST/u_logic/Z7hvx4 ), .ip2(n10168), .op(
        n10169) );
  not_ab_or_c_or_d U12040 ( .ip1(\CORTEXM0DS_INST/u_logic/L9hvx4 ), .ip2(
        n10170), .ip3(n10207), .ip4(n10169), .op(n10173) );
  nand4_1 U12041 ( .ip1(\CORTEXM0DS_INST/u_logic/L9hvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Z7hvx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/B5hvx4 ), .ip4(n10171), .op(n10172) );
  nand2_1 U12042 ( .ip1(n12017), .ip2(n10172), .op(n11838) );
  not_ab_or_c_or_d U12043 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [30]), .ip2(
        n11823), .ip3(n10173), .ip4(n11838), .op(n10175) );
  nand2_1 U12044 ( .ip1(n11824), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [6]), 
        .op(n10174) );
  nand3_1 U12045 ( .ip1(n10176), .ip2(n10175), .ip3(n10174), .op(n10177) );
  not_ab_or_c_or_d U12046 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [14]), .ip2(
        n11833), .ip3(n10178), .ip4(n10177), .op(n10179) );
  nor2_1 U12047 ( .ip1(n10179), .ip2(n11839), .op(n10181) );
  inv_1 U12048 ( .ip(n3485), .op(n10180) );
  not_ab_or_c_or_d U12049 ( .ip1(n11821), .ip2(n10182), .ip3(n10181), .ip4(
        n10180), .op(n10552) );
  nor2_1 U12050 ( .ip1(n10552), .ip2(n10400), .op(n10201) );
  nand2_1 U12051 ( .ip1(n10184), .ip2(n10183), .op(n10199) );
  nand2_1 U12052 ( .ip1(n11607), .ip2(n10185), .op(n10198) );
  nand2_1 U12053 ( .ip1(n11833), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [8]), 
        .op(n10195) );
  nor2_1 U12054 ( .ip1(n11790), .ip2(n10186), .op(n10192) );
  nand2_1 U12055 ( .ip1(n11824), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [0]), 
        .op(n10190) );
  nand2_1 U12056 ( .ip1(n11866), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [6]), 
        .op(n10189) );
  nand2_1 U12057 ( .ip1(n11799), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [6]), 
        .op(n10188) );
  nand2_1 U12058 ( .ip1(n11800), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [6]), 
        .op(n10187) );
  nand4_1 U12059 ( .ip1(n10190), .ip2(n10189), .ip3(n10188), .ip4(n10187), 
        .op(n10191) );
  not_ab_or_c_or_d U12060 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [16]), .ip2(
        n11827), .ip3(n10192), .ip4(n10191), .op(n10194) );
  nand2_1 U12061 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [6]), .ip2(n11801), 
        .op(n10193) );
  nand3_1 U12062 ( .ip1(n10195), .ip2(n10194), .ip3(n10193), .op(n10196) );
  nand2_1 U12063 ( .ip1(n11807), .ip2(n10196), .op(n10197) );
  and4_1 U12064 ( .ip1(n3514), .ip2(n10199), .ip3(n10198), .ip4(n10197), .op(
        n10550) );
  nor2_1 U12065 ( .ip1(n10550), .ip2(n10426), .op(n10200) );
  not_ab_or_c_or_d U12066 ( .ip1(n10560), .ip2(n10257), .ip3(n10201), .ip4(
        n10200), .op(n10222) );
  nor2_1 U12067 ( .ip1(n11790), .ip2(n10202), .op(n10214) );
  nand2_1 U12068 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [22]), .ip2(n11866), 
        .op(n10212) );
  inv_1 U12069 ( .ip(n11824), .op(n11814) );
  nor2_1 U12070 ( .ip1(n11814), .ip2(n10203), .op(n10206) );
  nor2_1 U12071 ( .ip1(n11795), .ip2(n10204), .op(n10205) );
  not_ab_or_c_or_d U12072 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [12]), .ip2(
        n11833), .ip3(n10206), .ip4(n10205), .op(n10211) );
  nor4_1 U12073 ( .ip1(\CORTEXM0DS_INST/u_logic/B5hvx4 ), .ip2(n10209), .ip3(
        n10208), .ip4(n10207), .op(n12637) );
  nand2_1 U12074 ( .ip1(\CORTEXM0DS_INST/u_logic/Psh2z4 [0]), .ip2(n12637), 
        .op(n10210) );
  nand3_1 U12075 ( .ip1(n10212), .ip2(n10211), .ip3(n10210), .op(n10213) );
  not_ab_or_c_or_d U12076 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [22]), .ip2(
        n11799), .ip3(n10214), .ip4(n10213), .op(n10215) );
  nor2_1 U12077 ( .ip1(n10215), .ip2(n11839), .op(n10218) );
  nor2_1 U12078 ( .ip1(n10216), .ip2(n11614), .op(n10217) );
  not_ab_or_c_or_d U12079 ( .ip1(n11607), .ip2(n10219), .ip3(n10218), .ip4(
        n10217), .op(n10220) );
  nand2_1 U12080 ( .ip1(n3554), .ip2(n10220), .op(n10556) );
  inv_1 U12081 ( .ip(n10395), .op(n10276) );
  nand2_1 U12082 ( .ip1(n10556), .ip2(n10276), .op(n10221) );
  nand2_1 U12083 ( .ip1(n10222), .ip2(n10221), .op(n11380) );
  inv_1 U12084 ( .ip(n10223), .op(n10226) );
  inv_1 U12085 ( .ip(n10224), .op(n10225) );
  not_ab_or_c_or_d U12086 ( .ip1(n12217), .ip2(n10226), .ip3(n10225), .ip4(
        n10565), .op(n10228) );
  nor2_1 U12087 ( .ip1(n12219), .ip2(n10855), .op(n10227) );
  not_ab_or_c_or_d U12088 ( .ip1(n10859), .ip2(n11380), .ip3(n10228), .ip4(
        n10227), .op(n10229) );
  nand2_1 U12089 ( .ip1(n10240), .ip2(n10229), .op(
        \CORTEXM0DS_INST/u_logic/Vihvx4 ) );
  nor2_1 U12090 ( .ip1(n10400), .ip2(n10384), .op(n10235) );
  nor2_1 U12091 ( .ip1(n10397), .ip2(n10230), .op(n10234) );
  nor2_1 U12092 ( .ip1(n10395), .ip2(n10383), .op(n10233) );
  nor2_1 U12093 ( .ip1(n10231), .ip2(n10426), .op(n10232) );
  nor4_1 U12094 ( .ip1(n10235), .ip2(n10234), .ip3(n10233), .ip4(n10232), .op(
        n11339) );
  nor2_1 U12095 ( .ip1(n11339), .ip2(n10562), .op(n10238) );
  nor3_1 U12096 ( .ip1(n12166), .ip2(n10251), .ip3(n10861), .op(n10405) );
  nor2_1 U12097 ( .ip1(n10245), .ip2(n10565), .op(n10236) );
  mux2_1 U12098 ( .ip1(n10405), .ip2(n10236), .s(\CORTEXM0DS_INST/vis_pc [17]), 
        .op(n10237) );
  not_ab_or_c_or_d U12099 ( .ip1(n10572), .ip2(n12182), .ip3(n10238), .ip4(
        n10237), .op(n10239) );
  nand2_1 U12100 ( .ip1(n10240), .ip2(n10239), .op(
        \CORTEXM0DS_INST/u_logic/Cjhvx4 ) );
  nor2_1 U12101 ( .ip1(n10395), .ip2(n10845), .op(n10244) );
  nand2_1 U12102 ( .ip1(n10848), .ip2(n10257), .op(n10242) );
  nand2_1 U12103 ( .ip1(n10850), .ip2(n10256), .op(n10241) );
  nand2_1 U12104 ( .ip1(n10242), .ip2(n10241), .op(n10243) );
  not_ab_or_c_or_d U12105 ( .ip1(n10561), .ip2(n10844), .ip3(n10244), .ip4(
        n10243), .op(n11329) );
  nor2_1 U12106 ( .ip1(n11329), .ip2(n10562), .op(n10249) );
  inv_1 U12107 ( .ip(n10861), .op(n10284) );
  nand3_1 U12108 ( .ip1(\CORTEXM0DS_INST/vis_pc [15]), .ip2(n10250), .ip3(
        n10284), .op(n10246) );
  not_ab_or_c_or_d U12109 ( .ip1(n12166), .ip2(n10246), .ip3(n10245), .ip4(
        n10565), .op(n10248) );
  nor2_1 U12110 ( .ip1(n12168), .ip2(n10855), .op(n10247) );
  or4_1 U12111 ( .ip1(n10249), .ip2(n10248), .ip3(n10247), .ip4(n10408), .op(
        \CORTEXM0DS_INST/u_logic/Jjhvx4 ) );
  nand2_1 U12112 ( .ip1(n12162), .ip2(n10572), .op(n10283) );
  inv_1 U12113 ( .ip(\CORTEXM0DS_INST/vis_pc [15]), .op(n12157) );
  inv_1 U12114 ( .ip(n10250), .op(n10253) );
  inv_1 U12115 ( .ip(n10251), .op(n10252) );
  not_ab_or_c_or_d U12116 ( .ip1(n12157), .ip2(n10253), .ip3(n10252), .ip4(
        n10861), .op(n10254) );
  not_ab_or_c_or_d U12117 ( .ip1(n5822), .ip2(\CORTEXM0DS_INST/vis_pc [15]), 
        .ip3(n10254), .ip4(n10408), .op(n10282) );
  not_ab_or_c_or_d U12118 ( .ip1(n11821), .ip2(n10255), .ip3(n3979), .ip4(
        n4241), .op(n10995) );
  inv_1 U12119 ( .ip(n10995), .op(n10424) );
  nand2_1 U12120 ( .ip1(n10424), .ip2(n10256), .op(n10280) );
  inv_1 U12121 ( .ip(n4408), .op(n10324) );
  nand2_1 U12122 ( .ip1(n10324), .ip2(n10257), .op(n10279) );
  inv_1 U12123 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [0]), .op(n11879) );
  nor2_1 U12124 ( .ip1(n11810), .ip2(n11879), .op(n10264) );
  nand2_1 U12125 ( .ip1(n11787), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [0]), 
        .op(n10262) );
  nor2_1 U12126 ( .ip1(n10258), .ip2(n11811), .op(n10260) );
  and2_1 U12127 ( .ip1(n10272), .ip2(\CORTEXM0DS_INST/u_logic/F2hvx4 ), .op(
        n10259) );
  not_ab_or_c_or_d U12128 ( .ip1(n11610), .ip2(
        \CORTEXM0DS_INST/u_logic/Czh2z4 [0]), .ip3(n10260), .ip4(n10259), .op(
        n10261) );
  nand3_1 U12129 ( .ip1(n10262), .ip2(n10261), .ip3(n3962), .op(n10263) );
  not_ab_or_c_or_d U12130 ( .ip1(n10265), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [0]), .ip3(n10264), .ip4(n10263), .op(
        n10425) );
  inv_1 U12131 ( .ip(n10425), .op(n11000) );
  nand2_1 U12132 ( .ip1(n10561), .ip2(n11000), .op(n10278) );
  nand2_1 U12133 ( .ip1(n11610), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [16]), 
        .op(n10275) );
  nor3_1 U12134 ( .ip1(n12440), .ip2(n12439), .ip3(n10266), .op(n10270) );
  nand2_1 U12135 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [16]), .ip2(n11609), 
        .op(n10268) );
  nand3_1 U12136 ( .ip1(n10268), .ip2(n3958), .ip3(n10267), .op(n10269) );
  not_ab_or_c_or_d U12137 ( .ip1(n11821), .ip2(n10271), .ip3(n10270), .ip4(
        n10269), .op(n10274) );
  nand2_1 U12138 ( .ip1(\CORTEXM0DS_INST/u_logic/Izgvx4 ), .ip2(n10272), .op(
        n10273) );
  nand3_1 U12139 ( .ip1(n10275), .ip2(n10274), .ip3(n10273), .op(n11004) );
  nand2_1 U12140 ( .ip1(n11004), .ip2(n10276), .op(n10277) );
  nand4_1 U12141 ( .ip1(n10280), .ip2(n10279), .ip3(n10278), .ip4(n10277), 
        .op(n11307) );
  nand2_1 U12142 ( .ip1(n10859), .ip2(n11307), .op(n10281) );
  nand3_1 U12143 ( .ip1(n10283), .ip2(n10282), .ip3(n10281), .op(
        \CORTEXM0DS_INST/u_logic/Qjhvx4 ) );
  nand2_1 U12144 ( .ip1(n10285), .ip2(n10284), .op(n10287) );
  not_ab_or_c_or_d U12145 ( .ip1(n10288), .ip2(n10287), .ip3(n10286), .ip4(
        n10565), .op(n10289) );
  not_ab_or_c_or_d U12146 ( .ip1(n10572), .ip2(n11302), .ip3(n10858), .ip4(
        n10289), .op(n10295) );
  nand2_1 U12147 ( .ip1(n10323), .ip2(n10560), .op(n10293) );
  nor2_1 U12148 ( .ip1(n10550), .ip2(n10296), .op(n10291) );
  nor2_1 U12149 ( .ip1(n10552), .ip2(n10311), .op(n10290) );
  not_ab_or_c_or_d U12150 ( .ip1(n10556), .ip2(n10331), .ip3(n10291), .ip4(
        n10290), .op(n10292) );
  nand3_1 U12151 ( .ip1(n10293), .ip2(n10292), .ip3(n10314), .op(n11300) );
  nand2_1 U12152 ( .ip1(n10859), .ip2(n11300), .op(n10294) );
  nand2_1 U12153 ( .ip1(n10295), .ip2(n10294), .op(
        \CORTEXM0DS_INST/u_logic/Xjhvx4 ) );
  nor2_1 U12154 ( .ip1(n4348), .ip2(n10310), .op(n10298) );
  nor2_1 U12155 ( .ip1(n10367), .ip2(n10296), .op(n10297) );
  ab_or_c_or_d U12156 ( .ip1(n10370), .ip2(n10322), .ip3(n10298), .ip4(n10297), 
        .op(n10299) );
  not_ab_or_c_or_d U12157 ( .ip1(n10366), .ip2(n10323), .ip3(n10330), .ip4(
        n10299), .op(n11282) );
  nor2_1 U12158 ( .ip1(n11282), .ip2(n10562), .op(n10305) );
  or2_1 U12159 ( .ip1(\CORTEXM0DS_INST/vis_pc [10]), .ip2(
        \CORTEXM0DS_INST/vis_pc [11]), .op(n10301) );
  or2_1 U12160 ( .ip1(n10307), .ip2(\CORTEXM0DS_INST/vis_pc [11]), .op(n10300)
         );
  nand2_1 U12161 ( .ip1(n10301), .ip2(n10300), .op(n10303) );
  nor2_1 U12162 ( .ip1(n10303), .ip2(n10302), .op(n10304) );
  not_ab_or_c_or_d U12163 ( .ip1(n10572), .ip2(n12147), .ip3(n10305), .ip4(
        n10304), .op(n10306) );
  nand2_1 U12164 ( .ip1(n10306), .ip2(n10573), .op(
        \CORTEXM0DS_INST/u_logic/Ekhvx4 ) );
  not_ab_or_c_or_d U12165 ( .ip1(n12122), .ip2(n10308), .ip3(n10307), .ip4(
        n10565), .op(n10309) );
  not_ab_or_c_or_d U12166 ( .ip1(n10572), .ip2(n12126), .ip3(n10858), .ip4(
        n10309), .op(n10318) );
  nand2_1 U12167 ( .ip1(n10387), .ip2(n10323), .op(n10316) );
  nor2_1 U12168 ( .ip1(n10310), .ip2(n10383), .op(n10313) );
  nor2_1 U12169 ( .ip1(n10311), .ip2(n10384), .op(n10312) );
  not_ab_or_c_or_d U12170 ( .ip1(n10325), .ip2(n10389), .ip3(n10313), .ip4(
        n10312), .op(n10315) );
  nand3_1 U12171 ( .ip1(n10316), .ip2(n10315), .ip3(n10314), .op(n11256) );
  nand2_1 U12172 ( .ip1(n10859), .ip2(n11256), .op(n10317) );
  nand2_1 U12173 ( .ip1(n10318), .ip2(n10317), .op(
        \CORTEXM0DS_INST/u_logic/Lkhvx4 ) );
  inv_1 U12174 ( .ip(n10319), .op(n10321) );
  not_ab_or_c_or_d U12175 ( .ip1(n12113), .ip2(n10321), .ip3(n10320), .ip4(
        n10565), .op(n10333) );
  nand2_1 U12176 ( .ip1(n10424), .ip2(n10322), .op(n10328) );
  nand2_1 U12177 ( .ip1(n10324), .ip2(n10323), .op(n10327) );
  nand2_1 U12178 ( .ip1(n11000), .ip2(n10325), .op(n10326) );
  nand3_1 U12179 ( .ip1(n10328), .ip2(n10327), .ip3(n10326), .op(n10329) );
  not_ab_or_c_or_d U12180 ( .ip1(n11004), .ip2(n10331), .ip3(n10330), .ip4(
        n10329), .op(n11522) );
  nor2_1 U12181 ( .ip1(n11522), .ip2(n10562), .op(n10332) );
  not_ab_or_c_or_d U12182 ( .ip1(n10572), .ip2(n12117), .ip3(n10333), .ip4(
        n10332), .op(n10334) );
  nand2_1 U12183 ( .ip1(n10334), .ip2(n10573), .op(
        \CORTEXM0DS_INST/u_logic/Skhvx4 ) );
  nand2_1 U12184 ( .ip1(n12299), .ip2(n10572), .op(n10345) );
  inv_1 U12185 ( .ip(\CORTEXM0DS_INST/vis_pc [6]), .op(n12302) );
  inv_1 U12186 ( .ip(n10349), .op(n10337) );
  inv_1 U12187 ( .ip(n10335), .op(n10336) );
  not_ab_or_c_or_d U12188 ( .ip1(n12302), .ip2(n10337), .ip3(n10336), .ip4(
        n10861), .op(n10338) );
  not_ab_or_c_or_d U12189 ( .ip1(n5822), .ip2(\CORTEXM0DS_INST/vis_pc [6]), 
        .ip3(n10858), .ip4(n10338), .op(n10344) );
  inv_1 U12190 ( .ip(n10996), .op(n10849) );
  nand2_1 U12191 ( .ip1(n10849), .ip2(n10414), .op(n10342) );
  nor2_1 U12192 ( .ip1(n4130), .ip2(n10994), .op(n10340) );
  nor2_1 U12193 ( .ip1(n4150), .ip2(n10382), .op(n10339) );
  not_ab_or_c_or_d U12194 ( .ip1(n10416), .ip2(n11003), .ip3(n10340), .ip4(
        n10339), .op(n10341) );
  nand3_1 U12195 ( .ip1(n10342), .ip2(n10341), .ip3(n10371), .op(n11470) );
  nand2_1 U12196 ( .ip1(n10859), .ip2(n11470), .op(n10343) );
  nand3_1 U12197 ( .ip1(n10345), .ip2(n10344), .ip3(n10343), .op(
        \CORTEXM0DS_INST/u_logic/Zkhvx4 ) );
  nand2_1 U12198 ( .ip1(n12243), .ip2(n10572), .op(n10354) );
  nor2_1 U12199 ( .ip1(n10550), .ip2(n10382), .op(n10347) );
  nor2_1 U12200 ( .ip1(n10552), .ip2(n10994), .op(n10346) );
  ab_or_c_or_d U12201 ( .ip1(n10556), .ip2(n11003), .ip3(n10347), .ip4(n10346), 
        .op(n10348) );
  not_ab_or_c_or_d U12202 ( .ip1(n10560), .ip2(n10849), .ip3(n11002), .ip4(
        n10348), .op(n11412) );
  nor2_1 U12203 ( .ip1(n11412), .ip2(n10562), .op(n10352) );
  not_ab_or_c_or_d U12204 ( .ip1(n12244), .ip2(n10350), .ip3(n10349), .ip4(
        n10861), .op(n10351) );
  not_ab_or_c_or_d U12205 ( .ip1(n5822), .ip2(\CORTEXM0DS_INST/vis_pc [5]), 
        .ip3(n10352), .ip4(n10351), .op(n10353) );
  nand3_1 U12206 ( .ip1(n10354), .ip2(n10353), .ip3(n10573), .op(
        \CORTEXM0DS_INST/u_logic/Glhvx4 ) );
  nor2_1 U12207 ( .ip1(n10376), .ip2(n10375), .op(n10374) );
  nor2_1 U12208 ( .ip1(\CORTEXM0DS_INST/vis_pc [4]), .ip2(n10374), .op(n10355)
         );
  not_ab_or_c_or_d U12209 ( .ip1(\CORTEXM0DS_INST/vis_pc [4]), .ip2(n10374), 
        .ip3(n10355), .ip4(n10565), .op(n10364) );
  inv_1 U12210 ( .ip(n10994), .op(n10851) );
  nor2_1 U12211 ( .ip1(n10356), .ip2(n10382), .op(n10359) );
  nor2_1 U12212 ( .ip1(n10357), .ip2(n10846), .op(n10358) );
  ab_or_c_or_d U12213 ( .ip1(n10360), .ip2(n10851), .ip3(n10359), .ip4(n10358), 
        .op(n10361) );
  not_ab_or_c_or_d U12214 ( .ip1(n10362), .ip2(n10849), .ip3(n11002), .ip4(
        n10361), .op(n11403) );
  nor2_1 U12215 ( .ip1(n11403), .ip2(n10562), .op(n10363) );
  not_ab_or_c_or_d U12216 ( .ip1(n10572), .ip2(n12230), .ip3(n10364), .ip4(
        n10363), .op(n10365) );
  nand2_1 U12217 ( .ip1(n10365), .ip2(n10573), .op(
        \CORTEXM0DS_INST/u_logic/Nlhvx4 ) );
  nand2_1 U12218 ( .ip1(n10849), .ip2(n10366), .op(n10373) );
  nor2_1 U12219 ( .ip1(n4348), .ip2(n10846), .op(n10369) );
  nor2_1 U12220 ( .ip1(n10367), .ip2(n10382), .op(n10368) );
  not_ab_or_c_or_d U12221 ( .ip1(n10370), .ip2(n10851), .ip3(n10369), .ip4(
        n10368), .op(n10372) );
  nand3_1 U12222 ( .ip1(n10373), .ip2(n10372), .ip3(n10371), .op(n11395) );
  not_ab_or_c_or_d U12223 ( .ip1(n10376), .ip2(n10375), .ip3(n10374), .ip4(
        n10565), .op(n10377) );
  not_ab_or_c_or_d U12224 ( .ip1(n10859), .ip2(n11395), .ip3(n10858), .ip4(
        n10377), .op(n10379) );
  nand2_1 U12225 ( .ip1(n11397), .ip2(n10572), .op(n10378) );
  nand2_1 U12226 ( .ip1(n10379), .ip2(n10378), .op(
        \CORTEXM0DS_INST/u_logic/Ulhvx4 ) );
  nand2_1 U12227 ( .ip1(\CORTEXM0DS_INST/vis_pc [0]), .ip2(n10860), .op(n10381) );
  not_ab_or_c_or_d U12228 ( .ip1(n12394), .ip2(n10381), .ip3(n10380), .ip4(
        n10565), .op(n10391) );
  inv_1 U12229 ( .ip(n10382), .op(n10999) );
  nor2_1 U12230 ( .ip1(n10846), .ip2(n10383), .op(n10386) );
  nor2_1 U12231 ( .ip1(n10994), .ip2(n10384), .op(n10385) );
  ab_or_c_or_d U12232 ( .ip1(n10849), .ip2(n10387), .ip3(n10386), .ip4(n10385), 
        .op(n10388) );
  not_ab_or_c_or_d U12233 ( .ip1(n10999), .ip2(n10389), .ip3(n11002), .ip4(
        n10388), .op(n11254) );
  nor2_1 U12234 ( .ip1(n11254), .ip2(n10562), .op(n10390) );
  not_ab_or_c_or_d U12235 ( .ip1(n10572), .ip2(n10392), .ip3(n10391), .ip4(
        n10390), .op(n10393) );
  nand2_1 U12236 ( .ip1(n10393), .ip2(n10573), .op(
        \CORTEXM0DS_INST/u_logic/Imhvx4 ) );
  nor2_1 U12237 ( .ip1(n10395), .ip2(n10394), .op(n10404) );
  nor2_1 U12238 ( .ip1(n10397), .ip2(n10396), .op(n10403) );
  nor2_1 U12239 ( .ip1(n10398), .ip2(n10426), .op(n10402) );
  nor2_1 U12240 ( .ip1(n10400), .ip2(n10399), .op(n10401) );
  nor4_1 U12241 ( .ip1(n10404), .ip2(n10403), .ip3(n10402), .ip4(n10401), .op(
        n11352) );
  nor2_1 U12242 ( .ip1(n11352), .ip2(n10562), .op(n10411) );
  inv_1 U12243 ( .ip(\CORTEXM0DS_INST/vis_pc [18]), .op(n12188) );
  nand2_1 U12244 ( .ip1(\CORTEXM0DS_INST/vis_pc [17]), .ip2(n10405), .op(
        n10407) );
  not_ab_or_c_or_d U12245 ( .ip1(n12188), .ip2(n10407), .ip3(n10406), .ip4(
        n10565), .op(n10410) );
  nor2_1 U12246 ( .ip1(n12189), .ip2(n10855), .op(n10409) );
  or4_1 U12247 ( .ip1(n10411), .ip2(n10410), .ip3(n10409), .ip4(n10408), .op(
        \CORTEXM0DS_INST/u_logic/Ithvx4 ) );
  nor2_1 U12248 ( .ip1(n4130), .ip2(n10553), .op(n10413) );
  nor2_1 U12249 ( .ip1(n4150), .ip2(n10551), .op(n10412) );
  ab_or_c_or_d U12250 ( .ip1(n10561), .ip2(n10414), .ip3(n10413), .ip4(n10412), 
        .op(n10415) );
  not_ab_or_c_or_d U12251 ( .ip1(n10416), .ip2(n10557), .ip3(n10559), .ip4(
        n10415), .op(n11625) );
  nor2_1 U12252 ( .ip1(n11625), .ip2(n10562), .op(n10420) );
  nor2_1 U12253 ( .ip1(n10417), .ip2(n10563), .op(n10566) );
  nor2_1 U12254 ( .ip1(\CORTEXM0DS_INST/vis_pc [30]), .ip2(n10566), .op(n10418) );
  not_ab_or_c_or_d U12255 ( .ip1(\CORTEXM0DS_INST/vis_pc [30]), .ip2(n10566), 
        .ip3(n10418), .ip4(n10565), .op(n10419) );
  not_ab_or_c_or_d U12256 ( .ip1(n10572), .ip2(n10421), .ip3(n10420), .ip4(
        n10419), .op(n10422) );
  nand2_1 U12257 ( .ip1(n10422), .ip2(n10573), .op(
        \CORTEXM0DS_INST/u_logic/Wthvx4 ) );
  nand2_1 U12258 ( .ip1(n10424), .ip2(n10423), .op(n10431) );
  nor2_1 U12259 ( .ip1(n10551), .ip2(n10425), .op(n10428) );
  nor2_1 U12260 ( .ip1(n4408), .ip2(n10426), .op(n10427) );
  not_ab_or_c_or_d U12261 ( .ip1(n10557), .ip2(n11004), .ip3(n10428), .ip4(
        n10427), .op(n10430) );
  inv_1 U12262 ( .ip(n10559), .op(n10429) );
  nand3_1 U12263 ( .ip1(n10431), .ip2(n10430), .ip3(n10429), .op(n11414) );
  nor2_1 U12264 ( .ip1(n12310), .ip2(n10855), .op(n10437) );
  inv_1 U12265 ( .ip(n10432), .op(n10435) );
  inv_1 U12266 ( .ip(n10433), .op(n10434) );
  not_ab_or_c_or_d U12267 ( .ip1(n12307), .ip2(n10435), .ip3(n10434), .ip4(
        n10565), .op(n10436) );
  not_ab_or_c_or_d U12268 ( .ip1(n10859), .ip2(n11414), .ip3(n10437), .ip4(
        n10436), .op(n10438) );
  nand2_1 U12269 ( .ip1(n10438), .ip2(n10573), .op(
        \CORTEXM0DS_INST/u_logic/Duhvx4 ) );
  nand2_1 U12270 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n12642), .op(
        n11088) );
  nor3_1 U12271 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n11088), .ip3(
        n10439), .op(n10487) );
  nor2_1 U12272 ( .ip1(n12332), .ip2(n10440), .op(n10449) );
  nand3_1 U12273 ( .ip1(n10767), .ip2(n10462), .ip3(n12280), .op(n10447) );
  nor3_1 U12274 ( .ip1(n11038), .ip2(n10782), .ip3(n10441), .op(n10508) );
  nor2_1 U12275 ( .ip1(n12580), .ip2(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .op(
        n10442) );
  not_ab_or_c_or_d U12276 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(
        n10742), .ip3(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip4(n10442), .op(
        n10443) );
  nand2_1 U12277 ( .ip1(n10508), .ip2(n10443), .op(n10446) );
  nand2_1 U12278 ( .ip1(n10819), .ip2(n11746), .op(n12630) );
  nand2_1 U12279 ( .ip1(n11202), .ip2(n10444), .op(n10445) );
  nand4_1 U12280 ( .ip1(n10447), .ip2(n10446), .ip3(n12630), .ip4(n10445), 
        .op(n10448) );
  not_ab_or_c_or_d U12281 ( .ip1(n10512), .ip2(n10615), .ip3(n10449), .ip4(
        n10448), .op(n10467) );
  nand3_1 U12282 ( .ip1(n12606), .ip2(n11744), .ip3(n10908), .op(n10466) );
  nand2_1 U12283 ( .ip1(n10766), .ip2(n12580), .op(n10450) );
  nand4_1 U12284 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n10452), .ip3(
        n10451), .ip4(n10450), .op(n10453) );
  nand4_1 U12285 ( .ip1(n10455), .ip2(n10454), .ip3(n10811), .ip4(n10453), 
        .op(n10465) );
  nor3_1 U12286 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(n10782), .ip3(
        n11053), .op(n10461) );
  inv_1 U12287 ( .ip(n10456), .op(n10458) );
  nand2_1 U12288 ( .ip1(n10457), .ip2(n10517), .op(n10698) );
  nor3_1 U12289 ( .ip1(n10459), .ip2(n10458), .ip3(n10698), .op(n10460) );
  not_ab_or_c_or_d U12290 ( .ip1(n10827), .ip2(n10462), .ip3(n10461), .ip4(
        n10460), .op(n10463) );
  or2_1 U12291 ( .ip1(n10463), .ip2(n12530), .op(n10464) );
  nand4_1 U12292 ( .ip1(n10467), .ip2(n10466), .ip3(n10465), .ip4(n10464), 
        .op(n10484) );
  and3_1 U12293 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n11745), .ip3(
        n10908), .op(n10641) );
  or2_1 U12294 ( .ip1(n10790), .ip2(n10641), .op(n10469) );
  or2_1 U12295 ( .ip1(\CORTEXM0DS_INST/u_logic/Ki8vx4 ), .ip2(n10641), .op(
        n10468) );
  nand2_1 U12296 ( .ip1(n10469), .ip2(n10468), .op(n10470) );
  nor2_1 U12297 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n10470), .op(
        n10483) );
  nor3_1 U12298 ( .ip1(n10471), .ip2(n10865), .ip3(n12095), .op(n10971) );
  not_ab_or_c_or_d U12299 ( .ip1(n10473), .ip2(n12530), .ip3(n10472), .ip4(
        n10971), .op(n10481) );
  nor3_1 U12300 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip3(n10943), .op(n10478) );
  and2_1 U12301 ( .ip1(n12642), .ip2(n10719), .op(n10476) );
  nand4_1 U12302 ( .ip1(n10476), .ip2(n10500), .ip3(n10475), .ip4(n10474), 
        .op(n10477) );
  nor4_1 U12303 ( .ip1(n10970), .ip2(n10810), .ip3(n10478), .ip4(n10477), .op(
        n10480) );
  or2_1 U12304 ( .ip1(n10903), .ip2(n10479), .op(n10689) );
  nand4_1 U12305 ( .ip1(n10481), .ip2(n10480), .ip3(n11758), .ip4(n10689), 
        .op(n10482) );
  not_ab_or_c_or_d U12306 ( .ip1(n12686), .ip2(n10484), .ip3(n10483), .ip4(
        n10482), .op(n10485) );
  not_ab_or_c_or_d U12307 ( .ip1(n5938), .ip2(n11754), .ip3(1'b0), .ip4(n10485), .op(n10486) );
  or2_1 U12308 ( .ip1(n10487), .ip2(n10486), .op(
        \CORTEXM0DS_INST/u_logic/Yuhvx4 ) );
  nor2_1 U12309 ( .ip1(n12625), .ip2(n10488), .op(n10829) );
  nor2_1 U12310 ( .ip1(n11206), .ip2(n6210), .op(n10647) );
  inv_1 U12311 ( .ip(n10647), .op(n10496) );
  or2_1 U12312 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n10489), .op(
        n10593) );
  or2_1 U12313 ( .ip1(n10593), .ip2(n11231), .op(n10493) );
  nand2_1 U12314 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n10490), .op(
        n10491) );
  or2_1 U12315 ( .ip1(n10491), .ip2(n11231), .op(n10492) );
  nand2_1 U12316 ( .ip1(n10493), .ip2(n10492), .op(n10494) );
  not_ab_or_c_or_d U12317 ( .ip1(n10829), .ip2(n10496), .ip3(n10495), .ip4(
        n10494), .op(n10499) );
  nand3_1 U12318 ( .ip1(n11654), .ip2(n11077), .ip3(n10949), .op(n10497) );
  nand3_1 U12319 ( .ip1(n10499), .ip2(n10498), .ip3(n10497), .op(n10545) );
  nor3_1 U12320 ( .ip1(n10908), .ip2(n12618), .ip3(n10500), .op(n10544) );
  nand2_1 U12321 ( .ip1(n12584), .ip2(n10882), .op(n10502) );
  or2_1 U12322 ( .ip1(n10502), .ip2(n10501), .op(n10503) );
  nand2_1 U12323 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n10503), .op(
        n10748) );
  nand2_1 U12324 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/R89vx4 ), .op(n10784) );
  inv_1 U12325 ( .ip(n10784), .op(n10618) );
  nor2_1 U12326 ( .ip1(n10748), .ip2(n10618), .op(n10504) );
  not_ab_or_c_or_d U12327 ( .ip1(n10757), .ip2(n10505), .ip3(n10504), .ip4(
        n10612), .op(n10507) );
  nor4_1 U12328 ( .ip1(\CORTEXM0DS_INST/u_logic/Ho8vx4 ), .ip2(n10507), .ip3(
        n12075), .ip4(n10506), .op(n10509) );
  not_ab_or_c_or_d U12329 ( .ip1(n10511), .ip2(n10510), .ip3(n10509), .ip4(
        n10508), .op(n10521) );
  nand3_1 U12330 ( .ip1(n10512), .ip2(n12530), .ip3(n9754), .op(n10520) );
  nand3_1 U12331 ( .ip1(n10517), .ip2(n12337), .ip3(n10750), .op(n10514) );
  nand4_1 U12332 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip3(n10811), .ip4(n12580), .op(
        n10513) );
  nand3_1 U12333 ( .ip1(n10515), .ip2(n10514), .ip3(n10513), .op(n10516) );
  nand2_1 U12334 ( .ip1(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip2(n10516), .op(
        n10519) );
  nand2_1 U12335 ( .ip1(n10517), .ip2(n10782), .op(n10518) );
  nand4_1 U12336 ( .ip1(n10521), .ip2(n10520), .ip3(n10519), .ip4(n10518), 
        .op(n10525) );
  nand2_1 U12337 ( .ip1(n11754), .ip2(n12625), .op(n12335) );
  nor3_1 U12338 ( .ip1(n10676), .ip2(n12335), .ip3(n11130), .op(n10524) );
  inv_1 U12339 ( .ip(n10601), .op(n10522) );
  not_ab_or_c_or_d U12340 ( .ip1(n10865), .ip2(n10522), .ip3(
        \CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip4(n10900), .op(n10523) );
  not_ab_or_c_or_d U12341 ( .ip1(n10728), .ip2(n10525), .ip3(n10524), .ip4(
        n10523), .op(n10542) );
  nand2_1 U12342 ( .ip1(n12606), .ip2(n10726), .op(n10902) );
  inv_1 U12343 ( .ip(n10902), .op(n10529) );
  or2_1 U12344 ( .ip1(n10813), .ip2(n12588), .op(n10528) );
  nand2_1 U12345 ( .ip1(n11032), .ip2(n10526), .op(n11043) );
  or2_1 U12346 ( .ip1(n11043), .ip2(n12588), .op(n10527) );
  nand2_1 U12347 ( .ip1(n10528), .ip2(n10527), .op(n10530) );
  or2_1 U12348 ( .ip1(n10529), .ip2(n10530), .op(n10533) );
  or2_1 U12349 ( .ip1(n10531), .ip2(n10530), .op(n10532) );
  nand2_1 U12350 ( .ip1(n10533), .ip2(n10532), .op(n10534) );
  nor2_1 U12351 ( .ip1(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip2(n10534), .op(
        n10536) );
  nor3_1 U12352 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n10665), .ip3(
        n10666), .op(n10535) );
  not_ab_or_c_or_d U12353 ( .ip1(n10537), .ip2(
        \CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip3(n10536), .ip4(n10535), .op(
        n10541) );
  nand4_1 U12354 ( .ip1(n10539), .ip2(n10538), .ip3(n10959), .ip4(n10908), 
        .op(n10540) );
  nand3_1 U12355 ( .ip1(n10542), .ip2(n10541), .ip3(n10540), .op(n10543) );
  not_ab_or_c_or_d U12356 ( .ip1(n12338), .ip2(n10545), .ip3(n10544), .ip4(
        n10543), .op(n10546) );
  mux2_1 U12357 ( .ip1(n10547), .ip2(n10546), .s(n12642), .op(n10548) );
  nand2_1 U12358 ( .ip1(n10549), .ip2(n10548), .op(
        \CORTEXM0DS_INST/u_logic/Mvhvx4 ) );
  nor2_1 U12359 ( .ip1(n10551), .ip2(n10550), .op(n10555) );
  nor2_1 U12360 ( .ip1(n10553), .ip2(n10552), .op(n10554) );
  ab_or_c_or_d U12361 ( .ip1(n10557), .ip2(n10556), .ip3(n10555), .ip4(n10554), 
        .op(n10558) );
  not_ab_or_c_or_d U12362 ( .ip1(n10561), .ip2(n10560), .ip3(n10559), .ip4(
        n10558), .op(n11631) );
  nor2_1 U12363 ( .ip1(n11631), .ip2(n10562), .op(n10570) );
  inv_1 U12364 ( .ip(n10563), .op(n10564) );
  nand2_1 U12365 ( .ip1(\CORTEXM0DS_INST/vis_pc [28]), .ip2(n10564), .op(
        n10567) );
  not_ab_or_c_or_d U12366 ( .ip1(n10568), .ip2(n10567), .ip3(n10566), .ip4(
        n10565), .op(n10569) );
  not_ab_or_c_or_d U12367 ( .ip1(n10572), .ip2(n10571), .ip3(n10570), .ip4(
        n10569), .op(n10574) );
  nand2_1 U12368 ( .ip1(n10574), .ip2(n10573), .op(
        \CORTEXM0DS_INST/u_logic/Tvhvx4 ) );
  nor2_1 U12369 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Z6gvx4 ), .op(n10579) );
  nor2_1 U12370 ( .ip1(n10575), .ip2(n10816), .op(n10577) );
  not_ab_or_c_or_d U12371 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(
        n12686), .ip3(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip4(n11729), .op(
        n10576) );
  not_ab_or_c_or_d U12372 ( .ip1(n11074), .ip2(n10579), .ip3(n10577), .ip4(
        n10576), .op(n10578) );
  nor2_1 U12373 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10578), .op(
        n10585) );
  inv_1 U12374 ( .ip(n10579), .op(n10580) );
  nand2_1 U12375 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n11074), .op(
        n10815) );
  or2_1 U12376 ( .ip1(n10580), .ip2(n10815), .op(n10582) );
  nand2_1 U12377 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n10734), .op(
        n10594) );
  or2_1 U12378 ( .ip1(n10594), .ip2(n10815), .op(n10581) );
  nand2_1 U12379 ( .ip1(n10582), .ip2(n10581), .op(n10583) );
  nor4_1 U12380 ( .ip1(n10586), .ip2(n10585), .ip3(n10584), .ip4(n10583), .op(
        n10644) );
  nor2_1 U12381 ( .ip1(n12686), .ip2(n12621), .op(n10591) );
  nand3_1 U12382 ( .ip1(n11077), .ip2(n10949), .ip3(n12338), .op(n11713) );
  nor2_1 U12383 ( .ip1(n10587), .ip2(n11713), .op(n10590) );
  not_ab_or_c_or_d U12384 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(
        n10588), .ip3(n12096), .ip4(n11730), .op(n10589) );
  not_ab_or_c_or_d U12385 ( .ip1(n10591), .ip2(n11725), .ip3(n10590), .ip4(
        n10589), .op(n10643) );
  nor3_1 U12386 ( .ip1(n12614), .ip2(n10592), .ip3(n12325), .op(n10640) );
  nand2_1 U12387 ( .ip1(n12072), .ip2(n10593), .op(n10637) );
  inv_1 U12388 ( .ip(n10594), .op(n10596) );
  not_ab_or_c_or_d U12389 ( .ip1(n10820), .ip2(n10596), .ip3(
        \CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip4(n10595), .op(n10598) );
  nor3_1 U12390 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n10598), .ip3(
        n10597), .op(n10636) );
  nand2_1 U12391 ( .ip1(n12075), .ip2(n10811), .op(n10603) );
  nand2_1 U12392 ( .ip1(n5100), .ip2(n10831), .op(n10602) );
  nor3_1 U12393 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n10599), .ip3(
        n10770), .op(n10600) );
  not_ab_or_c_or_d U12394 ( .ip1(n10603), .ip2(n10602), .ip3(n10601), .ip4(
        n10600), .op(n10634) );
  nor2_1 U12395 ( .ip1(\CORTEXM0DS_INST/u_logic/R89vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/K79vx4 ), .op(n10876) );
  inv_1 U12396 ( .ip(n10876), .op(n10692) );
  inv_1 U12397 ( .ip(n12279), .op(n10604) );
  not_ab_or_c_or_d U12398 ( .ip1(n12584), .ip2(n10692), .ip3(n12580), .ip4(
        n10604), .op(n10611) );
  nor4_1 U12399 ( .ip1(\CORTEXM0DS_INST/u_logic/Sh9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip3(n9754), .ip4(n12073), .op(
        n10610) );
  not_ab_or_c_or_d U12400 ( .ip1(n10606), .ip2(n10784), .ip3(n12588), .ip4(
        n10605), .op(n10609) );
  not_ab_or_c_or_d U12401 ( .ip1(n10612), .ip2(n10607), .ip3(n11038), .ip4(
        n12592), .op(n10608) );
  nor4_1 U12402 ( .ip1(n10611), .ip2(n10610), .ip3(n10609), .ip4(n10608), .op(
        n10633) );
  nor3_1 U12403 ( .ip1(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip2(n10613), .ip3(
        n10612), .op(n10614) );
  not_ab_or_c_or_d U12404 ( .ip1(n10617), .ip2(n10616), .ip3(n10615), .ip4(
        n10614), .op(n10621) );
  nand3_1 U12405 ( .ip1(\CORTEXM0DS_INST/u_logic/K79vx4 ), .ip2(n10618), .ip3(
        n10806), .op(n10620) );
  nand2_1 U12406 ( .ip1(n10871), .ip2(n11039), .op(n10619) );
  nand4_1 U12407 ( .ip1(n10621), .ip2(n12686), .ip3(n10620), .ip4(n10619), 
        .op(n10630) );
  or2_1 U12408 ( .ip1(n11028), .ip2(n12329), .op(n10624) );
  or2_1 U12409 ( .ip1(n10622), .ip2(n12329), .op(n10623) );
  nand2_1 U12410 ( .ip1(n10624), .ip2(n10623), .op(n10629) );
  or2_1 U12411 ( .ip1(n11053), .ip2(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .op(
        n10627) );
  nand2_1 U12412 ( .ip1(n10757), .ip2(n12328), .op(n10625) );
  or2_1 U12413 ( .ip1(n10625), .ip2(\CORTEXM0DS_INST/u_logic/Aj9vx4 ), .op(
        n10626) );
  nand2_1 U12414 ( .ip1(n10627), .ip2(n10626), .op(n10628) );
  not_ab_or_c_or_d U12415 ( .ip1(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .ip2(
        n10630), .ip3(n10629), .ip4(n10628), .op(n10632) );
  nand3_1 U12416 ( .ip1(n10820), .ip2(n10776), .ip3(n11077), .op(n10631) );
  nand4_1 U12417 ( .ip1(n10634), .ip2(n10633), .ip3(n10632), .ip4(n10631), 
        .op(n10635) );
  not_ab_or_c_or_d U12418 ( .ip1(n11744), .ip2(n10637), .ip3(n10636), .ip4(
        n10635), .op(n10638) );
  nor2_1 U12419 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n10638), .op(
        n10639) );
  not_ab_or_c_or_d U12420 ( .ip1(n12082), .ip2(n10641), .ip3(n10640), .ip4(
        n10639), .op(n10642) );
  nand3_1 U12421 ( .ip1(n10644), .ip2(n10643), .ip3(n10642), .op(n10645) );
  mux2_1 U12422 ( .ip1(n10645), .ip2(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .s(
        n5938), .op(\CORTEXM0DS_INST/u_logic/Hwhvx4 ) );
  nand2_1 U12423 ( .ip1(n10776), .ip2(n11177), .op(n10660) );
  inv_1 U12424 ( .ip(n10646), .op(n10656) );
  nand2_1 U12425 ( .ip1(n11725), .ip2(n12686), .op(n12617) );
  not_ab_or_c_or_d U12426 ( .ip1(n10648), .ip2(n11700), .ip3(n10647), .ip4(
        n12617), .op(n10655) );
  nor3_1 U12427 ( .ip1(n10665), .ip2(n12651), .ip3(n10649), .op(n10651) );
  nor3_1 U12428 ( .ip1(\CORTEXM0DS_INST/u_logic/Rkgvx4 ), .ip2(n10865), .ip3(
        \CORTEXM0DS_INST/u_logic/Z6gvx4 ), .op(n10650) );
  nor2_1 U12429 ( .ip1(n10651), .ip2(n10650), .op(n10653) );
  nor2_1 U12430 ( .ip1(n10653), .ip2(n10652), .op(n10654) );
  not_ab_or_c_or_d U12431 ( .ip1(n10656), .ip2(n11771), .ip3(n10655), .ip4(
        n10654), .op(n10659) );
  nand2_1 U12432 ( .ip1(n10657), .ip2(n12338), .op(n10658) );
  nand3_1 U12433 ( .ip1(n10660), .ip2(n10659), .ip3(n10658), .op(n10740) );
  nor2_1 U12434 ( .ip1(n12616), .ip2(n12618), .op(n10662) );
  not_ab_or_c_or_d U12435 ( .ip1(n10906), .ip2(n10908), .ip3(n10662), .ip4(
        n10661), .op(n10663) );
  nor2_1 U12436 ( .ip1(n10663), .ip2(n10949), .op(n10739) );
  nand2_1 U12437 ( .ip1(n11074), .ip2(n11771), .op(n10664) );
  nand2_1 U12438 ( .ip1(n10900), .ip2(n10664), .op(n10914) );
  or2_1 U12439 ( .ip1(n12326), .ip2(n10665), .op(n10668) );
  or2_1 U12440 ( .ip1(n10666), .ip2(n10665), .op(n10667) );
  nand2_1 U12441 ( .ip1(n10668), .ip2(n10667), .op(n10675) );
  or2_1 U12442 ( .ip1(n10669), .ip2(n10950), .op(n10673) );
  nand2_1 U12443 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n10670), .op(
        n10671) );
  or2_1 U12444 ( .ip1(n10671), .ip2(n10950), .op(n10672) );
  nand2_1 U12445 ( .ip1(n10673), .ip2(n10672), .op(n10674) );
  not_ab_or_c_or_d U12446 ( .ip1(n12094), .ip2(n10914), .ip3(n10675), .ip4(
        n10674), .op(n10737) );
  inv_1 U12447 ( .ip(n10676), .op(n11201) );
  nor3_1 U12448 ( .ip1(n10679), .ip2(n10678), .ip3(n10677), .op(n10683) );
  or2_1 U12449 ( .ip1(n12621), .ip2(n12686), .op(n10681) );
  or2_1 U12450 ( .ip1(n12335), .ip2(n12686), .op(n10680) );
  nand2_1 U12451 ( .ip1(n10681), .ip2(n10680), .op(n10682) );
  not_ab_or_c_or_d U12452 ( .ip1(n11201), .ip2(n11038), .ip3(n10683), .ip4(
        n10682), .op(n10684) );
  nor3_1 U12453 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Rkgvx4 ), .ip3(n10684), .op(n10687) );
  nor2_1 U12454 ( .ip1(n10927), .ip2(n10685), .op(n10686) );
  not_ab_or_c_or_d U12455 ( .ip1(n11744), .ip2(n11698), .ip3(n10687), .ip4(
        n10686), .op(n10691) );
  nand3_1 U12456 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n10830), .ip3(
        n6210), .op(n10688) );
  nand4_1 U12457 ( .ip1(n10691), .ip2(n10690), .ip3(n10689), .ip4(n10688), 
        .op(n10725) );
  nor4_1 U12458 ( .ip1(n12554), .ip2(n12558), .ip3(n10692), .ip4(n10875), .op(
        n10695) );
  not_ab_or_c_or_d U12459 ( .ip1(\CORTEXM0DS_INST/u_logic/R89vx4 ), .ip2(
        n12588), .ip3(n10868), .ip4(n10693), .op(n10694) );
  not_ab_or_c_or_d U12460 ( .ip1(n10728), .ip2(n10696), .ip3(n10695), .ip4(
        n10694), .op(n10697) );
  nor2_1 U12461 ( .ip1(n10697), .ip2(n12592), .op(n10724) );
  nand3_1 U12462 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip3(n12580), .op(n10699) );
  not_ab_or_c_or_d U12463 ( .ip1(n10700), .ip2(n10699), .ip3(n10712), .ip4(
        n10698), .op(n10704) );
  nor2_1 U12464 ( .ip1(n10706), .ip2(n10701), .op(n10873) );
  nand2_1 U12465 ( .ip1(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip2(n12580), .op(
        n10702) );
  and3_1 U12466 ( .ip1(n10873), .ip2(\CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip3(
        n10702), .op(n10703) );
  not_ab_or_c_or_d U12467 ( .ip1(n10705), .ip2(
        \CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip3(n10704), .ip4(n10703), .op(
        n10722) );
  nor2_1 U12468 ( .ip1(n10707), .ip2(n10706), .op(n10709) );
  or2_1 U12469 ( .ip1(n10708), .ip2(n10709), .op(n10711) );
  or2_1 U12470 ( .ip1(n10726), .ip2(n10709), .op(n10710) );
  nand2_1 U12471 ( .ip1(n10711), .ip2(n10710), .op(n10721) );
  inv_1 U12472 ( .ip(n10712), .op(n10718) );
  nor2_1 U12473 ( .ip1(n11183), .ip2(n12352), .op(n10716) );
  not_ab_or_c_or_d U12474 ( .ip1(n10830), .ip2(n10713), .ip3(1'b0), .ip4(n5938), .op(n10814) );
  nand3_1 U12475 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n11170), .ip3(
        n12095), .op(n10973) );
  or2_1 U12476 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n10800), .op(
        n10714) );
  nand3_1 U12477 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10874), .ip3(
        n11730), .op(n10772) );
  nand4_1 U12478 ( .ip1(n10814), .ip2(n10973), .ip3(n10714), .ip4(n10772), 
        .op(n10715) );
  not_ab_or_c_or_d U12479 ( .ip1(n10718), .ip2(n10717), .ip3(n10716), .ip4(
        n10715), .op(n10720) );
  nand4_1 U12480 ( .ip1(n10722), .ip2(n10721), .ip3(n10720), .ip4(n10719), 
        .op(n10723) );
  not_ab_or_c_or_d U12481 ( .ip1(n12338), .ip2(n10725), .ip3(n10724), .ip4(
        n10723), .op(n10736) );
  nand3_1 U12482 ( .ip1(n10726), .ip2(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip3(
        n12647), .op(n10732) );
  nand3_1 U12483 ( .ip1(n10729), .ip2(n10728), .ip3(n10727), .op(n10730) );
  nand3_1 U12484 ( .ip1(n10732), .ip2(n10731), .ip3(n10730), .op(n10733) );
  nand2_1 U12485 ( .ip1(n10734), .ip2(n10733), .op(n10735) );
  nand3_1 U12486 ( .ip1(n10737), .ip2(n10736), .ip3(n10735), .op(n10738) );
  not_ab_or_c_or_d U12487 ( .ip1(n11650), .ip2(n10740), .ip3(n10739), .ip4(
        n10738), .op(n10741) );
  not_ab_or_c_or_d U12488 ( .ip1(n5938), .ip2(n12095), .ip3(1'b0), .ip4(n10741), .op(\CORTEXM0DS_INST/u_logic/Owhvx4 ) );
  nor2_1 U12489 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n10742), .op(
        n10744) );
  not_ab_or_c_or_d U12490 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(
        n10745), .ip3(n10744), .ip4(n10743), .op(n10747) );
  nand3_1 U12491 ( .ip1(n10748), .ip2(n10747), .ip3(n10746), .op(n10754) );
  not_ab_or_c_or_d U12492 ( .ip1(n10751), .ip2(n10750), .ip3(
        \CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip4(n10749), .op(n10752) );
  not_ab_or_c_or_d U12493 ( .ip1(n10827), .ip2(n10754), .ip3(n10753), .ip4(
        n10752), .op(n10755) );
  nor2_1 U12494 ( .ip1(\CORTEXM0DS_INST/u_logic/Ho8vx4 ), .ip2(n10755), .op(
        n10798) );
  inv_1 U12495 ( .ip(n10756), .op(n10928) );
  not_ab_or_c_or_d U12496 ( .ip1(n10758), .ip2(n10928), .ip3(n10757), .ip4(
        n12592), .op(n10765) );
  or2_1 U12497 ( .ip1(n10759), .ip2(n12530), .op(n10763) );
  nand2_1 U12498 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n10760), .op(
        n10761) );
  or2_1 U12499 ( .ip1(n10761), .ip2(n12530), .op(n10762) );
  nand2_1 U12500 ( .ip1(n10763), .ip2(n10762), .op(n10764) );
  not_ab_or_c_or_d U12501 ( .ip1(n10766), .ip2(
        \CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip3(n10765), .ip4(n10764), .op(
        n10769) );
  or2_1 U12502 ( .ip1(n11139), .ip2(n10767), .op(n10768) );
  not_ab_or_c_or_d U12503 ( .ip1(n10769), .ip2(n10768), .ip3(n12329), .ip4(
        n11038), .op(n10797) );
  nor2_1 U12504 ( .ip1(n10771), .ip2(n10770), .op(n10774) );
  nor2_1 U12505 ( .ip1(n11089), .ip2(n10772), .op(n10773) );
  nor2_1 U12506 ( .ip1(n10774), .ip2(n10773), .op(n10775) );
  nor2_1 U12507 ( .ip1(n10820), .ip2(n10775), .op(n10796) );
  nand2_1 U12508 ( .ip1(n10776), .ip2(n12082), .op(n10777) );
  nand2_1 U12509 ( .ip1(n12652), .ip2(n10777), .op(n10780) );
  not_ab_or_c_or_d U12510 ( .ip1(n11650), .ip2(n10780), .ip3(n10779), .ip4(
        n10778), .op(n10794) );
  nor3_1 U12511 ( .ip1(n11754), .ip2(n11751), .ip3(n10781), .op(n10789) );
  nor2_1 U12512 ( .ip1(n10782), .ip2(n11053), .op(n10788) );
  nor4_1 U12513 ( .ip1(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip3(n12592), .ip4(n12073), .op(
        n10787) );
  nand2_1 U12514 ( .ip1(n10784), .ip2(n10783), .op(n10785) );
  not_ab_or_c_or_d U12515 ( .ip1(n12584), .ip2(n10785), .ip3(
        \CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip4(n12073), .op(n10786) );
  nor4_1 U12516 ( .ip1(n10789), .ip2(n10788), .ip3(n10787), .ip4(n10786), .op(
        n10793) );
  nand3_1 U12517 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10790), .ip3(
        n10894), .op(n10791) );
  nand4_1 U12518 ( .ip1(n10794), .ip2(n10793), .ip3(n10792), .ip4(n10791), 
        .op(n10795) );
  nor4_1 U12519 ( .ip1(n10798), .ip2(n10797), .ip3(n10796), .ip4(n10795), .op(
        n10799) );
  nor2_1 U12520 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n10799), .op(
        n10842) );
  or2_1 U12521 ( .ip1(n10800), .ip2(n10949), .op(n10804) );
  nand3_1 U12522 ( .ip1(n10801), .ip2(n10908), .ip3(n12625), .op(n10802) );
  or2_1 U12523 ( .ip1(n10802), .ip2(n10949), .op(n10803) );
  nand2_1 U12524 ( .ip1(n10804), .ip2(n10803), .op(n10841) );
  inv_1 U12525 ( .ip(n11700), .op(n11662) );
  nor3_1 U12526 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n11662), .ip3(
        n12647), .op(n10805) );
  not_ab_or_c_or_d U12527 ( .ip1(n10806), .ip2(n11730), .ip3(
        \CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip4(n10805), .op(n10809) );
  inv_1 U12528 ( .ip(n10807), .op(n10808) );
  nor2_1 U12529 ( .ip1(n10809), .ip2(n10808), .op(n10840) );
  nor2_1 U12530 ( .ip1(n12033), .ip2(n10810), .op(n12342) );
  inv_1 U12531 ( .ip(n12330), .op(n11067) );
  nand4_1 U12532 ( .ip1(n10830), .ip2(n11067), .ip3(n11730), .ip4(n10811), 
        .op(n10812) );
  and4_1 U12533 ( .ip1(n10814), .ip2(n12342), .ip3(n10813), .ip4(n10812), .op(
        n10838) );
  not_ab_or_c_or_d U12534 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Ho8vx4 ), .ip3(n6210), .ip4(n10815), .op(
        n10818) );
  nor2_1 U12535 ( .ip1(n11212), .ip2(n10816), .op(n10817) );
  nor4_1 U12536 ( .ip1(n11198), .ip2(n10819), .ip3(n10818), .ip4(n10817), .op(
        n10837) );
  nor2_1 U12537 ( .ip1(n10820), .ip2(n10902), .op(n10826) );
  or2_1 U12538 ( .ip1(n10821), .ip2(n11211), .op(n10884) );
  nand2_1 U12539 ( .ip1(n11077), .ip2(n10822), .op(n10823) );
  or2_1 U12540 ( .ip1(n10823), .ip2(n11211), .op(n10824) );
  nand2_1 U12541 ( .ip1(n10884), .ip2(n10824), .op(n10825) );
  not_ab_or_c_or_d U12542 ( .ip1(n11726), .ip2(n11736), .ip3(n10826), .ip4(
        n10825), .op(n10836) );
  not_ab_or_c_or_d U12543 ( .ip1(\CORTEXM0DS_INST/u_logic/P39vx4 ), .ip2(
        n10829), .ip3(n10828), .ip4(n10827), .op(n10833) );
  nand3_1 U12544 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n10830), .ip3(
        n12329), .op(n10832) );
  nand4_1 U12545 ( .ip1(n10833), .ip2(n10832), .ip3(n5100), .ip4(n10831), .op(
        n10834) );
  nand2_1 U12546 ( .ip1(n11032), .ip2(n10834), .op(n10835) );
  nand4_1 U12547 ( .ip1(n10838), .ip2(n10837), .ip3(n10836), .ip4(n10835), 
        .op(n10839) );
  nor4_1 U12548 ( .ip1(n10842), .ip2(n10841), .ip3(n10840), .ip4(n10839), .op(
        n10843) );
  not_ab_or_c_or_d U12549 ( .ip1(n5938), .ip2(n6210), .ip3(1'b0), .ip4(n10843), 
        .op(\CORTEXM0DS_INST/u_logic/Vwhvx4 ) );
  nand2_1 U12550 ( .ip1(n10844), .ip2(n10999), .op(n10854) );
  nor2_1 U12551 ( .ip1(n10846), .ip2(n10845), .op(n10847) );
  not_ab_or_c_or_d U12552 ( .ip1(n10849), .ip2(n10848), .ip3(n11002), .ip4(
        n10847), .op(n10853) );
  nand2_1 U12553 ( .ip1(n10851), .ip2(n10850), .op(n10852) );
  nand3_1 U12554 ( .ip1(n10854), .ip2(n10853), .ip3(n10852), .op(n11485) );
  nor2_1 U12555 ( .ip1(n10856), .ip2(n10855), .op(n10857) );
  not_ab_or_c_or_d U12556 ( .ip1(n10859), .ip2(n11485), .ip3(n10858), .ip4(
        n10857), .op(n10863) );
  mux2_1 U12557 ( .ip1(n10861), .ip2(n10860), .s(\CORTEXM0DS_INST/vis_pc [0]), 
        .op(n10862) );
  nand2_1 U12558 ( .ip1(n10863), .ip2(n10862), .op(
        \CORTEXM0DS_INST/u_logic/Cxhvx4 ) );
  nand2_1 U12559 ( .ip1(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip2(n10864), .op(
        n5021) );
  inv_1 U12560 ( .ip(n11758), .op(n10867) );
  nor3_1 U12561 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10865), .ip3(
        n12686), .op(n10866) );
  nor2_1 U12562 ( .ip1(n10867), .ip2(n10866), .op(n5022) );
  nor4_1 U12563 ( .ip1(n10871), .ip2(n10870), .ip3(n10869), .ip4(n10868), .op(
        n10872) );
  not_ab_or_c_or_d U12564 ( .ip1(n10874), .ip2(n12078), .ip3(n10873), .ip4(
        n10872), .op(n10923) );
  or2_1 U12565 ( .ip1(\CORTEXM0DS_INST/u_logic/D69vx4 ), .ip2(n10875), .op(
        n10878) );
  or2_1 U12566 ( .ip1(n10876), .ip2(n10875), .op(n10877) );
  nand2_1 U12567 ( .ip1(n10878), .ip2(n10877), .op(n10890) );
  nor3_1 U12568 ( .ip1(n12278), .ip2(n10879), .ip3(n10950), .op(n10889) );
  nor2_1 U12569 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n10900), .op(
        n10946) );
  nand2_1 U12570 ( .ip1(n10880), .ip2(n10946), .op(n10948) );
  nand3_1 U12571 ( .ip1(n10881), .ip2(\CORTEXM0DS_INST/u_logic/Ih8vx4 ), .ip3(
        n11038), .op(n10886) );
  nand3_1 U12572 ( .ip1(n10883), .ip2(n12584), .ip3(n10882), .op(n10885) );
  nand4_1 U12573 ( .ip1(n10948), .ip2(n10886), .ip3(n10885), .ip4(n10884), 
        .op(n10887) );
  nor4_1 U12574 ( .ip1(n10890), .ip2(n10889), .ip3(n10888), .ip4(n10887), .op(
        n10922) );
  nor3_1 U12575 ( .ip1(n11105), .ip2(n11079), .ip3(n10891), .op(n12046) );
  and3_1 U12576 ( .ip1(n12096), .ip2(\CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip3(
        n12046), .op(n12050) );
  nor2_1 U12577 ( .ip1(n11183), .ip2(n10892), .op(n10893) );
  not_ab_or_c_or_d U12578 ( .ip1(n12050), .ip2(n12625), .ip3(n10893), .ip4(
        n11199), .op(n10897) );
  nand2_1 U12579 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n10894), .op(
        n10895) );
  nand2_1 U12580 ( .ip1(n6210), .ip2(n10895), .op(n10896) );
  not_ab_or_c_or_d U12581 ( .ip1(n10897), .ip2(n10896), .ip3(n10900), .ip4(
        n11730), .op(n10913) );
  nand2_1 U12582 ( .ip1(n10899), .ip2(n10898), .op(n10901) );
  not_ab_or_c_or_d U12583 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(
        n10901), .ip3(n11754), .ip4(n10900), .op(n10905) );
  nor3_1 U12584 ( .ip1(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip2(n10903), .ip3(
        n10902), .op(n10904) );
  not_ab_or_c_or_d U12585 ( .ip1(n10906), .ip2(n12625), .ip3(n10905), .ip4(
        n10904), .op(n10907) );
  or2_1 U12586 ( .ip1(n10907), .ip2(n10908), .op(n10911) );
  or2_1 U12587 ( .ip1(n10909), .ip2(n10908), .op(n10910) );
  nand2_1 U12588 ( .ip1(n10911), .ip2(n10910), .op(n10912) );
  not_ab_or_c_or_d U12589 ( .ip1(n10915), .ip2(n10914), .ip3(n10913), .ip4(
        n10912), .op(n10921) );
  nand4_1 U12590 ( .ip1(n10919), .ip2(n10918), .ip3(n10917), .ip4(n10916), 
        .op(n10920) );
  nand4_1 U12591 ( .ip1(n10923), .ip2(n10922), .ip3(n10921), .ip4(n10920), 
        .op(n10924) );
  mux2_1 U12592 ( .ip1(n10924), .ip2(\CORTEXM0DS_INST/u_logic/Cn8vx4 ), .s(
        n5938), .op(\CORTEXM0DS_INST/u_logic/Xxhvx4 ) );
  nor2_1 U12593 ( .ip1(n12588), .ip2(n10925), .op(n10929) );
  nor4_1 U12594 ( .ip1(n10929), .ip2(n10928), .ip3(n10927), .ip4(n10926), .op(
        n10931) );
  not_ab_or_c_or_d U12595 ( .ip1(n10933), .ip2(n10932), .ip3(n10931), .ip4(
        n10930), .op(n10962) );
  nand3_1 U12596 ( .ip1(n11130), .ip2(n10934), .ip3(n12325), .op(n10958) );
  not_ab_or_c_or_d U12597 ( .ip1(n10936), .ip2(n10935), .ip3(n12618), .ip4(
        n12352), .op(n10957) );
  nand2_1 U12598 ( .ip1(n10937), .ip2(n11074), .op(n11131) );
  or2_1 U12599 ( .ip1(n11131), .ip2(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .op(
        n10942) );
  nand2_1 U12600 ( .ip1(n10939), .ip2(n10938), .op(n10940) );
  or2_1 U12601 ( .ip1(n10940), .ip2(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .op(
        n10941) );
  nand2_1 U12602 ( .ip1(n10942), .ip2(n10941), .op(n10955) );
  inv_1 U12603 ( .ip(n11169), .op(n10944) );
  nor3_1 U12604 ( .ip1(\CORTEXM0DS_INST/u_logic/Q5gvx4 ), .ip2(n10944), .ip3(
        n10943), .op(n10945) );
  nor2_1 U12605 ( .ip1(n10946), .ip2(n10945), .op(n10947) );
  nor2_1 U12606 ( .ip1(n10947), .ip2(n11212), .op(n10954) );
  nor2_1 U12607 ( .ip1(n10949), .ip2(n10948), .op(n10953) );
  nor2_1 U12608 ( .ip1(n10951), .ip2(n10950), .op(n10952) );
  or4_1 U12609 ( .ip1(n10955), .ip2(n10954), .ip3(n10953), .ip4(n10952), .op(
        n10956) );
  not_ab_or_c_or_d U12610 ( .ip1(n6210), .ip2(n10958), .ip3(n10957), .ip4(
        n10956), .op(n10961) );
  nand3_1 U12611 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n11195), .ip3(
        n10959), .op(n10960) );
  nand3_1 U12612 ( .ip1(n10962), .ip2(n10961), .ip3(n10960), .op(n10963) );
  mux2_1 U12613 ( .ip1(n10963), .ip2(\CORTEXM0DS_INST/u_logic/Dw8vx4 ), .s(
        n5938), .op(\CORTEXM0DS_INST/u_logic/Lyhvx4 ) );
  nor2_1 U12614 ( .ip1(n10964), .ip2(n12295), .op(n10968) );
  not_ab_or_c_or_d U12615 ( .ip1(n10966), .ip2(n10965), .ip3(n12155), .ip4(
        n12305), .op(n10967) );
  not_ab_or_c_or_d U12616 ( .ip1(n12300), .ip2(n11535), .ip3(n10968), .ip4(
        n10967), .op(\CORTEXM0DS_INST/u_logic/N1447 ) );
  nand3_1 U12617 ( .ip1(n11199), .ip2(n10969), .ip3(n12625), .op(n12351) );
  nor2_1 U12618 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n12351), .op(
        n11720) );
  not_ab_or_c_or_d U12619 ( .ip1(n10972), .ip2(n10971), .ip3(n10970), .ip4(
        n11720), .op(n10974) );
  nand3_1 U12620 ( .ip1(n10974), .ip2(n10973), .ip3(n11222), .op(n3217) );
  nand2_1 U12621 ( .ip1(\CORTEXM0DS_INST/vis_ipsr [3]), .ip2(n4831), .op(
        n10979) );
  nand2_1 U12622 ( .ip1(n3217), .ip2(n10975), .op(n11778) );
  nor2_1 U12623 ( .ip1(n5938), .ip2(n11778), .op(n11025) );
  nand2_1 U12624 ( .ip1(n11025), .ip2(n11388), .op(n10978) );
  inv_1 U12625 ( .ip(n4831), .op(n12393) );
  inv_1 U12626 ( .ip(n12078), .op(n11190) );
  nand2_1 U12627 ( .ip1(n10976), .ip2(n11190), .op(n12027) );
  nand2_1 U12628 ( .ip1(n12393), .ip2(n12027), .op(n12025) );
  nor2_1 U12629 ( .ip1(n12446), .ip2(n12025), .op(n10983) );
  nand2_1 U12630 ( .ip1(\CORTEXM0DS_INST/u_logic/Lrevx4 ), .ip2(n10983), .op(
        n10977) );
  nand3_1 U12631 ( .ip1(n10979), .ip2(n10978), .ip3(n10977), .op(
        \CORTEXM0DS_INST/u_logic/L8mvx4 ) );
  inv_1 U12632 ( .ip(n11025), .op(n11005) );
  nor2_1 U12633 ( .ip1(n11254), .ip2(n11005), .op(n10982) );
  nor2_1 U12634 ( .ip1(n10980), .ip2(n12393), .op(n10981) );
  ab_or_c_or_d U12635 ( .ip1(n10983), .ip2(\CORTEXM0DS_INST/u_logic/Bqevx4 ), 
        .ip3(n10982), .ip4(n10981), .op(\CORTEXM0DS_INST/u_logic/U9mvx4 ) );
  nand2_1 U12636 ( .ip1(n4831), .ip2(\CORTEXM0DS_INST/vis_ipsr [4]), .op(
        n10986) );
  nand2_1 U12637 ( .ip1(n11025), .ip2(n11395), .op(n10985) );
  nand2_1 U12638 ( .ip1(\CORTEXM0DS_INST/u_logic/Vsevx4 ), .ip2(n10983), .op(
        n10984) );
  nand3_1 U12639 ( .ip1(n10986), .ip2(n10985), .ip3(n10984), .op(
        \CORTEXM0DS_INST/u_logic/Pamvx4 ) );
  nor2_1 U12640 ( .ip1(n11403), .ip2(n11005), .op(n10988) );
  inv_1 U12641 ( .ip(\CORTEXM0DS_INST/u_logic/Fuevx4 ), .op(n12559) );
  nor3_1 U12642 ( .ip1(n12446), .ip2(n12559), .ip3(n12025), .op(n10987) );
  ab_or_c_or_d U12643 ( .ip1(n4831), .ip2(\CORTEXM0DS_INST/vis_ipsr [5]), 
        .ip3(n10988), .ip4(n10987), .op(\CORTEXM0DS_INST/u_logic/Wamvx4 ) );
  nand2_1 U12644 ( .ip1(\CORTEXM0DS_INST/u_logic/G8fvx4 ), .ip2(n10989), .op(
        n10990) );
  nand3_1 U12645 ( .ip1(n10990), .ip2(n4816), .ip3(n12024), .op(
        \CORTEXM0DS_INST/u_logic/G8nvx4 ) );
  inv_1 U12646 ( .ip(\CORTEXM0DS_INST/u_logic/Roevx4 ), .op(n12539) );
  nor3_1 U12647 ( .ip1(n12446), .ip2(n12539), .ip3(n12025), .op(n10993) );
  nor2_1 U12648 ( .ip1(n10991), .ip2(n12393), .op(n10992) );
  ab_or_c_or_d U12649 ( .ip1(n11025), .ip2(n11485), .ip3(n10993), .ip4(n10992), 
        .op(\CORTEXM0DS_INST/u_logic/Acnvx4 ) );
  nor2_1 U12650 ( .ip1(n10995), .ip2(n10994), .op(n10998) );
  nor2_1 U12651 ( .ip1(n4408), .ip2(n10996), .op(n10997) );
  ab_or_c_or_d U12652 ( .ip1(n11000), .ip2(n10999), .ip3(n10998), .ip4(n10997), 
        .op(n11001) );
  not_ab_or_c_or_d U12653 ( .ip1(n11004), .ip2(n11003), .ip3(n11002), .ip4(
        n11001), .op(n11473) );
  nor2_1 U12654 ( .ip1(n11473), .ip2(n11005), .op(n11007) );
  nand2_1 U12655 ( .ip1(\CORTEXM0DS_INST/u_logic/Hnevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Xlevx4 ), .op(n12454) );
  nor2_1 U12656 ( .ip1(n12454), .ip2(n12025), .op(n11006) );
  ab_or_c_or_d U12657 ( .ip1(n4831), .ip2(\CORTEXM0DS_INST/vis_ipsr [0]), 
        .ip3(n11007), .ip4(n11006), .op(\CORTEXM0DS_INST/u_logic/Ocnvx4 ) );
  nand2_1 U12658 ( .ip1(n11768), .ip2(n11008), .op(n11776) );
  nand2_1 U12659 ( .ip1(n11776), .ip2(n11778), .op(n11633) );
  inv_1 U12660 ( .ip(n11633), .op(n11783) );
  nor2_1 U12661 ( .ip1(n11009), .ip2(n11776), .op(n11011) );
  nor2_1 U12662 ( .ip1(n11467), .ip2(n11778), .op(n11010) );
  ab_or_c_or_d U12663 ( .ip1(n11783), .ip2(n11012), .ip3(n11011), .ip4(n11010), 
        .op(n11015) );
  not_ab_or_c_or_d U12664 ( .ip1(n11013), .ip2(n11783), .ip3(1'b0), .ip4(n5938), .op(n11014) );
  mux2_1 U12665 ( .ip1(\CORTEXM0DS_INST/vis_apsr [0]), .ip2(n11015), .s(n11014), .op(\CORTEXM0DS_INST/u_logic/Rhnvx4 ) );
  nor2_1 U12666 ( .ip1(n11016), .ip2(n11473), .op(n11020) );
  nor2_1 U12667 ( .ip1(n11018), .ip2(n11017), .op(n11019) );
  ab_or_c_or_d U12668 ( .ip1(n11025), .ip2(n11414), .ip3(n11020), .ip4(n11019), 
        .op(n11027) );
  nor2_1 U12669 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Mcgvx4 ), .op(n11021) );
  not_ab_or_c_or_d U12670 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(
        n11022), .ip3(n11202), .ip4(n11021), .op(n11023) );
  nor3_1 U12671 ( .ip1(n11023), .ip2(LOCKUP_top_out), .ip3(n12091), .op(n11024) );
  nor2_1 U12672 ( .ip1(n11025), .ip2(n11024), .op(n11026) );
  mux2_1 U12673 ( .ip1(n11027), .ip2(\CORTEXM0DS_INST/cm0_xpsr[24] ), .s(
        n11026), .op(\CORTEXM0DS_INST/u_logic/Ojnvx4 ) );
  nor2_1 U12674 ( .ip1(n11790), .ip2(n12635), .op(n4712) );
  inv_1 U12675 ( .ip(n3227), .op(n12638) );
  mux2_1 U12676 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [31]), .ip2(n12638), 
        .s(n4712), .op(\CORTEXM0DS_INST/u_logic/Vkmvx4 ) );
  inv_1 U12677 ( .ip(n3226), .op(n4711) );
  mux2_1 U12678 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [29]), .ip2(n4711), .s(
        n4712), .op(\CORTEXM0DS_INST/u_logic/Jlmvx4 ) );
  nand2_1 U12679 ( .ip1(n11827), .ip2(\CORTEXM0DS_INST/u_logic/Mf8vx4 ), .op(
        n4708) );
  mux2_1 U12680 ( .ip1(n12638), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [23]), 
        .s(n4708), .op(\CORTEXM0DS_INST/u_logic/Rimvx4 ) );
  mux2_1 U12681 ( .ip1(n4711), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [21]), .s(
        n4708), .op(\CORTEXM0DS_INST/u_logic/Fjmvx4 ) );
  and2_1 U12682 ( .ip1(n11833), .ip2(\CORTEXM0DS_INST/u_logic/Mf8vx4 ), .op(
        n4706) );
  mux2_1 U12683 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [15]), .ip2(n12638), 
        .s(n4706), .op(\CORTEXM0DS_INST/u_logic/Ngmvx4 ) );
  mux2_1 U12684 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [13]), .ip2(n4711), .s(
        n4706), .op(\CORTEXM0DS_INST/u_logic/Bhmvx4 ) );
  nand2_1 U12685 ( .ip1(n11824), .ip2(\CORTEXM0DS_INST/u_logic/Mf8vx4 ), .op(
        n4704) );
  mux2_1 U12686 ( .ip1(n12638), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [7]), .s(
        n4704), .op(\CORTEXM0DS_INST/u_logic/Jemvx4 ) );
  mux2_1 U12687 ( .ip1(n4711), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [5]), .s(
        n4704), .op(\CORTEXM0DS_INST/u_logic/Xemvx4 ) );
  or2_1 U12688 ( .ip1(n11028), .ip2(n12330), .op(n11031) );
  or2_1 U12689 ( .ip1(n11029), .ip2(n12330), .op(n11030) );
  nand2_1 U12690 ( .ip1(n11031), .ip2(n11030), .op(n11111) );
  nand3_1 U12691 ( .ip1(n11033), .ip2(n12328), .ip3(n11032), .op(n11109) );
  nor2_1 U12692 ( .ip1(n9754), .ip2(n11109), .op(n11037) );
  inv_1 U12693 ( .ip(\CORTEXM0DS_INST/u_logic/Lrevx4 ), .op(n12549) );
  nand2_1 U12694 ( .ip1(n11184), .ip2(n11164), .op(n11034) );
  nand2_1 U12695 ( .ip1(n11035), .ip2(n11034), .op(n11121) );
  nand2_1 U12696 ( .ip1(\CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip2(n11121), .op(
        n11146) );
  nor2_1 U12697 ( .ip1(n12549), .ip2(n11146), .op(n11036) );
  not_ab_or_c_or_d U12698 ( .ip1(\CORTEXM0DS_INST/u_logic/I29vx4 ), .ip2(
        n11111), .ip3(n11037), .ip4(n11036), .op(n11087) );
  nand3_1 U12699 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n11725), .ip3(
        n11038), .op(n11042) );
  nand4_1 U12700 ( .ip1(n11040), .ip2(n11039), .ip3(n12530), .ip4(n12338), 
        .op(n11041) );
  and4_1 U12701 ( .ip1(n11044), .ip2(n11043), .ip3(n11042), .ip4(n11041), .op(
        n11140) );
  nor2_1 U12702 ( .ip1(n11140), .ip2(n12550), .op(n11083) );
  inv_1 U12703 ( .ip(n11045), .op(n11048) );
  mux2_1 U12704 ( .ip1(n11048), .ip2(n11045), .s(n11047), .op(n11059) );
  nand2_1 U12705 ( .ip1(\CORTEXM0DS_INST/u_logic/R89vx4 ), .ip2(n11059), .op(
        n11114) );
  fulladder U12706 ( .a(\CORTEXM0DS_INST/u_logic/B19vx4 ), .b(
        \CORTEXM0DS_INST/u_logic/I29vx4 ), .ci(
        \CORTEXM0DS_INST/u_logic/Uz8vx4 ), .co(n11062), .s(n11046) );
  fulladder U12707 ( .a(\CORTEXM0DS_INST/u_logic/W49vx4 ), .b(
        \CORTEXM0DS_INST/u_logic/P39vx4 ), .ci(n11046), .co(n11061), .s(n11047) );
  nand2_1 U12708 ( .ip1(\CORTEXM0DS_INST/u_logic/K79vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/D69vx4 ), .op(n11050) );
  nand2_1 U12709 ( .ip1(n11048), .ip2(n11047), .op(n11049) );
  nand2_1 U12710 ( .ip1(n11050), .ip2(n11049), .op(n11060) );
  inv_1 U12711 ( .ip(n11051), .op(n11113) );
  nor2_1 U12712 ( .ip1(n11114), .ip2(n11113), .op(n11117) );
  nand3_1 U12713 ( .ip1(n11117), .ip2(n11061), .ip3(n11062), .op(n11058) );
  or2_1 U12714 ( .ip1(n11052), .ip2(n11054), .op(n11057) );
  inv_1 U12715 ( .ip(n11053), .op(n11055) );
  or2_1 U12716 ( .ip1(n11055), .ip2(n11054), .op(n11056) );
  nand2_1 U12717 ( .ip1(n11057), .ip2(n11056), .op(n11136) );
  or2_1 U12718 ( .ip1(n11058), .ip2(n11136), .op(n11066) );
  mux2_1 U12719 ( .ip1(n12570), .ip2(\CORTEXM0DS_INST/u_logic/R89vx4 ), .s(
        n11059), .op(n11138) );
  nor2_1 U12720 ( .ip1(n11139), .ip2(n11138), .op(n11137) );
  inv_1 U12721 ( .ip(n11137), .op(n11112) );
  nor2_1 U12722 ( .ip1(n11113), .ip2(n11112), .op(n11116) );
  fulladder U12723 ( .a(n11062), .b(n11061), .ci(n11060), .co(n11064), .s(
        n11051) );
  nand2_1 U12724 ( .ip1(n11062), .ip2(n11061), .op(n11063) );
  mux2_1 U12725 ( .ip1(n11064), .ip2(n11063), .s(n11117), .op(n11096) );
  nand2_1 U12726 ( .ip1(n11116), .ip2(n11096), .op(n11099) );
  or2_1 U12727 ( .ip1(n11099), .ip2(n11136), .op(n11065) );
  nand2_1 U12728 ( .ip1(n11066), .ip2(n11065), .op(n11082) );
  nand2_1 U12729 ( .ip1(n11068), .ip2(n11067), .op(n12054) );
  and2_1 U12730 ( .ip1(n11069), .ip2(n12054), .op(n11072) );
  nand2_1 U12731 ( .ip1(n11072), .ip2(n11070), .op(n11071) );
  nand2_1 U12732 ( .ip1(n12329), .ip2(n11071), .op(n11093) );
  not_ab_or_c_or_d U12733 ( .ip1(n11072), .ip2(
        \CORTEXM0DS_INST/u_logic/Ud9vx4 ), .ip3(n12580), .ip4(n11093), .op(
        n11081) );
  nand2_1 U12734 ( .ip1(n11073), .ip2(\CORTEXM0DS_INST/u_logic/Qm9vx4 ), .op(
        n11078) );
  and2_1 U12735 ( .ip1(n11661), .ip2(n11074), .op(n11076) );
  not_ab_or_c_or_d U12736 ( .ip1(n11660), .ip2(n11077), .ip3(n11076), .ip4(
        n11075), .op(n12049) );
  not_ab_or_c_or_d U12737 ( .ip1(n11079), .ip2(n11078), .ip3(n12049), .ip4(
        n12046), .op(n11080) );
  nor4_1 U12738 ( .ip1(n11083), .ip2(n11082), .ip3(n11081), .ip4(n11080), .op(
        n11086) );
  nand4_1 U12739 ( .ip1(n11087), .ip2(n11086), .ip3(n11085), .ip4(n11084), 
        .op(n11091) );
  inv_1 U12740 ( .ip(n11088), .op(n12645) );
  nand3_1 U12741 ( .ip1(n11089), .ip2(n12645), .ip3(n11161), .op(n11090) );
  nand2_1 U12742 ( .ip1(n4627), .ip2(n11090), .op(n11151) );
  mux2_1 U12743 ( .ip1(\CORTEXM0DS_INST/u_logic/Un9vx4 ), .ip2(n11091), .s(
        n11151), .op(\CORTEXM0DS_INST/u_logic/N2mvx4 ) );
  inv_1 U12744 ( .ip(n11109), .op(n12058) );
  not_ab_or_c_or_d U12745 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(
        n12544), .ip3(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip4(n11729), .op(
        n11134) );
  inv_1 U12746 ( .ip(\CORTEXM0DS_INST/u_logic/Bqevx4 ), .op(n12545) );
  nor2_1 U12747 ( .ip1(n12545), .ip2(n11146), .op(n11092) );
  not_ab_or_c_or_d U12748 ( .ip1(n12058), .ip2(
        \CORTEXM0DS_INST/u_logic/R89vx4 ), .ip3(n11134), .ip4(n11092), .op(
        n11103) );
  inv_1 U12749 ( .ip(n11093), .op(n11143) );
  nor3_1 U12750 ( .ip1(\CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip2(n12049), .ip3(
        n11105), .op(n11095) );
  nor2_1 U12751 ( .ip1(n11140), .ip2(n12544), .op(n11094) );
  not_ab_or_c_or_d U12752 ( .ip1(n11143), .ip2(
        \CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip3(n11095), .ip4(n11094), .op(
        n11102) );
  or2_1 U12753 ( .ip1(n11116), .ip2(n11096), .op(n11098) );
  inv_1 U12754 ( .ip(n11136), .op(n11097) );
  nand3_1 U12755 ( .ip1(n11099), .ip2(n11098), .ip3(n11097), .op(n11101) );
  nand2_1 U12756 ( .ip1(\CORTEXM0DS_INST/u_logic/B19vx4 ), .ip2(n11111), .op(
        n11100) );
  nand4_1 U12757 ( .ip1(n11103), .ip2(n11102), .ip3(n11101), .ip4(n11100), 
        .op(n11104) );
  nand2_1 U12758 ( .ip1(n11104), .ip2(n11151), .op(n11108) );
  inv_1 U12759 ( .ip(n12049), .op(n11144) );
  nand2_1 U12760 ( .ip1(n11105), .ip2(n11144), .op(n11106) );
  nand2_1 U12761 ( .ip1(n11151), .ip2(n11106), .op(n11127) );
  nand2_1 U12762 ( .ip1(\CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip2(n11127), .op(
        n11107) );
  nand2_1 U12763 ( .ip1(n11108), .ip2(n11107), .op(
        \CORTEXM0DS_INST/u_logic/U2mvx4 ) );
  nor2_1 U12764 ( .ip1(n12564), .ip2(n11109), .op(n11110) );
  not_ab_or_c_or_d U12765 ( .ip1(n11111), .ip2(
        \CORTEXM0DS_INST/u_logic/Uz8vx4 ), .ip3(n11134), .ip4(n11110), .op(
        n11125) );
  and3_1 U12766 ( .ip1(n11114), .ip2(n11113), .ip3(n11112), .op(n11115) );
  nor4_1 U12767 ( .ip1(n11136), .ip2(n11117), .ip3(n11116), .ip4(n11115), .op(
        n11119) );
  inv_1 U12768 ( .ip(\CORTEXM0DS_INST/u_logic/B19vx4 ), .op(n12540) );
  nor2_1 U12769 ( .ip1(n11140), .ip2(n12540), .op(n11118) );
  not_ab_or_c_or_d U12770 ( .ip1(n11143), .ip2(
        \CORTEXM0DS_INST/u_logic/R89vx4 ), .ip3(n11119), .ip4(n11118), .op(
        n11124) );
  nand2_1 U12771 ( .ip1(n11120), .ip2(n11144), .op(n11123) );
  nand3_1 U12772 ( .ip1(\CORTEXM0DS_INST/u_logic/Roevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip3(n11121), .op(n11122) );
  nand4_1 U12773 ( .ip1(n11125), .ip2(n11124), .ip3(n11123), .ip4(n11122), 
        .op(n11126) );
  nand2_1 U12774 ( .ip1(n11126), .ip2(n11151), .op(n11129) );
  nand2_1 U12775 ( .ip1(\CORTEXM0DS_INST/u_logic/Ml9vx4 ), .ip2(n11127), .op(
        n11128) );
  nand2_1 U12776 ( .ip1(n11129), .ip2(n11128), .op(
        \CORTEXM0DS_INST/u_logic/Jdnvx4 ) );
  nand4_1 U12777 ( .ip1(n11132), .ip2(n11131), .ip3(n11130), .ip4(n12325), 
        .op(n11133) );
  not_ab_or_c_or_d U12778 ( .ip1(n11135), .ip2(n12588), .ip3(n11134), .ip4(
        n11133), .op(n11150) );
  not_ab_or_c_or_d U12779 ( .ip1(n11139), .ip2(n11138), .ip3(n11137), .ip4(
        n11136), .op(n11142) );
  nor2_1 U12780 ( .ip1(n11140), .ip2(n12535), .op(n11141) );
  not_ab_or_c_or_d U12781 ( .ip1(n11143), .ip2(
        \CORTEXM0DS_INST/u_logic/K79vx4 ), .ip3(n11142), .ip4(n11141), .op(
        n11149) );
  nand2_1 U12782 ( .ip1(n11145), .ip2(n11144), .op(n11148) );
  inv_1 U12783 ( .ip(\CORTEXM0DS_INST/u_logic/Hnevx4 ), .op(n12534) );
  or2_1 U12784 ( .ip1(n12534), .ip2(n11146), .op(n11147) );
  nand4_1 U12785 ( .ip1(n11150), .ip2(n11149), .ip3(n11148), .ip4(n11147), 
        .op(n11152) );
  mux2_1 U12786 ( .ip1(\CORTEXM0DS_INST/u_logic/Ik9vx4 ), .ip2(n11152), .s(
        n11151), .op(\CORTEXM0DS_INST/u_logic/Tinvx4 ) );
  mux2_1 U12787 ( .ip1(n11153), .ip2(\CORTEXM0DS_INST/u_logic/Zph2z4 [1]), .s(
        n4585), .op(\CORTEXM0DS_INST/u_logic/X9kvx4 ) );
  mux2_1 U12788 ( .ip1(n12286), .ip2(\CORTEXM0DS_INST/u_logic/Zph2z4 [0]), .s(
        n4585), .op(\CORTEXM0DS_INST/u_logic/Ufnvx4 ) );
  nand2_1 U12789 ( .ip1(n11549), .ip2(n12659), .op(n11157) );
  nor3_1 U12790 ( .ip1(n11155), .ip2(n11154), .ip3(n11719), .op(n11156) );
  nand3_1 U12791 ( .ip1(n11157), .ip2(n11156), .ip3(n11451), .op(n11577) );
  nor2_1 U12792 ( .ip1(n11237), .ip2(n11158), .op(n11234) );
  nor2_1 U12793 ( .ip1(n11238), .ip2(n11159), .op(n11233) );
  nor2_1 U12794 ( .ip1(n11239), .ip2(n11160), .op(n11232) );
  nand2_1 U12795 ( .ip1(n11161), .ip2(\CORTEXM0DS_INST/u_logic/Whgvx4 ), .op(
        n11167) );
  nand2_1 U12796 ( .ip1(n11162), .ip2(n12335), .op(n11163) );
  nand2_1 U12797 ( .ip1(n11164), .ip2(n11163), .op(n11165) );
  nand3_1 U12798 ( .ip1(n11167), .ip2(n11166), .ip3(n11165), .op(n11228) );
  nor2_1 U12799 ( .ip1(n6210), .ip2(n11168), .op(n11176) );
  or2_1 U12800 ( .ip1(n11169), .ip2(n11170), .op(n11172) );
  or2_1 U12801 ( .ip1(n12686), .ip2(n11170), .op(n11171) );
  nand2_1 U12802 ( .ip1(n11172), .ip2(n11171), .op(n11173) );
  nor2_1 U12803 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n11173), .op(
        n11174) );
  not_ab_or_c_or_d U12804 ( .ip1(n11177), .ip2(n11176), .ip3(n11175), .ip4(
        n11174), .op(n11178) );
  nor2_1 U12805 ( .ip1(n11178), .ip2(n12618), .op(n11227) );
  nor2_1 U12806 ( .ip1(n12072), .ip2(n11750), .op(n11179) );
  not_ab_or_c_or_d U12807 ( .ip1(n11182), .ip2(n11181), .ip3(n11180), .ip4(
        n11179), .op(n11225) );
  inv_1 U12808 ( .ip(n11183), .op(n11194) );
  and2_1 U12809 ( .ip1(n11184), .ip2(n11660), .op(n11185) );
  or2_1 U12810 ( .ip1(n12082), .ip2(n11185), .op(n11188) );
  or2_1 U12811 ( .ip1(n11186), .ip2(n11185), .op(n11187) );
  nand2_1 U12812 ( .ip1(n11188), .ip2(n11187), .op(n11189) );
  nor2_1 U12813 ( .ip1(n11189), .ip2(n12625), .op(n11193) );
  nor3_1 U12814 ( .ip1(\CORTEXM0DS_INST/u_logic/Nggvx4 ), .ip2(n11191), .ip3(
        n11190), .op(n11192) );
  ab_or_c_or_d U12815 ( .ip1(n11195), .ip2(n11194), .ip3(n11193), .ip4(n11192), 
        .op(n11196) );
  not_ab_or_c_or_d U12816 ( .ip1(n11199), .ip2(n11198), .ip3(n11197), .ip4(
        n11196), .op(n11224) );
  nand3_1 U12817 ( .ip1(n11654), .ip2(n11200), .ip3(n11698), .op(n11204) );
  nand2_1 U12818 ( .ip1(n11202), .ip2(n11201), .op(n11203) );
  nand2_1 U12819 ( .ip1(n11204), .ip2(n11203), .op(n11221) );
  or3_1 U12820 ( .ip1(n12095), .ip2(n12653), .ip3(n12613), .op(n11205) );
  or2_1 U12821 ( .ip1(n11205), .ip2(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .op(
        n11210) );
  nand3_1 U12822 ( .ip1(n11207), .ip2(n11206), .ip3(n11736), .op(n11208) );
  or2_1 U12823 ( .ip1(n11208), .ip2(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .op(
        n11209) );
  nand2_1 U12824 ( .ip1(n11210), .ip2(n11209), .op(n11220) );
  nor3_1 U12825 ( .ip1(n12625), .ip2(n11212), .ip3(n11211), .op(n11216) );
  nor2_1 U12826 ( .ip1(n11214), .ip2(n11213), .op(n11215) );
  not_ab_or_c_or_d U12827 ( .ip1(n11217), .ip2(n10865), .ip3(n11216), .ip4(
        n11215), .op(n11218) );
  nor2_1 U12828 ( .ip1(n11218), .ip2(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .op(
        n11219) );
  not_ab_or_c_or_d U12829 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(
        n11221), .ip3(n11220), .ip4(n11219), .op(n11223) );
  nand4_1 U12830 ( .ip1(n11225), .ip2(n11224), .ip3(n11223), .ip4(n11222), 
        .op(n11226) );
  not_ab_or_c_or_d U12831 ( .ip1(n11229), .ip2(n11228), .ip3(n11227), .ip4(
        n11226), .op(n11230) );
  nor2_1 U12832 ( .ip1(n5938), .ip2(n11230), .op(n11235) );
  nand2_1 U12833 ( .ip1(n11235), .ip2(n11231), .op(n11250) );
  nor4_1 U12834 ( .ip1(n11234), .ip2(n11233), .ip3(n11232), .ip4(n11250), .op(
        n11496) );
  nand2_1 U12835 ( .ip1(n11235), .ip2(n11556), .op(n11490) );
  nor2_1 U12836 ( .ip1(n11496), .ip2(n11490), .op(n11494) );
  inv_1 U12837 ( .ip(n11236), .op(n11249) );
  inv_1 U12838 ( .ip(n11237), .op(n11244) );
  nand2_1 U12839 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [2]), .ip2(n11244), 
        .op(n11242) );
  inv_1 U12840 ( .ip(n11238), .op(n11243) );
  nand2_1 U12841 ( .ip1(\CORTEXM0DS_INST/u_logic/Wv9vx4 ), .ip2(n11243), .op(
        n11241) );
  inv_1 U12842 ( .ip(n11239), .op(n11245) );
  nand2_1 U12843 ( .ip1(\CORTEXM0DS_INST/u_logic/Nt8vx4 ), .ip2(n11245), .op(
        n11240) );
  nand4_1 U12844 ( .ip1(n11249), .ip2(n11242), .ip3(n11241), .ip4(n11240), 
        .op(n11491) );
  nor2_1 U12845 ( .ip1(n11250), .ip2(n11491), .op(n11503) );
  nand2_1 U12846 ( .ip1(\CORTEXM0DS_INST/u_logic/Bx9vx4 ), .ip2(n11243), .op(
        n11248) );
  nand2_1 U12847 ( .ip1(\CORTEXM0DS_INST/u_logic/Tjh2z4 [3]), .ip2(n11244), 
        .op(n11247) );
  nand2_1 U12848 ( .ip1(\CORTEXM0DS_INST/u_logic/Vu8vx4 ), .ip2(n11245), .op(
        n11246) );
  nand4_1 U12849 ( .ip1(n11249), .ip2(n11248), .ip3(n11247), .ip4(n11246), 
        .op(n11501) );
  nor2_1 U12850 ( .ip1(n11250), .ip2(n11501), .op(n11492) );
  nor2_1 U12851 ( .ip1(n11503), .ip2(n11492), .op(n11557) );
  nand2_1 U12852 ( .ip1(n11494), .ip2(n11557), .op(n11525) );
  nor2_1 U12853 ( .ip1(\CORTEXM0DS_INST/u_logic/O7evx4 ), .ip2(n11525), .op(
        n11469) );
  buf_1 U12854 ( .ip(n11469), .op(n11554) );
  mux2_1 U12855 ( .ip1(\CORTEXM0DS_INST/vis_msp [7]), .ip2(n11577), .s(n11554), 
        .op(\CORTEXM0DS_INST/u_logic/Plivx4 ) );
  not_ab_or_c_or_d U12856 ( .ip1(n11549), .ip2(n12667), .ip3(n11252), .ip4(
        n11251), .op(n11253) );
  nand2_1 U12857 ( .ip1(n11254), .ip2(n11253), .op(n11578) );
  mux2_1 U12858 ( .ip1(\CORTEXM0DS_INST/vis_msp [0]), .ip2(n11578), .s(n11554), 
        .op(\CORTEXM0DS_INST/u_logic/Eqivx4 ) );
  inv_1 U12859 ( .ip(n11255), .op(n12660) );
  not_ab_or_c_or_d U12860 ( .ip1(n11549), .ip2(n12660), .ip3(n11257), .ip4(
        n11256), .op(n11258) );
  nand2_1 U12861 ( .ip1(n11259), .ip2(n11258), .op(n11579) );
  mux2_1 U12862 ( .ip1(\CORTEXM0DS_INST/vis_msp [8]), .ip2(n11579), .s(n11469), 
        .op(\CORTEXM0DS_INST/u_logic/Tuivx4 ) );
  inv_1 U12863 ( .ip(n11260), .op(n12661) );
  nor2_1 U12864 ( .ip1(n11511), .ip2(n11261), .op(n11262) );
  not_ab_or_c_or_d U12865 ( .ip1(n11549), .ip2(n12661), .ip3(n11263), .ip4(
        n11262), .op(n11268) );
  nor2_1 U12866 ( .ip1(n11434), .ip2(n11264), .op(n11266) );
  not_ab_or_c_or_d U12867 ( .ip1(n12137), .ip2(n11534), .ip3(n11266), .ip4(
        n11265), .op(n11267) );
  nand3_1 U12868 ( .ip1(n11268), .ip2(n11267), .ip3(n11451), .op(n11580) );
  mux2_1 U12869 ( .ip1(\CORTEXM0DS_INST/vis_msp [9]), .ip2(n11580), .s(n11469), 
        .op(\CORTEXM0DS_INST/u_logic/Izivx4 ) );
  nand2_1 U12870 ( .ip1(n12147), .ip2(n11534), .op(n11284) );
  inv_1 U12871 ( .ip(n11269), .op(n12662) );
  or2_1 U12872 ( .ip1(n12141), .ip2(n11270), .op(n11272) );
  or2_1 U12873 ( .ip1(n11511), .ip2(n11270), .op(n11271) );
  nand2_1 U12874 ( .ip1(n11272), .ip2(n11271), .op(n11273) );
  or2_1 U12875 ( .ip1(n11513), .ip2(n11273), .op(n11276) );
  inv_1 U12876 ( .ip(n12141), .op(n11274) );
  or2_1 U12877 ( .ip1(n11274), .ip2(n11273), .op(n11275) );
  nand2_1 U12878 ( .ip1(n11276), .ip2(n11275), .op(n11278) );
  or2_1 U12879 ( .ip1(n11277), .ip2(n11278), .op(n11280) );
  or2_1 U12880 ( .ip1(n11434), .ip2(n11278), .op(n11279) );
  nand2_1 U12881 ( .ip1(n11280), .ip2(n11279), .op(n11281) );
  not_ab_or_c_or_d U12882 ( .ip1(n11549), .ip2(n12662), .ip3(n11548), .ip4(
        n11281), .op(n11283) );
  nand3_1 U12883 ( .ip1(n11284), .ip2(n11283), .ip3(n11282), .op(n11581) );
  mux2_1 U12884 ( .ip1(\CORTEXM0DS_INST/vis_msp [10]), .ip2(n11581), .s(n11469), .op(\CORTEXM0DS_INST/u_logic/X3jvx4 ) );
  inv_1 U12885 ( .ip(n11285), .op(n12663) );
  nor2_1 U12886 ( .ip1(n11511), .ip2(n11286), .op(n11287) );
  not_ab_or_c_or_d U12887 ( .ip1(n11549), .ip2(n12663), .ip3(n11288), .ip4(
        n11287), .op(n11294) );
  nor2_1 U12888 ( .ip1(n11434), .ip2(n11289), .op(n11291) );
  not_ab_or_c_or_d U12889 ( .ip1(n11292), .ip2(n11534), .ip3(n11291), .ip4(
        n11290), .op(n11293) );
  nand3_1 U12890 ( .ip1(n11294), .ip2(n11293), .ip3(n11451), .op(n11582) );
  mux2_1 U12891 ( .ip1(\CORTEXM0DS_INST/vis_msp [11]), .ip2(n11582), .s(n11469), .op(\CORTEXM0DS_INST/u_logic/M8jvx4 ) );
  nor2_1 U12892 ( .ip1(n11295), .ip2(n11331), .op(n11296) );
  not_ab_or_c_or_d U12893 ( .ip1(n11298), .ip2(n11538), .ip3(n11297), .ip4(
        n11296), .op(n11304) );
  nor2_1 U12894 ( .ip1(n11434), .ip2(n11299), .op(n11301) );
  not_ab_or_c_or_d U12895 ( .ip1(n11302), .ip2(n11534), .ip3(n11301), .ip4(
        n11300), .op(n11303) );
  nand3_1 U12896 ( .ip1(n11304), .ip2(n11303), .ip3(n11451), .op(n11583) );
  mux2_1 U12897 ( .ip1(\CORTEXM0DS_INST/vis_msp [12]), .ip2(n11583), .s(n11469), .op(\CORTEXM0DS_INST/u_logic/Bdjvx4 ) );
  nand2_1 U12898 ( .ip1(n11305), .ip2(n11538), .op(n11315) );
  nand2_1 U12899 ( .ip1(n11451), .ip2(n11306), .op(n11528) );
  not_ab_or_c_or_d U12900 ( .ip1(n12162), .ip2(n11534), .ip3(n11528), .ip4(
        n11307), .op(n11314) );
  inv_1 U12901 ( .ip(n11308), .op(n11312) );
  nor2_1 U12902 ( .ip1(n11434), .ip2(n11309), .op(n11310) );
  not_ab_or_c_or_d U12903 ( .ip1(n11549), .ip2(n11312), .ip3(n11311), .ip4(
        n11310), .op(n11313) );
  nand3_1 U12904 ( .ip1(n11315), .ip2(n11314), .ip3(n11313), .op(n11584) );
  mux2_1 U12905 ( .ip1(\CORTEXM0DS_INST/vis_msp [14]), .ip2(n11584), .s(n11469), .op(\CORTEXM0DS_INST/u_logic/Qhjvx4 ) );
  inv_1 U12906 ( .ip(n11528), .op(n11377) );
  inv_1 U12907 ( .ip(n11316), .op(n12668) );
  nor2_1 U12908 ( .ip1(n11530), .ip2(n12168), .op(n11327) );
  or2_1 U12909 ( .ip1(n11511), .ip2(n11317), .op(n11318) );
  nand2_1 U12910 ( .ip1(n11323), .ip2(n11318), .op(n11320) );
  or2_1 U12911 ( .ip1(n11513), .ip2(n11320), .op(n11322) );
  inv_1 U12912 ( .ip(n11319), .op(n12171) );
  or2_1 U12913 ( .ip1(n12171), .ip2(n11320), .op(n11321) );
  nand2_1 U12914 ( .ip1(n11322), .ip2(n11321), .op(n11325) );
  nor2_1 U12915 ( .ip1(n11323), .ip2(n11537), .op(n11324) );
  nor2_1 U12916 ( .ip1(n11325), .ip2(n11324), .op(n11326) );
  not_ab_or_c_or_d U12917 ( .ip1(n11549), .ip2(n12668), .ip3(n11327), .ip4(
        n11326), .op(n11328) );
  nand3_1 U12918 ( .ip1(n11377), .ip2(n11329), .ip3(n11328), .op(n11585) );
  mux2_1 U12919 ( .ip1(\CORTEXM0DS_INST/vis_msp [15]), .ip2(n11585), .s(n11469), .op(\CORTEXM0DS_INST/u_logic/Fmjvx4 ) );
  nor2_1 U12920 ( .ip1(n11434), .ip2(n11330), .op(n11335) );
  nor2_1 U12921 ( .ip1(n12666), .ip2(n11331), .op(n11334) );
  nor2_1 U12922 ( .ip1(n11511), .ip2(n11332), .op(n11333) );
  nor4_1 U12923 ( .ip1(n11336), .ip2(n11335), .ip3(n11334), .ip4(n11333), .op(
        n11338) );
  nand2_1 U12924 ( .ip1(n12182), .ip2(n11534), .op(n11337) );
  nand4_1 U12925 ( .ip1(n11339), .ip2(n11377), .ip3(n11338), .ip4(n11337), 
        .op(n11586) );
  mux2_1 U12926 ( .ip1(\CORTEXM0DS_INST/vis_msp [16]), .ip2(n11586), .s(n11469), .op(\CORTEXM0DS_INST/u_logic/Uqjvx4 ) );
  or2_1 U12927 ( .ip1(n11511), .ip2(n11340), .op(n11341) );
  nand2_1 U12928 ( .ip1(n11346), .ip2(n11341), .op(n11343) );
  or2_1 U12929 ( .ip1(n11513), .ip2(n11343), .op(n11345) );
  inv_1 U12930 ( .ip(n11342), .op(n12192) );
  or2_1 U12931 ( .ip1(n12192), .ip2(n11343), .op(n11344) );
  nand2_1 U12932 ( .ip1(n11345), .ip2(n11344), .op(n11348) );
  nor2_1 U12933 ( .ip1(n11346), .ip2(n11537), .op(n11347) );
  nor2_1 U12934 ( .ip1(n11348), .ip2(n11347), .op(n11349) );
  not_ab_or_c_or_d U12935 ( .ip1(n11549), .ip2(n12672), .ip3(n11350), .ip4(
        n11349), .op(n11351) );
  nand3_1 U12936 ( .ip1(n11377), .ip2(n11352), .ip3(n11351), .op(n11587) );
  mux2_1 U12937 ( .ip1(\CORTEXM0DS_INST/vis_msp [17]), .ip2(n11587), .s(n11469), .op(\CORTEXM0DS_INST/u_logic/Jvjvx4 ) );
  nand2_1 U12938 ( .ip1(n11353), .ip2(n11538), .op(n11362) );
  nor3_1 U12939 ( .ip1(n11355), .ip2(n11528), .ip3(n11354), .op(n11361) );
  inv_1 U12940 ( .ip(n11356), .op(n12670) );
  nor2_1 U12941 ( .ip1(n11434), .ip2(n11357), .op(n11358) );
  not_ab_or_c_or_d U12942 ( .ip1(n11549), .ip2(n12670), .ip3(n11359), .ip4(
        n11358), .op(n11360) );
  nand3_1 U12943 ( .ip1(n11362), .ip2(n11361), .ip3(n11360), .op(n11588) );
  mux2_1 U12944 ( .ip1(\CORTEXM0DS_INST/vis_msp [18]), .ip2(n11588), .s(n11469), .op(\CORTEXM0DS_INST/u_logic/Yzjvx4 ) );
  or2_1 U12945 ( .ip1(n11366), .ip2(n11363), .op(n11365) );
  or2_1 U12946 ( .ip1(n11511), .ip2(n11363), .op(n11364) );
  nand2_1 U12947 ( .ip1(n11365), .ip2(n11364), .op(n11367) );
  or2_1 U12948 ( .ip1(n11513), .ip2(n11367), .op(n11369) );
  inv_1 U12949 ( .ip(n11366), .op(n12212) );
  or2_1 U12950 ( .ip1(n12212), .ip2(n11367), .op(n11368) );
  nand2_1 U12951 ( .ip1(n11369), .ip2(n11368), .op(n11371) );
  or2_1 U12952 ( .ip1(n11370), .ip2(n11371), .op(n11373) );
  or2_1 U12953 ( .ip1(n11434), .ip2(n11371), .op(n11372) );
  nand2_1 U12954 ( .ip1(n11373), .ip2(n11372), .op(n11375) );
  not_ab_or_c_or_d U12955 ( .ip1(n11549), .ip2(n12674), .ip3(n11375), .ip4(
        n11374), .op(n11378) );
  or2_1 U12956 ( .ip1(n12209), .ip2(n11530), .op(n11376) );
  nand3_1 U12957 ( .ip1(n11378), .ip2(n11377), .ip3(n11376), .op(n11589) );
  mux2_1 U12958 ( .ip1(\CORTEXM0DS_INST/vis_msp [19]), .ip2(n11589), .s(n11469), .op(\CORTEXM0DS_INST/u_logic/N4kvx4 ) );
  nand2_1 U12959 ( .ip1(n11379), .ip2(n11538), .op(n11387) );
  nor3_1 U12960 ( .ip1(n11381), .ip2(n11528), .ip3(n11380), .op(n11386) );
  nor2_1 U12961 ( .ip1(n11434), .ip2(n11382), .op(n11383) );
  not_ab_or_c_or_d U12962 ( .ip1(n11549), .ip2(n12676), .ip3(n11384), .ip4(
        n11383), .op(n11385) );
  nand3_1 U12963 ( .ip1(n11387), .ip2(n11386), .ip3(n11385), .op(n11590) );
  mux2_1 U12964 ( .ip1(\CORTEXM0DS_INST/vis_msp [20]), .ip2(n11590), .s(n11469), .op(\CORTEXM0DS_INST/u_logic/C9kvx4 ) );
  not_ab_or_c_or_d U12965 ( .ip1(n11390), .ip2(n11534), .ip3(n11389), .ip4(
        n11388), .op(n11394) );
  nand2_1 U12966 ( .ip1(n11549), .ip2(n12673), .op(n11393) );
  nand2_1 U12967 ( .ip1(n11548), .ip2(n11769), .op(n11392) );
  nand2_1 U12968 ( .ip1(n11481), .ip2(\CORTEXM0DS_INST/vis_ipsr [3]), .op(
        n11391) );
  nand4_1 U12969 ( .ip1(n11394), .ip2(n11393), .ip3(n11392), .ip4(n11391), 
        .op(n11591) );
  mux2_1 U12970 ( .ip1(\CORTEXM0DS_INST/vis_msp [1]), .ip2(n11591), .s(n11469), 
        .op(\CORTEXM0DS_INST/u_logic/Ydkvx4 ) );
  not_ab_or_c_or_d U12971 ( .ip1(n11397), .ip2(n11534), .ip3(n11396), .ip4(
        n11395), .op(n11398) );
  nand2_1 U12972 ( .ip1(n11399), .ip2(n11398), .op(n11592) );
  mux2_1 U12973 ( .ip1(\CORTEXM0DS_INST/vis_msp [2]), .ip2(n11592), .s(n11469), 
        .op(\CORTEXM0DS_INST/u_logic/Nikvx4 ) );
  not_ab_or_c_or_d U12974 ( .ip1(n12230), .ip2(n11534), .ip3(n11548), .ip4(
        n11400), .op(n11402) );
  nand3_1 U12975 ( .ip1(n11403), .ip2(n11402), .ip3(n11401), .op(n11593) );
  mux2_1 U12976 ( .ip1(\CORTEXM0DS_INST/vis_msp [3]), .ip2(n11593), .s(n11554), 
        .op(\CORTEXM0DS_INST/u_logic/Cnkvx4 ) );
  nor2_1 U12977 ( .ip1(n11511), .ip2(n11404), .op(n11405) );
  not_ab_or_c_or_d U12978 ( .ip1(n11549), .ip2(n12677), .ip3(n11548), .ip4(
        n11405), .op(n11411) );
  nand2_1 U12979 ( .ip1(n12243), .ip2(n11534), .op(n11410) );
  nand2_1 U12980 ( .ip1(n11434), .ip2(n11406), .op(n11407) );
  nand2_1 U12981 ( .ip1(n11408), .ip2(n11407), .op(n11409) );
  nand4_1 U12982 ( .ip1(n11412), .ip2(n11411), .ip3(n11410), .ip4(n11409), 
        .op(n11594) );
  mux2_1 U12983 ( .ip1(\CORTEXM0DS_INST/vis_msp [4]), .ip2(n11594), .s(n11469), 
        .op(\CORTEXM0DS_INST/u_logic/Rrkvx4 ) );
  nand2_1 U12984 ( .ip1(n11549), .ip2(n11413), .op(n11418) );
  nor3_1 U12985 ( .ip1(n11416), .ip2(n11415), .ip3(n11414), .op(n11417) );
  nand3_1 U12986 ( .ip1(n11418), .ip2(n11417), .ip3(n11451), .op(n11595) );
  mux2_1 U12987 ( .ip1(\CORTEXM0DS_INST/vis_msp [22]), .ip2(n11595), .s(n11469), .op(\CORTEXM0DS_INST/u_logic/Gwkvx4 ) );
  nor3_1 U12988 ( .ip1(n11421), .ip2(n11420), .ip3(n11419), .op(n11426) );
  nand2_1 U12989 ( .ip1(n11538), .ip2(n11422), .op(n11425) );
  nand2_1 U12990 ( .ip1(n11549), .ip2(n11423), .op(n11424) );
  nand4_1 U12991 ( .ip1(n11426), .ip2(n11451), .ip3(n11425), .ip4(n11424), 
        .op(n11596) );
  mux2_1 U12992 ( .ip1(\CORTEXM0DS_INST/vis_msp [23]), .ip2(n11596), .s(n11554), .op(\CORTEXM0DS_INST/u_logic/O0lvx4 ) );
  inv_1 U12993 ( .ip(n11427), .op(n11428) );
  or2_1 U12994 ( .ip1(n11513), .ip2(n11428), .op(n11430) );
  or2_1 U12995 ( .ip1(n11431), .ip2(n11428), .op(n11429) );
  nand2_1 U12996 ( .ip1(n11430), .ip2(n11429), .op(n11433) );
  nor2_1 U12997 ( .ip1(n11538), .ip2(n11431), .op(n11432) );
  not_ab_or_c_or_d U12998 ( .ip1(n11435), .ip2(n11434), .ip3(n11433), .ip4(
        n11432), .op(n11436) );
  not_ab_or_c_or_d U12999 ( .ip1(n11549), .ip2(n11437), .ip3(n11548), .ip4(
        n11436), .op(n11439) );
  nand3_1 U13000 ( .ip1(n11440), .ip2(n11439), .ip3(n11438), .op(n11597) );
  mux2_1 U13001 ( .ip1(\CORTEXM0DS_INST/vis_msp [24]), .ip2(n11597), .s(n11469), .op(\CORTEXM0DS_INST/u_logic/D5lvx4 ) );
  not_ab_or_c_or_d U13002 ( .ip1(n11549), .ip2(n11442), .ip3(n11548), .ip4(
        n11441), .op(n11444) );
  nand3_1 U13003 ( .ip1(n11445), .ip2(n11444), .ip3(n11443), .op(n11598) );
  mux2_1 U13004 ( .ip1(\CORTEXM0DS_INST/vis_msp [25]), .ip2(n11598), .s(n11469), .op(\CORTEXM0DS_INST/u_logic/S9lvx4 ) );
  not_ab_or_c_or_d U13005 ( .ip1(n11549), .ip2(n11447), .ip3(n11548), .ip4(
        n11446), .op(n11449) );
  nand3_1 U13006 ( .ip1(n11779), .ip2(n11449), .ip3(n11448), .op(n11601) );
  mux2_1 U13007 ( .ip1(\CORTEXM0DS_INST/vis_msp [27]), .ip2(n11601), .s(n11469), .op(\CORTEXM0DS_INST/u_logic/Helvx4 ) );
  nand2_1 U13008 ( .ip1(\CORTEXM0DS_INST/vis_apsr [2]), .ip2(n11450), .op(
        n11453) );
  nand3_1 U13009 ( .ip1(n11453), .ip2(n11452), .ip3(n11451), .op(n11454) );
  not_ab_or_c_or_d U13010 ( .ip1(n11549), .ip2(n11456), .ip3(n11455), .ip4(
        n11454), .op(n11460) );
  nand2_1 U13011 ( .ip1(n11457), .ip2(n11537), .op(n11458) );
  nand4_1 U13012 ( .ip1(n11631), .ip2(n11460), .ip3(n11459), .ip4(n11458), 
        .op(n11602) );
  mux2_1 U13013 ( .ip1(\CORTEXM0DS_INST/vis_msp [28]), .ip2(n11602), .s(n11554), .op(\CORTEXM0DS_INST/u_logic/Djlvx4 ) );
  inv_1 U13014 ( .ip(n11461), .op(n11462) );
  nand2_1 U13015 ( .ip1(n11462), .ip2(n11625), .op(n11617) );
  mux2_1 U13016 ( .ip1(\CORTEXM0DS_INST/vis_msp [29]), .ip2(n11617), .s(n11469), .op(\CORTEXM0DS_INST/u_logic/Rjlvx4 ) );
  inv_1 U13017 ( .ip(n11463), .op(n11468) );
  nand2_1 U13018 ( .ip1(n11549), .ip2(n11464), .op(n11465) );
  nand4_1 U13019 ( .ip1(n11468), .ip2(n11467), .ip3(n11466), .ip4(n11465), 
        .op(n11606) );
  mux2_1 U13020 ( .ip1(\CORTEXM0DS_INST/vis_msp [26]), .ip2(n11606), .s(n11469), .op(\CORTEXM0DS_INST/u_logic/Yjlvx4 ) );
  or2_1 U13021 ( .ip1(n11471), .ip2(n11470), .op(n11605) );
  mux2_1 U13022 ( .ip1(\CORTEXM0DS_INST/vis_msp [5]), .ip2(n11605), .s(n11554), 
        .op(\CORTEXM0DS_INST/u_logic/Fklvx4 ) );
  nand3_1 U13023 ( .ip1(n11496), .ip2(n11556), .ip3(n11557), .op(n11489) );
  buf_1 U13024 ( .ip(n11489), .op(n11560) );
  mux2_1 U13025 ( .ip1(n11577), .ip2(\CORTEXM0DS_INST/cm0_r12 [9]), .s(n11560), 
        .op(\CORTEXM0DS_INST/u_logic/Blivx4 ) );
  mux2_1 U13026 ( .ip1(n11578), .ip2(\CORTEXM0DS_INST/cm0_r12 [2]), .s(n11489), 
        .op(\CORTEXM0DS_INST/u_logic/Qpivx4 ) );
  mux2_1 U13027 ( .ip1(n11579), .ip2(\CORTEXM0DS_INST/cm0_r12 [10]), .s(n11489), .op(\CORTEXM0DS_INST/u_logic/Fuivx4 ) );
  mux2_1 U13028 ( .ip1(n11580), .ip2(\CORTEXM0DS_INST/cm0_r12 [11]), .s(n11489), .op(\CORTEXM0DS_INST/u_logic/Uyivx4 ) );
  mux2_1 U13029 ( .ip1(n11581), .ip2(\CORTEXM0DS_INST/cm0_r12 [12]), .s(n11489), .op(\CORTEXM0DS_INST/u_logic/J3jvx4 ) );
  mux2_1 U13030 ( .ip1(n11582), .ip2(\CORTEXM0DS_INST/cm0_r12 [13]), .s(n11489), .op(\CORTEXM0DS_INST/u_logic/Y7jvx4 ) );
  mux2_1 U13031 ( .ip1(n11583), .ip2(\CORTEXM0DS_INST/cm0_r12 [14]), .s(n11489), .op(\CORTEXM0DS_INST/u_logic/Ncjvx4 ) );
  mux2_1 U13032 ( .ip1(n11584), .ip2(\CORTEXM0DS_INST/cm0_r12 [16]), .s(n11489), .op(\CORTEXM0DS_INST/u_logic/Chjvx4 ) );
  mux2_1 U13033 ( .ip1(n11585), .ip2(\CORTEXM0DS_INST/cm0_r12 [17]), .s(n11489), .op(\CORTEXM0DS_INST/u_logic/Rljvx4 ) );
  mux2_1 U13034 ( .ip1(n11586), .ip2(\CORTEXM0DS_INST/cm0_r12 [18]), .s(n11560), .op(\CORTEXM0DS_INST/u_logic/Gqjvx4 ) );
  mux2_1 U13035 ( .ip1(n11587), .ip2(\CORTEXM0DS_INST/cm0_r12 [19]), .s(n11489), .op(\CORTEXM0DS_INST/u_logic/Vujvx4 ) );
  mux2_1 U13036 ( .ip1(n11588), .ip2(\CORTEXM0DS_INST/cm0_r12 [20]), .s(n11560), .op(\CORTEXM0DS_INST/u_logic/Kzjvx4 ) );
  mux2_1 U13037 ( .ip1(n11589), .ip2(\CORTEXM0DS_INST/cm0_r12 [21]), .s(n11489), .op(\CORTEXM0DS_INST/u_logic/Z3kvx4 ) );
  mux2_1 U13038 ( .ip1(n11590), .ip2(\CORTEXM0DS_INST/cm0_r12 [22]), .s(n11489), .op(\CORTEXM0DS_INST/u_logic/O8kvx4 ) );
  mux2_1 U13039 ( .ip1(n11591), .ip2(\CORTEXM0DS_INST/cm0_r12 [3]), .s(n11489), 
        .op(\CORTEXM0DS_INST/u_logic/Kdkvx4 ) );
  mux2_1 U13040 ( .ip1(n11592), .ip2(\CORTEXM0DS_INST/cm0_r12 [4]), .s(n11489), 
        .op(\CORTEXM0DS_INST/u_logic/Zhkvx4 ) );
  mux2_1 U13041 ( .ip1(n11593), .ip2(\CORTEXM0DS_INST/cm0_r12 [5]), .s(n11489), 
        .op(\CORTEXM0DS_INST/u_logic/Omkvx4 ) );
  mux2_1 U13042 ( .ip1(n11594), .ip2(\CORTEXM0DS_INST/cm0_r12 [6]), .s(n11489), 
        .op(\CORTEXM0DS_INST/u_logic/Drkvx4 ) );
  mux2_1 U13043 ( .ip1(n11595), .ip2(\CORTEXM0DS_INST/cm0_r12 [24]), .s(n11560), .op(\CORTEXM0DS_INST/u_logic/Svkvx4 ) );
  mux2_1 U13044 ( .ip1(n11596), .ip2(\CORTEXM0DS_INST/cm0_r12 [25]), .s(n11489), .op(\CORTEXM0DS_INST/u_logic/A0lvx4 ) );
  mux2_1 U13045 ( .ip1(n11597), .ip2(\CORTEXM0DS_INST/cm0_r12 [26]), .s(n11489), .op(\CORTEXM0DS_INST/u_logic/P4lvx4 ) );
  mux2_1 U13046 ( .ip1(n11598), .ip2(\CORTEXM0DS_INST/cm0_r12 [27]), .s(n11489), .op(\CORTEXM0DS_INST/u_logic/E9lvx4 ) );
  mux2_1 U13047 ( .ip1(n11601), .ip2(\CORTEXM0DS_INST/cm0_r12 [29]), .s(n11560), .op(\CORTEXM0DS_INST/u_logic/Tdlvx4 ) );
  mux2_1 U13048 ( .ip1(n11602), .ip2(\CORTEXM0DS_INST/cm0_r12 [30]), .s(n11489), .op(\CORTEXM0DS_INST/u_logic/Pilvx4 ) );
  nand2_1 U13049 ( .ip1(n11549), .ip2(n11472), .op(n11484) );
  inv_1 U13050 ( .ip(n11473), .op(n11474) );
  not_ab_or_c_or_d U13051 ( .ip1(n11476), .ip2(n11534), .ip3(n11475), .ip4(
        n11474), .op(n11483) );
  nor3_1 U13052 ( .ip1(n11479), .ip2(n11478), .ip3(n11477), .op(n11480) );
  not_ab_or_c_or_d U13053 ( .ip1(n11481), .ip2(\CORTEXM0DS_INST/vis_ipsr [0]), 
        .ip3(n11548), .ip4(n11480), .op(n11482) );
  nand3_1 U13054 ( .ip1(n11484), .ip2(n11483), .ip3(n11482), .op(n11603) );
  mux2_1 U13055 ( .ip1(n11603), .ip2(\CORTEXM0DS_INST/cm0_r12 [0]), .s(n11489), 
        .op(\CORTEXM0DS_INST/u_logic/Mrlvx4 ) );
  not_ab_or_c_or_d U13056 ( .ip1(n11549), .ip2(n12669), .ip3(n11486), .ip4(
        n11485), .op(n11488) );
  nand2_1 U13057 ( .ip1(n11488), .ip2(n11487), .op(n11604) );
  mux2_1 U13058 ( .ip1(n11604), .ip2(\CORTEXM0DS_INST/cm0_r12 [1]), .s(n11489), 
        .op(\CORTEXM0DS_INST/u_logic/Trlvx4 ) );
  mux2_1 U13059 ( .ip1(n11605), .ip2(\CORTEXM0DS_INST/cm0_r12 [7]), .s(n11560), 
        .op(\CORTEXM0DS_INST/u_logic/Aslvx4 ) );
  mux2_1 U13060 ( .ip1(n11606), .ip2(\CORTEXM0DS_INST/cm0_r12 [28]), .s(n11560), .op(\CORTEXM0DS_INST/u_logic/Hslvx4 ) );
  mux2_1 U13061 ( .ip1(n11617), .ip2(\CORTEXM0DS_INST/cm0_r12 [31]), .s(n11560), .op(\CORTEXM0DS_INST/u_logic/Oslvx4 ) );
  inv_1 U13062 ( .ip(n11496), .op(n11555) );
  nand2_1 U13063 ( .ip1(n11555), .ip2(n11490), .op(n11504) );
  nand2_1 U13064 ( .ip1(n11492), .ip2(n11491), .op(n11563) );
  nor2_1 U13065 ( .ip1(n11504), .ip2(n11563), .op(n11493) );
  mux2_1 U13066 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [9]), .ip2(n11577), .s(n11493), 
        .op(\CORTEXM0DS_INST/u_logic/Ukivx4 ) );
  buf_1 U13067 ( .ip(n11493), .op(n11561) );
  mux2_1 U13068 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [2]), .ip2(n11578), .s(n11561), 
        .op(\CORTEXM0DS_INST/u_logic/Jpivx4 ) );
  mux2_1 U13069 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [10]), .ip2(n11579), .s(n11493), .op(\CORTEXM0DS_INST/u_logic/Ytivx4 ) );
  mux2_1 U13070 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [11]), .ip2(n11580), .s(n11493), .op(\CORTEXM0DS_INST/u_logic/Nyivx4 ) );
  mux2_1 U13071 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [12]), .ip2(n11581), .s(n11493), .op(\CORTEXM0DS_INST/u_logic/C3jvx4 ) );
  mux2_1 U13072 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [13]), .ip2(n11582), .s(n11493), .op(\CORTEXM0DS_INST/u_logic/R7jvx4 ) );
  mux2_1 U13073 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [14]), .ip2(n11583), .s(n11493), .op(\CORTEXM0DS_INST/u_logic/Gcjvx4 ) );
  mux2_1 U13074 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [16]), .ip2(n11584), .s(n11493), .op(\CORTEXM0DS_INST/u_logic/Vgjvx4 ) );
  mux2_1 U13075 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [17]), .ip2(n11585), .s(n11493), .op(\CORTEXM0DS_INST/u_logic/Kljvx4 ) );
  mux2_1 U13076 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [18]), .ip2(n11586), .s(n11493), .op(\CORTEXM0DS_INST/u_logic/Zpjvx4 ) );
  mux2_1 U13077 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [19]), .ip2(n11587), .s(n11493), .op(\CORTEXM0DS_INST/u_logic/Oujvx4 ) );
  mux2_1 U13078 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [20]), .ip2(n11588), .s(n11493), .op(\CORTEXM0DS_INST/u_logic/Dzjvx4 ) );
  mux2_1 U13079 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [21]), .ip2(n11589), .s(n11561), .op(\CORTEXM0DS_INST/u_logic/S3kvx4 ) );
  mux2_1 U13080 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [22]), .ip2(n11590), .s(n11493), .op(\CORTEXM0DS_INST/u_logic/H8kvx4 ) );
  mux2_1 U13081 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [3]), .ip2(n11591), .s(n11493), 
        .op(\CORTEXM0DS_INST/u_logic/Ddkvx4 ) );
  mux2_1 U13082 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [4]), .ip2(n11592), .s(n11493), 
        .op(\CORTEXM0DS_INST/u_logic/Shkvx4 ) );
  mux2_1 U13083 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [5]), .ip2(n11593), .s(n11561), 
        .op(\CORTEXM0DS_INST/u_logic/Hmkvx4 ) );
  mux2_1 U13084 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [6]), .ip2(n11594), .s(n11493), 
        .op(\CORTEXM0DS_INST/u_logic/Wqkvx4 ) );
  mux2_1 U13085 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [24]), .ip2(n11595), .s(n11493), .op(\CORTEXM0DS_INST/u_logic/Lvkvx4 ) );
  mux2_1 U13086 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [25]), .ip2(n11596), .s(n11493), .op(\CORTEXM0DS_INST/u_logic/Tzkvx4 ) );
  mux2_1 U13087 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [26]), .ip2(n11597), .s(n11493), .op(\CORTEXM0DS_INST/u_logic/I4lvx4 ) );
  mux2_1 U13088 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [27]), .ip2(n11598), .s(n11493), .op(\CORTEXM0DS_INST/u_logic/X8lvx4 ) );
  mux2_1 U13089 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [29]), .ip2(n11601), .s(n11493), .op(\CORTEXM0DS_INST/u_logic/Mdlvx4 ) );
  mux2_1 U13090 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [30]), .ip2(n11602), .s(n11493), .op(\CORTEXM0DS_INST/u_logic/Iilvx4 ) );
  mux2_1 U13091 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [0]), .ip2(n11603), .s(n11561), 
        .op(\CORTEXM0DS_INST/u_logic/Dqlvx4 ) );
  mux2_1 U13092 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [1]), .ip2(n11604), .s(n11561), 
        .op(\CORTEXM0DS_INST/u_logic/Kqlvx4 ) );
  mux2_1 U13093 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [7]), .ip2(n11605), .s(n11561), 
        .op(\CORTEXM0DS_INST/u_logic/Rqlvx4 ) );
  mux2_1 U13094 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [28]), .ip2(n11606), .s(n11561), .op(\CORTEXM0DS_INST/u_logic/Yqlvx4 ) );
  mux2_1 U13095 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [31]), .ip2(n11617), .s(n11561), .op(\CORTEXM0DS_INST/u_logic/Frlvx4 ) );
  inv_1 U13096 ( .ip(n11494), .op(n11506) );
  nor2_1 U13097 ( .ip1(n11506), .ip2(n11563), .op(n11495) );
  mux2_1 U13098 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [9]), .ip2(n11577), .s(n11495), 
        .op(\CORTEXM0DS_INST/u_logic/Gkivx4 ) );
  buf_1 U13099 ( .ip(n11495), .op(n11566) );
  mux2_1 U13100 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [2]), .ip2(n11578), .s(n11566), 
        .op(\CORTEXM0DS_INST/u_logic/Voivx4 ) );
  mux2_1 U13101 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [10]), .ip2(n11579), .s(n11495), .op(\CORTEXM0DS_INST/u_logic/Ktivx4 ) );
  mux2_1 U13102 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [11]), .ip2(n11580), .s(n11495), .op(\CORTEXM0DS_INST/u_logic/Zxivx4 ) );
  mux2_1 U13103 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [12]), .ip2(n11581), .s(n11495), .op(\CORTEXM0DS_INST/u_logic/O2jvx4 ) );
  mux2_1 U13104 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [13]), .ip2(n11582), .s(n11495), .op(\CORTEXM0DS_INST/u_logic/D7jvx4 ) );
  mux2_1 U13105 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [14]), .ip2(n11583), .s(n11495), .op(\CORTEXM0DS_INST/u_logic/Sbjvx4 ) );
  mux2_1 U13106 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [16]), .ip2(n11584), .s(n11495), .op(\CORTEXM0DS_INST/u_logic/Hgjvx4 ) );
  mux2_1 U13107 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [17]), .ip2(n11585), .s(n11495), .op(\CORTEXM0DS_INST/u_logic/Wkjvx4 ) );
  mux2_1 U13108 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [18]), .ip2(n11586), .s(n11495), .op(\CORTEXM0DS_INST/u_logic/Lpjvx4 ) );
  mux2_1 U13109 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [19]), .ip2(n11587), .s(n11495), .op(\CORTEXM0DS_INST/u_logic/Aujvx4 ) );
  mux2_1 U13110 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [20]), .ip2(n11588), .s(n11495), .op(\CORTEXM0DS_INST/u_logic/Pyjvx4 ) );
  mux2_1 U13111 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [21]), .ip2(n11589), .s(n11566), .op(\CORTEXM0DS_INST/u_logic/E3kvx4 ) );
  mux2_1 U13112 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [22]), .ip2(n11590), .s(n11495), .op(\CORTEXM0DS_INST/u_logic/T7kvx4 ) );
  mux2_1 U13113 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [3]), .ip2(n11591), .s(n11495), 
        .op(\CORTEXM0DS_INST/u_logic/Pckvx4 ) );
  mux2_1 U13114 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [4]), .ip2(n11592), .s(n11495), 
        .op(\CORTEXM0DS_INST/u_logic/Ehkvx4 ) );
  mux2_1 U13115 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [5]), .ip2(n11593), .s(n11566), 
        .op(\CORTEXM0DS_INST/u_logic/Tlkvx4 ) );
  mux2_1 U13116 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [6]), .ip2(n11594), .s(n11495), 
        .op(\CORTEXM0DS_INST/u_logic/Iqkvx4 ) );
  mux2_1 U13117 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [24]), .ip2(n11595), .s(n11495), .op(\CORTEXM0DS_INST/u_logic/Xukvx4 ) );
  mux2_1 U13118 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [25]), .ip2(n11596), .s(n11495), .op(\CORTEXM0DS_INST/u_logic/Fzkvx4 ) );
  mux2_1 U13119 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [26]), .ip2(n11597), .s(n11495), .op(\CORTEXM0DS_INST/u_logic/U3lvx4 ) );
  mux2_1 U13120 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [27]), .ip2(n11598), .s(n11495), .op(\CORTEXM0DS_INST/u_logic/J8lvx4 ) );
  mux2_1 U13121 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [29]), .ip2(n11601), .s(n11495), .op(\CORTEXM0DS_INST/u_logic/Yclvx4 ) );
  mux2_1 U13122 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [30]), .ip2(n11602), .s(n11495), .op(\CORTEXM0DS_INST/u_logic/Uhlvx4 ) );
  mux2_1 U13123 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [0]), .ip2(n11603), .s(n11566), 
        .op(\CORTEXM0DS_INST/u_logic/Lnlvx4 ) );
  mux2_1 U13124 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [1]), .ip2(n11604), .s(n11566), 
        .op(\CORTEXM0DS_INST/u_logic/Snlvx4 ) );
  mux2_1 U13125 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [7]), .ip2(n11605), .s(n11566), 
        .op(\CORTEXM0DS_INST/u_logic/Znlvx4 ) );
  mux2_1 U13126 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [28]), .ip2(n11606), .s(n11566), .op(\CORTEXM0DS_INST/u_logic/Golvx4 ) );
  mux2_1 U13127 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [31]), .ip2(n11617), .s(n11566), .op(\CORTEXM0DS_INST/u_logic/Nolvx4 ) );
  nand2_1 U13128 ( .ip1(n11496), .ip2(n11556), .op(n11508) );
  nor2_1 U13129 ( .ip1(n11508), .ip2(n11563), .op(n11497) );
  mux2_1 U13130 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [9]), .ip2(n11577), .s(n11497), 
        .op(\CORTEXM0DS_INST/u_logic/Zjivx4 ) );
  buf_1 U13131 ( .ip(n11497), .op(n11567) );
  mux2_1 U13132 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [2]), .ip2(n11578), .s(n11567), 
        .op(\CORTEXM0DS_INST/u_logic/Ooivx4 ) );
  mux2_1 U13133 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [10]), .ip2(n11579), .s(n11497), .op(\CORTEXM0DS_INST/u_logic/Dtivx4 ) );
  mux2_1 U13134 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [11]), .ip2(n11580), .s(n11497), .op(\CORTEXM0DS_INST/u_logic/Sxivx4 ) );
  mux2_1 U13135 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [12]), .ip2(n11581), .s(n11497), .op(\CORTEXM0DS_INST/u_logic/H2jvx4 ) );
  mux2_1 U13136 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [13]), .ip2(n11582), .s(n11497), .op(\CORTEXM0DS_INST/u_logic/W6jvx4 ) );
  mux2_1 U13137 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [14]), .ip2(n11583), .s(n11497), .op(\CORTEXM0DS_INST/u_logic/Lbjvx4 ) );
  mux2_1 U13138 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [16]), .ip2(n11584), .s(n11497), .op(\CORTEXM0DS_INST/u_logic/Agjvx4 ) );
  mux2_1 U13139 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [17]), .ip2(n11585), .s(n11497), .op(\CORTEXM0DS_INST/u_logic/Pkjvx4 ) );
  mux2_1 U13140 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [18]), .ip2(n11586), .s(n11497), .op(\CORTEXM0DS_INST/u_logic/Epjvx4 ) );
  mux2_1 U13141 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [19]), .ip2(n11587), .s(n11497), .op(\CORTEXM0DS_INST/u_logic/Ttjvx4 ) );
  mux2_1 U13142 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [20]), .ip2(n11588), .s(n11497), .op(\CORTEXM0DS_INST/u_logic/Iyjvx4 ) );
  mux2_1 U13143 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [21]), .ip2(n11589), .s(n11567), .op(\CORTEXM0DS_INST/u_logic/X2kvx4 ) );
  mux2_1 U13144 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [22]), .ip2(n11590), .s(n11497), .op(\CORTEXM0DS_INST/u_logic/M7kvx4 ) );
  mux2_1 U13145 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [3]), .ip2(n11591), .s(n11497), 
        .op(\CORTEXM0DS_INST/u_logic/Ickvx4 ) );
  mux2_1 U13146 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [4]), .ip2(n11592), .s(n11497), 
        .op(\CORTEXM0DS_INST/u_logic/Xgkvx4 ) );
  mux2_1 U13147 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [5]), .ip2(n11593), .s(n11567), 
        .op(\CORTEXM0DS_INST/u_logic/Mlkvx4 ) );
  mux2_1 U13148 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [6]), .ip2(n11594), .s(n11497), 
        .op(\CORTEXM0DS_INST/u_logic/Bqkvx4 ) );
  mux2_1 U13149 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [24]), .ip2(n11595), .s(n11497), .op(\CORTEXM0DS_INST/u_logic/Qukvx4 ) );
  mux2_1 U13150 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [25]), .ip2(n11596), .s(n11567), .op(\CORTEXM0DS_INST/u_logic/Yykvx4 ) );
  mux2_1 U13151 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [26]), .ip2(n11597), .s(n11497), .op(\CORTEXM0DS_INST/u_logic/N3lvx4 ) );
  mux2_1 U13152 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [27]), .ip2(n11598), .s(n11497), .op(\CORTEXM0DS_INST/u_logic/C8lvx4 ) );
  mux2_1 U13153 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [29]), .ip2(n11601), .s(n11497), .op(\CORTEXM0DS_INST/u_logic/Rclvx4 ) );
  mux2_1 U13154 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [30]), .ip2(n11602), .s(n11567), .op(\CORTEXM0DS_INST/u_logic/Nhlvx4 ) );
  mux2_1 U13155 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [0]), .ip2(n11603), .s(n11497), 
        .op(\CORTEXM0DS_INST/u_logic/Cmlvx4 ) );
  mux2_1 U13156 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [1]), .ip2(n11604), .s(n11497), 
        .op(\CORTEXM0DS_INST/u_logic/Jmlvx4 ) );
  mux2_1 U13157 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [7]), .ip2(n11605), .s(n11567), 
        .op(\CORTEXM0DS_INST/u_logic/Qmlvx4 ) );
  mux2_1 U13158 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [28]), .ip2(n11606), .s(n11567), .op(\CORTEXM0DS_INST/u_logic/Xmlvx4 ) );
  mux2_1 U13159 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [31]), .ip2(n11617), .s(n11567), .op(\CORTEXM0DS_INST/u_logic/Enlvx4 ) );
  nand2_1 U13160 ( .ip1(n11503), .ip2(n11501), .op(n11569) );
  nor2_1 U13161 ( .ip1(n11504), .ip2(n11569), .op(n11498) );
  mux2_1 U13162 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [9]), .ip2(n11577), .s(n11498), 
        .op(\CORTEXM0DS_INST/u_logic/Sjivx4 ) );
  mux2_1 U13163 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [2]), .ip2(n11578), .s(n11498), 
        .op(\CORTEXM0DS_INST/u_logic/Hoivx4 ) );
  mux2_1 U13164 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [10]), .ip2(n11579), .s(n11498), .op(\CORTEXM0DS_INST/u_logic/Wsivx4 ) );
  mux2_1 U13165 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [11]), .ip2(n11580), .s(n11498), .op(\CORTEXM0DS_INST/u_logic/Lxivx4 ) );
  mux2_1 U13166 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [12]), .ip2(n11581), .s(n11498), .op(\CORTEXM0DS_INST/u_logic/A2jvx4 ) );
  mux2_1 U13167 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [13]), .ip2(n11582), .s(n11498), .op(\CORTEXM0DS_INST/u_logic/P6jvx4 ) );
  mux2_1 U13168 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [14]), .ip2(n11583), .s(n11498), .op(\CORTEXM0DS_INST/u_logic/Ebjvx4 ) );
  mux2_1 U13169 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [16]), .ip2(n11584), .s(n11498), .op(\CORTEXM0DS_INST/u_logic/Tfjvx4 ) );
  mux2_1 U13170 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [17]), .ip2(n11585), .s(n11498), .op(\CORTEXM0DS_INST/u_logic/Ikjvx4 ) );
  mux2_1 U13171 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [18]), .ip2(n11586), .s(n11498), .op(\CORTEXM0DS_INST/u_logic/Xojvx4 ) );
  mux2_1 U13172 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [19]), .ip2(n11587), .s(n11498), .op(\CORTEXM0DS_INST/u_logic/Mtjvx4 ) );
  buf_1 U13173 ( .ip(n11498), .op(n11568) );
  mux2_1 U13174 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [20]), .ip2(n11588), .s(n11568), .op(\CORTEXM0DS_INST/u_logic/Byjvx4 ) );
  mux2_1 U13175 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [21]), .ip2(n11589), .s(n11568), .op(\CORTEXM0DS_INST/u_logic/Q2kvx4 ) );
  mux2_1 U13176 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [22]), .ip2(n11590), .s(n11498), .op(\CORTEXM0DS_INST/u_logic/F7kvx4 ) );
  mux2_1 U13177 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [3]), .ip2(n11591), .s(n11498), 
        .op(\CORTEXM0DS_INST/u_logic/Bckvx4 ) );
  mux2_1 U13178 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [4]), .ip2(n11592), .s(n11498), 
        .op(\CORTEXM0DS_INST/u_logic/Qgkvx4 ) );
  mux2_1 U13179 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [5]), .ip2(n11593), .s(n11498), 
        .op(\CORTEXM0DS_INST/u_logic/Flkvx4 ) );
  mux2_1 U13180 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [6]), .ip2(n11594), .s(n11498), 
        .op(\CORTEXM0DS_INST/u_logic/Upkvx4 ) );
  mux2_1 U13181 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [24]), .ip2(n11595), .s(n11498), .op(\CORTEXM0DS_INST/u_logic/Jukvx4 ) );
  mux2_1 U13182 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [25]), .ip2(n11596), .s(n11568), .op(\CORTEXM0DS_INST/u_logic/Rykvx4 ) );
  mux2_1 U13183 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [26]), .ip2(n11597), .s(n11498), .op(\CORTEXM0DS_INST/u_logic/G3lvx4 ) );
  mux2_1 U13184 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [27]), .ip2(n11598), .s(n11498), .op(\CORTEXM0DS_INST/u_logic/V7lvx4 ) );
  mux2_1 U13185 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [29]), .ip2(n11601), .s(n11568), .op(\CORTEXM0DS_INST/u_logic/Kclvx4 ) );
  mux2_1 U13186 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [30]), .ip2(n11602), .s(n11568), .op(\CORTEXM0DS_INST/u_logic/Ghlvx4 ) );
  mux2_1 U13187 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [0]), .ip2(n11603), .s(n11498), 
        .op(\CORTEXM0DS_INST/u_logic/Eulvx4 ) );
  mux2_1 U13188 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [1]), .ip2(n11604), .s(n11498), 
        .op(\CORTEXM0DS_INST/u_logic/Lulvx4 ) );
  mux2_1 U13189 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [7]), .ip2(n11605), .s(n11568), 
        .op(\CORTEXM0DS_INST/u_logic/Sulvx4 ) );
  mux2_1 U13190 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [28]), .ip2(n11606), .s(n11568), .op(\CORTEXM0DS_INST/u_logic/Zulvx4 ) );
  mux2_1 U13191 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [31]), .ip2(n11617), .s(n11568), .op(\CORTEXM0DS_INST/u_logic/Gvlvx4 ) );
  nor2_1 U13192 ( .ip1(n11506), .ip2(n11569), .op(n11499) );
  mux2_1 U13193 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [9]), .ip2(n11577), .s(n11499), 
        .op(\CORTEXM0DS_INST/u_logic/Ejivx4 ) );
  buf_1 U13194 ( .ip(n11499), .op(n11572) );
  mux2_1 U13195 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [2]), .ip2(n11578), .s(n11572), 
        .op(\CORTEXM0DS_INST/u_logic/Tnivx4 ) );
  mux2_1 U13196 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [10]), .ip2(n11579), .s(n11499), .op(\CORTEXM0DS_INST/u_logic/Isivx4 ) );
  mux2_1 U13197 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [11]), .ip2(n11580), .s(n11499), .op(\CORTEXM0DS_INST/u_logic/Xwivx4 ) );
  mux2_1 U13198 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [12]), .ip2(n11581), .s(n11499), .op(\CORTEXM0DS_INST/u_logic/M1jvx4 ) );
  mux2_1 U13199 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [13]), .ip2(n11582), .s(n11499), .op(\CORTEXM0DS_INST/u_logic/B6jvx4 ) );
  mux2_1 U13200 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [14]), .ip2(n11583), .s(n11499), .op(\CORTEXM0DS_INST/u_logic/Qajvx4 ) );
  mux2_1 U13201 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [16]), .ip2(n11584), .s(n11499), .op(\CORTEXM0DS_INST/u_logic/Ffjvx4 ) );
  mux2_1 U13202 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [17]), .ip2(n11585), .s(n11499), .op(\CORTEXM0DS_INST/u_logic/Ujjvx4 ) );
  mux2_1 U13203 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [18]), .ip2(n11586), .s(n11499), .op(\CORTEXM0DS_INST/u_logic/Jojvx4 ) );
  mux2_1 U13204 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [19]), .ip2(n11587), .s(n11499), .op(\CORTEXM0DS_INST/u_logic/Ysjvx4 ) );
  mux2_1 U13205 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [20]), .ip2(n11588), .s(n11499), .op(\CORTEXM0DS_INST/u_logic/Nxjvx4 ) );
  mux2_1 U13206 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [21]), .ip2(n11589), .s(n11572), .op(\CORTEXM0DS_INST/u_logic/C2kvx4 ) );
  mux2_1 U13207 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [22]), .ip2(n11590), .s(n11499), .op(\CORTEXM0DS_INST/u_logic/R6kvx4 ) );
  mux2_1 U13208 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [3]), .ip2(n11591), .s(n11499), 
        .op(\CORTEXM0DS_INST/u_logic/Nbkvx4 ) );
  mux2_1 U13209 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [4]), .ip2(n11592), .s(n11499), 
        .op(\CORTEXM0DS_INST/u_logic/Cgkvx4 ) );
  mux2_1 U13210 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [5]), .ip2(n11593), .s(n11572), 
        .op(\CORTEXM0DS_INST/u_logic/Rkkvx4 ) );
  mux2_1 U13211 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [6]), .ip2(n11594), .s(n11499), 
        .op(\CORTEXM0DS_INST/u_logic/Gpkvx4 ) );
  mux2_1 U13212 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [24]), .ip2(n11595), .s(n11499), .op(\CORTEXM0DS_INST/u_logic/Vtkvx4 ) );
  mux2_1 U13213 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [25]), .ip2(n11596), .s(n11572), .op(\CORTEXM0DS_INST/u_logic/Dykvx4 ) );
  mux2_1 U13214 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [26]), .ip2(n11597), .s(n11499), .op(\CORTEXM0DS_INST/u_logic/S2lvx4 ) );
  mux2_1 U13215 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [27]), .ip2(n11598), .s(n11499), .op(\CORTEXM0DS_INST/u_logic/H7lvx4 ) );
  mux2_1 U13216 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [29]), .ip2(n11601), .s(n11499), .op(\CORTEXM0DS_INST/u_logic/Wblvx4 ) );
  mux2_1 U13217 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [30]), .ip2(n11602), .s(n11572), .op(\CORTEXM0DS_INST/u_logic/Sglvx4 ) );
  mux2_1 U13218 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [0]), .ip2(n11603), .s(n11499), 
        .op(\CORTEXM0DS_INST/u_logic/Wwlvx4 ) );
  mux2_1 U13219 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [1]), .ip2(n11604), .s(n11499), 
        .op(\CORTEXM0DS_INST/u_logic/Dxlvx4 ) );
  mux2_1 U13220 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [7]), .ip2(n11605), .s(n11572), 
        .op(\CORTEXM0DS_INST/u_logic/Kxlvx4 ) );
  mux2_1 U13221 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [28]), .ip2(n11606), .s(n11572), .op(\CORTEXM0DS_INST/u_logic/Rxlvx4 ) );
  mux2_1 U13222 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [31]), .ip2(n11617), .s(n11572), .op(\CORTEXM0DS_INST/u_logic/Yxlvx4 ) );
  nor2_1 U13223 ( .ip1(n11508), .ip2(n11569), .op(n11500) );
  mux2_1 U13224 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [9]), .ip2(n11577), .s(n11500), 
        .op(\CORTEXM0DS_INST/u_logic/Xiivx4 ) );
  mux2_1 U13225 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [2]), .ip2(n11578), .s(n11500), 
        .op(\CORTEXM0DS_INST/u_logic/Mnivx4 ) );
  mux2_1 U13226 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [10]), .ip2(n11579), .s(n11500), .op(\CORTEXM0DS_INST/u_logic/Bsivx4 ) );
  mux2_1 U13227 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [11]), .ip2(n11580), .s(n11500), .op(\CORTEXM0DS_INST/u_logic/Qwivx4 ) );
  mux2_1 U13228 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [12]), .ip2(n11581), .s(n11500), .op(\CORTEXM0DS_INST/u_logic/F1jvx4 ) );
  mux2_1 U13229 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [13]), .ip2(n11582), .s(n11500), .op(\CORTEXM0DS_INST/u_logic/U5jvx4 ) );
  mux2_1 U13230 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [14]), .ip2(n11583), .s(n11500), .op(\CORTEXM0DS_INST/u_logic/Jajvx4 ) );
  mux2_1 U13231 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [16]), .ip2(n11584), .s(n11500), .op(\CORTEXM0DS_INST/u_logic/Yejvx4 ) );
  mux2_1 U13232 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [17]), .ip2(n11585), .s(n11500), .op(\CORTEXM0DS_INST/u_logic/Njjvx4 ) );
  mux2_1 U13233 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [18]), .ip2(n11586), .s(n11500), .op(\CORTEXM0DS_INST/u_logic/Cojvx4 ) );
  mux2_1 U13234 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [19]), .ip2(n11587), .s(n11500), .op(\CORTEXM0DS_INST/u_logic/Rsjvx4 ) );
  buf_1 U13235 ( .ip(n11500), .op(n11573) );
  mux2_1 U13236 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [20]), .ip2(n11588), .s(n11573), .op(\CORTEXM0DS_INST/u_logic/Gxjvx4 ) );
  mux2_1 U13237 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [21]), .ip2(n11589), .s(n11573), .op(\CORTEXM0DS_INST/u_logic/V1kvx4 ) );
  mux2_1 U13238 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [22]), .ip2(n11590), .s(n11500), .op(\CORTEXM0DS_INST/u_logic/K6kvx4 ) );
  mux2_1 U13239 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [3]), .ip2(n11591), .s(n11500), 
        .op(\CORTEXM0DS_INST/u_logic/Gbkvx4 ) );
  mux2_1 U13240 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [4]), .ip2(n11592), .s(n11500), 
        .op(\CORTEXM0DS_INST/u_logic/Vfkvx4 ) );
  mux2_1 U13241 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [5]), .ip2(n11593), .s(n11500), 
        .op(\CORTEXM0DS_INST/u_logic/Kkkvx4 ) );
  mux2_1 U13242 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [6]), .ip2(n11594), .s(n11500), 
        .op(\CORTEXM0DS_INST/u_logic/Zokvx4 ) );
  mux2_1 U13243 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [24]), .ip2(n11595), .s(n11500), .op(\CORTEXM0DS_INST/u_logic/Otkvx4 ) );
  mux2_1 U13244 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [25]), .ip2(n11596), .s(n11573), .op(\CORTEXM0DS_INST/u_logic/Wxkvx4 ) );
  mux2_1 U13245 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [26]), .ip2(n11597), .s(n11500), .op(\CORTEXM0DS_INST/u_logic/L2lvx4 ) );
  mux2_1 U13246 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [27]), .ip2(n11598), .s(n11500), .op(\CORTEXM0DS_INST/u_logic/A7lvx4 ) );
  mux2_1 U13247 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [29]), .ip2(n11601), .s(n11573), .op(\CORTEXM0DS_INST/u_logic/Pblvx4 ) );
  mux2_1 U13248 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [30]), .ip2(n11602), .s(n11573), .op(\CORTEXM0DS_INST/u_logic/Lglvx4 ) );
  mux2_1 U13249 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [0]), .ip2(n11603), .s(n11500), 
        .op(\CORTEXM0DS_INST/u_logic/Fylvx4 ) );
  mux2_1 U13250 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [1]), .ip2(n11604), .s(n11500), 
        .op(\CORTEXM0DS_INST/u_logic/Mylvx4 ) );
  mux2_1 U13251 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [7]), .ip2(n11605), .s(n11573), 
        .op(\CORTEXM0DS_INST/u_logic/Tylvx4 ) );
  mux2_1 U13252 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [28]), .ip2(n11606), .s(n11573), .op(\CORTEXM0DS_INST/u_logic/Azlvx4 ) );
  mux2_1 U13253 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [31]), .ip2(n11617), .s(n11573), .op(\CORTEXM0DS_INST/u_logic/Hzlvx4 ) );
  inv_1 U13254 ( .ip(n11501), .op(n11502) );
  nand2_1 U13255 ( .ip1(n11503), .ip2(n11502), .op(n11576) );
  nor2_1 U13256 ( .ip1(n11504), .ip2(n11576), .op(n11505) );
  mux2_1 U13257 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [9]), .ip2(n11577), .s(n11505), 
        .op(\CORTEXM0DS_INST/u_logic/Qiivx4 ) );
  buf_1 U13258 ( .ip(n11505), .op(n11574) );
  mux2_1 U13259 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [2]), .ip2(n11578), .s(n11574), 
        .op(\CORTEXM0DS_INST/u_logic/Fnivx4 ) );
  mux2_1 U13260 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [10]), .ip2(n11579), .s(n11505), .op(\CORTEXM0DS_INST/u_logic/Urivx4 ) );
  mux2_1 U13261 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [11]), .ip2(n11580), .s(n11505), .op(\CORTEXM0DS_INST/u_logic/Jwivx4 ) );
  mux2_1 U13262 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [12]), .ip2(n11581), .s(n11505), .op(\CORTEXM0DS_INST/u_logic/Y0jvx4 ) );
  mux2_1 U13263 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [13]), .ip2(n11582), .s(n11505), .op(\CORTEXM0DS_INST/u_logic/N5jvx4 ) );
  mux2_1 U13264 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [14]), .ip2(n11583), .s(n11505), .op(\CORTEXM0DS_INST/u_logic/Cajvx4 ) );
  mux2_1 U13265 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [16]), .ip2(n11584), .s(n11505), .op(\CORTEXM0DS_INST/u_logic/Rejvx4 ) );
  mux2_1 U13266 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [17]), .ip2(n11585), .s(n11505), .op(\CORTEXM0DS_INST/u_logic/Gjjvx4 ) );
  mux2_1 U13267 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [18]), .ip2(n11586), .s(n11505), .op(\CORTEXM0DS_INST/u_logic/Vnjvx4 ) );
  mux2_1 U13268 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [19]), .ip2(n11587), .s(n11505), .op(\CORTEXM0DS_INST/u_logic/Ksjvx4 ) );
  mux2_1 U13269 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [20]), .ip2(n11588), .s(n11505), .op(\CORTEXM0DS_INST/u_logic/Zwjvx4 ) );
  mux2_1 U13270 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [21]), .ip2(n11589), .s(n11574), .op(\CORTEXM0DS_INST/u_logic/O1kvx4 ) );
  mux2_1 U13271 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [22]), .ip2(n11590), .s(n11505), .op(\CORTEXM0DS_INST/u_logic/D6kvx4 ) );
  mux2_1 U13272 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [3]), .ip2(n11591), .s(n11505), 
        .op(\CORTEXM0DS_INST/u_logic/Zakvx4 ) );
  mux2_1 U13273 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [4]), .ip2(n11592), .s(n11505), 
        .op(\CORTEXM0DS_INST/u_logic/Ofkvx4 ) );
  mux2_1 U13274 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [5]), .ip2(n11593), .s(n11574), 
        .op(\CORTEXM0DS_INST/u_logic/Dkkvx4 ) );
  mux2_1 U13275 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [6]), .ip2(n11594), .s(n11505), 
        .op(\CORTEXM0DS_INST/u_logic/Sokvx4 ) );
  mux2_1 U13276 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [24]), .ip2(n11595), .s(n11505), .op(\CORTEXM0DS_INST/u_logic/Htkvx4 ) );
  mux2_1 U13277 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [25]), .ip2(n11596), .s(n11574), .op(\CORTEXM0DS_INST/u_logic/Pxkvx4 ) );
  mux2_1 U13278 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [26]), .ip2(n11597), .s(n11505), .op(\CORTEXM0DS_INST/u_logic/E2lvx4 ) );
  mux2_1 U13279 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [27]), .ip2(n11598), .s(n11505), .op(\CORTEXM0DS_INST/u_logic/T6lvx4 ) );
  mux2_1 U13280 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [29]), .ip2(n11601), .s(n11505), .op(\CORTEXM0DS_INST/u_logic/Iblvx4 ) );
  mux2_1 U13281 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [30]), .ip2(n11602), .s(n11574), .op(\CORTEXM0DS_INST/u_logic/Eglvx4 ) );
  mux2_1 U13282 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [0]), .ip2(n11603), .s(n11505), 
        .op(\CORTEXM0DS_INST/u_logic/Ozlvx4 ) );
  mux2_1 U13283 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [1]), .ip2(n11604), .s(n11505), 
        .op(\CORTEXM0DS_INST/u_logic/Vzlvx4 ) );
  mux2_1 U13284 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [7]), .ip2(n11605), .s(n11574), 
        .op(\CORTEXM0DS_INST/u_logic/C0mvx4 ) );
  mux2_1 U13285 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [28]), .ip2(n11606), .s(n11574), .op(\CORTEXM0DS_INST/u_logic/J0mvx4 ) );
  mux2_1 U13286 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [31]), .ip2(n11617), .s(n11574), .op(\CORTEXM0DS_INST/u_logic/Q0mvx4 ) );
  nor2_1 U13287 ( .ip1(n11506), .ip2(n11576), .op(n11507) );
  mux2_1 U13288 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [9]), .ip2(n11577), .s(n11507), 
        .op(\CORTEXM0DS_INST/u_logic/Ciivx4 ) );
  mux2_1 U13289 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [2]), .ip2(n11578), .s(n11507), 
        .op(\CORTEXM0DS_INST/u_logic/Rmivx4 ) );
  mux2_1 U13290 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [10]), .ip2(n11579), .s(n11507), .op(\CORTEXM0DS_INST/u_logic/Grivx4 ) );
  mux2_1 U13291 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [11]), .ip2(n11580), .s(n11507), .op(\CORTEXM0DS_INST/u_logic/Vvivx4 ) );
  mux2_1 U13292 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [12]), .ip2(n11581), .s(n11507), .op(\CORTEXM0DS_INST/u_logic/K0jvx4 ) );
  mux2_1 U13293 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [13]), .ip2(n11582), .s(n11507), .op(\CORTEXM0DS_INST/u_logic/Z4jvx4 ) );
  mux2_1 U13294 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [14]), .ip2(n11583), .s(n11507), .op(\CORTEXM0DS_INST/u_logic/O9jvx4 ) );
  mux2_1 U13295 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [16]), .ip2(n11584), .s(n11507), .op(\CORTEXM0DS_INST/u_logic/Dejvx4 ) );
  mux2_1 U13296 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [17]), .ip2(n11585), .s(n11507), .op(\CORTEXM0DS_INST/u_logic/Sijvx4 ) );
  mux2_1 U13297 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [18]), .ip2(n11586), .s(n11507), .op(\CORTEXM0DS_INST/u_logic/Hnjvx4 ) );
  mux2_1 U13298 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [19]), .ip2(n11587), .s(n11507), .op(\CORTEXM0DS_INST/u_logic/Wrjvx4 ) );
  buf_1 U13299 ( .ip(n11507), .op(n11618) );
  mux2_1 U13300 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [20]), .ip2(n11588), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/Lwjvx4 ) );
  mux2_1 U13301 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [21]), .ip2(n11589), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/A1kvx4 ) );
  mux2_1 U13302 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [22]), .ip2(n11590), .s(n11507), .op(\CORTEXM0DS_INST/u_logic/P5kvx4 ) );
  mux2_1 U13303 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [3]), .ip2(n11591), .s(n11507), 
        .op(\CORTEXM0DS_INST/u_logic/Lakvx4 ) );
  mux2_1 U13304 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [4]), .ip2(n11592), .s(n11507), 
        .op(\CORTEXM0DS_INST/u_logic/Afkvx4 ) );
  mux2_1 U13305 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [5]), .ip2(n11593), .s(n11507), 
        .op(\CORTEXM0DS_INST/u_logic/Pjkvx4 ) );
  mux2_1 U13306 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [6]), .ip2(n11594), .s(n11507), 
        .op(\CORTEXM0DS_INST/u_logic/Eokvx4 ) );
  mux2_1 U13307 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [24]), .ip2(n11595), .s(n11507), .op(\CORTEXM0DS_INST/u_logic/Tskvx4 ) );
  mux2_1 U13308 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [25]), .ip2(n11596), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/Bxkvx4 ) );
  mux2_1 U13309 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [26]), .ip2(n11597), .s(n11507), .op(\CORTEXM0DS_INST/u_logic/Q1lvx4 ) );
  mux2_1 U13310 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [27]), .ip2(n11598), .s(n11507), .op(\CORTEXM0DS_INST/u_logic/F6lvx4 ) );
  mux2_1 U13311 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [29]), .ip2(n11601), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/Ualvx4 ) );
  mux2_1 U13312 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [30]), .ip2(n11602), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/Qflvx4 ) );
  mux2_1 U13313 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [0]), .ip2(n11603), .s(n11507), 
        .op(\CORTEXM0DS_INST/u_logic/Eenvx4 ) );
  mux2_1 U13314 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [1]), .ip2(n11604), .s(n11507), 
        .op(\CORTEXM0DS_INST/u_logic/Lenvx4 ) );
  mux2_1 U13315 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [7]), .ip2(n11605), .s(n11618), 
        .op(\CORTEXM0DS_INST/u_logic/Senvx4 ) );
  mux2_1 U13316 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [28]), .ip2(n11606), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/Zenvx4 ) );
  mux2_1 U13317 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [31]), .ip2(n11617), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/Gfnvx4 ) );
  nor2_1 U13318 ( .ip1(n11508), .ip2(n11576), .op(n11509) );
  mux2_1 U13319 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [9]), .ip2(n11577), .s(n11509), 
        .op(\CORTEXM0DS_INST/u_logic/Vhivx4 ) );
  buf_1 U13320 ( .ip(n11509), .op(n11621) );
  mux2_1 U13321 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [2]), .ip2(n11578), .s(n11621), 
        .op(\CORTEXM0DS_INST/u_logic/Kmivx4 ) );
  mux2_1 U13322 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [10]), .ip2(n11579), .s(n11509), .op(\CORTEXM0DS_INST/u_logic/Zqivx4 ) );
  mux2_1 U13323 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [11]), .ip2(n11580), .s(n11509), .op(\CORTEXM0DS_INST/u_logic/Ovivx4 ) );
  mux2_1 U13324 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [12]), .ip2(n11581), .s(n11509), .op(\CORTEXM0DS_INST/u_logic/D0jvx4 ) );
  mux2_1 U13325 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [13]), .ip2(n11582), .s(n11509), .op(\CORTEXM0DS_INST/u_logic/S4jvx4 ) );
  mux2_1 U13326 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [14]), .ip2(n11583), .s(n11509), .op(\CORTEXM0DS_INST/u_logic/H9jvx4 ) );
  mux2_1 U13327 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [16]), .ip2(n11584), .s(n11509), .op(\CORTEXM0DS_INST/u_logic/Wdjvx4 ) );
  mux2_1 U13328 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [17]), .ip2(n11585), .s(n11509), .op(\CORTEXM0DS_INST/u_logic/Lijvx4 ) );
  mux2_1 U13329 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [18]), .ip2(n11586), .s(n11509), .op(\CORTEXM0DS_INST/u_logic/Anjvx4 ) );
  mux2_1 U13330 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [19]), .ip2(n11587), .s(n11509), .op(\CORTEXM0DS_INST/u_logic/Prjvx4 ) );
  mux2_1 U13331 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [20]), .ip2(n11588), .s(n11509), .op(\CORTEXM0DS_INST/u_logic/Ewjvx4 ) );
  mux2_1 U13332 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [21]), .ip2(n11589), .s(n11621), .op(\CORTEXM0DS_INST/u_logic/T0kvx4 ) );
  mux2_1 U13333 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [22]), .ip2(n11590), .s(n11509), .op(\CORTEXM0DS_INST/u_logic/I5kvx4 ) );
  mux2_1 U13334 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [3]), .ip2(n11591), .s(n11509), 
        .op(\CORTEXM0DS_INST/u_logic/Eakvx4 ) );
  mux2_1 U13335 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [4]), .ip2(n11592), .s(n11509), 
        .op(\CORTEXM0DS_INST/u_logic/Tekvx4 ) );
  mux2_1 U13336 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [5]), .ip2(n11593), .s(n11621), 
        .op(\CORTEXM0DS_INST/u_logic/Ijkvx4 ) );
  mux2_1 U13337 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [6]), .ip2(n11594), .s(n11509), 
        .op(\CORTEXM0DS_INST/u_logic/Xnkvx4 ) );
  mux2_1 U13338 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [24]), .ip2(n11595), .s(n11509), .op(\CORTEXM0DS_INST/u_logic/Mskvx4 ) );
  mux2_1 U13339 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [25]), .ip2(n11596), .s(n11621), .op(\CORTEXM0DS_INST/u_logic/Uwkvx4 ) );
  mux2_1 U13340 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [26]), .ip2(n11597), .s(n11509), .op(\CORTEXM0DS_INST/u_logic/J1lvx4 ) );
  mux2_1 U13341 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [27]), .ip2(n11598), .s(n11509), .op(\CORTEXM0DS_INST/u_logic/Y5lvx4 ) );
  mux2_1 U13342 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [29]), .ip2(n11601), .s(n11509), .op(\CORTEXM0DS_INST/u_logic/Nalvx4 ) );
  mux2_1 U13343 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [30]), .ip2(n11602), .s(n11509), .op(\CORTEXM0DS_INST/u_logic/Jflvx4 ) );
  mux2_1 U13344 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [0]), .ip2(n11603), .s(n11509), 
        .op(\CORTEXM0DS_INST/u_logic/Bgnvx4 ) );
  mux2_1 U13345 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [7]), .ip2(n11605), .s(n11621), 
        .op(\CORTEXM0DS_INST/u_logic/Ignvx4 ) );
  mux2_1 U13346 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [31]), .ip2(n11617), .s(n11621), .op(\CORTEXM0DS_INST/u_logic/Wgnvx4 ) );
  mux2_1 U13347 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [28]), .ip2(n11606), .s(n11621), .op(\CORTEXM0DS_INST/u_logic/Dhnvx4 ) );
  mux2_1 U13348 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [1]), .ip2(n11604), .s(n11621), 
        .op(\CORTEXM0DS_INST/u_logic/Minvx4 ) );
  nand2_1 U13349 ( .ip1(n12117), .ip2(n11534), .op(n11524) );
  or2_1 U13350 ( .ip1(n11511), .ip2(n11510), .op(n11512) );
  nand2_1 U13351 ( .ip1(n11518), .ip2(n11512), .op(n11514) );
  or2_1 U13352 ( .ip1(n11513), .ip2(n11514), .op(n11517) );
  inv_1 U13353 ( .ip(n12114), .op(n11515) );
  or2_1 U13354 ( .ip1(n11515), .ip2(n11514), .op(n11516) );
  nand2_1 U13355 ( .ip1(n11517), .ip2(n11516), .op(n11520) );
  nor2_1 U13356 ( .ip1(n11518), .ip2(n11537), .op(n11519) );
  nor2_1 U13357 ( .ip1(n11520), .ip2(n11519), .op(n11521) );
  not_ab_or_c_or_d U13358 ( .ip1(n11549), .ip2(n12658), .ip3(n11548), .ip4(
        n11521), .op(n11523) );
  nand3_1 U13359 ( .ip1(n11524), .ip2(n11523), .ip3(n11522), .op(n11622) );
  nor2_1 U13360 ( .ip1(n11526), .ip2(n11525), .op(n11527) );
  mux2_1 U13361 ( .ip1(\CORTEXM0DS_INST/vis_psp [6]), .ip2(n11622), .s(n11527), 
        .op(\CORTEXM0DS_INST/u_logic/Hhivx4 ) );
  mux2_1 U13362 ( .ip1(\CORTEXM0DS_INST/vis_psp [7]), .ip2(n11577), .s(n11527), 
        .op(\CORTEXM0DS_INST/u_logic/Wlivx4 ) );
  mux2_1 U13363 ( .ip1(\CORTEXM0DS_INST/vis_psp [0]), .ip2(n11578), .s(n11527), 
        .op(\CORTEXM0DS_INST/u_logic/Lqivx4 ) );
  mux2_1 U13364 ( .ip1(\CORTEXM0DS_INST/vis_psp [8]), .ip2(n11579), .s(n11527), 
        .op(\CORTEXM0DS_INST/u_logic/Avivx4 ) );
  mux2_1 U13365 ( .ip1(\CORTEXM0DS_INST/vis_psp [9]), .ip2(n11580), .s(n11527), 
        .op(\CORTEXM0DS_INST/u_logic/Pzivx4 ) );
  mux2_1 U13366 ( .ip1(\CORTEXM0DS_INST/vis_psp [10]), .ip2(n11581), .s(n11527), .op(\CORTEXM0DS_INST/u_logic/E4jvx4 ) );
  mux2_1 U13367 ( .ip1(\CORTEXM0DS_INST/vis_psp [11]), .ip2(n11582), .s(n11527), .op(\CORTEXM0DS_INST/u_logic/T8jvx4 ) );
  mux2_1 U13368 ( .ip1(\CORTEXM0DS_INST/vis_psp [12]), .ip2(n11583), .s(n11527), .op(\CORTEXM0DS_INST/u_logic/Idjvx4 ) );
  mux2_1 U13369 ( .ip1(\CORTEXM0DS_INST/vis_psp [14]), .ip2(n11584), .s(n11527), .op(\CORTEXM0DS_INST/u_logic/Xhjvx4 ) );
  buf_1 U13370 ( .ip(n11527), .op(n11553) );
  mux2_1 U13371 ( .ip1(\CORTEXM0DS_INST/vis_psp [15]), .ip2(n11585), .s(n11553), .op(\CORTEXM0DS_INST/u_logic/Mmjvx4 ) );
  mux2_1 U13372 ( .ip1(\CORTEXM0DS_INST/vis_psp [16]), .ip2(n11586), .s(n11527), .op(\CORTEXM0DS_INST/u_logic/Brjvx4 ) );
  mux2_1 U13373 ( .ip1(\CORTEXM0DS_INST/vis_psp [17]), .ip2(n11587), .s(n11527), .op(\CORTEXM0DS_INST/u_logic/Qvjvx4 ) );
  mux2_1 U13374 ( .ip1(\CORTEXM0DS_INST/vis_psp [18]), .ip2(n11588), .s(n11553), .op(\CORTEXM0DS_INST/u_logic/F0kvx4 ) );
  mux2_1 U13375 ( .ip1(\CORTEXM0DS_INST/vis_psp [19]), .ip2(n11589), .s(n11527), .op(\CORTEXM0DS_INST/u_logic/U4kvx4 ) );
  mux2_1 U13376 ( .ip1(\CORTEXM0DS_INST/vis_psp [20]), .ip2(n11590), .s(n11527), .op(\CORTEXM0DS_INST/u_logic/J9kvx4 ) );
  mux2_1 U13377 ( .ip1(\CORTEXM0DS_INST/vis_psp [1]), .ip2(n11591), .s(n11527), 
        .op(\CORTEXM0DS_INST/u_logic/Fekvx4 ) );
  mux2_1 U13378 ( .ip1(\CORTEXM0DS_INST/vis_psp [2]), .ip2(n11592), .s(n11527), 
        .op(\CORTEXM0DS_INST/u_logic/Uikvx4 ) );
  mux2_1 U13379 ( .ip1(\CORTEXM0DS_INST/vis_psp [3]), .ip2(n11593), .s(n11527), 
        .op(\CORTEXM0DS_INST/u_logic/Jnkvx4 ) );
  mux2_1 U13380 ( .ip1(\CORTEXM0DS_INST/vis_psp [4]), .ip2(n11594), .s(n11527), 
        .op(\CORTEXM0DS_INST/u_logic/Yrkvx4 ) );
  mux2_1 U13381 ( .ip1(\CORTEXM0DS_INST/vis_psp [22]), .ip2(n11595), .s(n11527), .op(\CORTEXM0DS_INST/u_logic/Nwkvx4 ) );
  mux2_1 U13382 ( .ip1(\CORTEXM0DS_INST/vis_psp [23]), .ip2(n11596), .s(n11553), .op(\CORTEXM0DS_INST/u_logic/V0lvx4 ) );
  mux2_1 U13383 ( .ip1(\CORTEXM0DS_INST/vis_psp [24]), .ip2(n11597), .s(n11527), .op(\CORTEXM0DS_INST/u_logic/K5lvx4 ) );
  mux2_1 U13384 ( .ip1(\CORTEXM0DS_INST/vis_psp [25]), .ip2(n11598), .s(n11527), .op(\CORTEXM0DS_INST/u_logic/Z9lvx4 ) );
  mux2_1 U13385 ( .ip1(\CORTEXM0DS_INST/vis_psp [27]), .ip2(n11601), .s(n11553), .op(\CORTEXM0DS_INST/u_logic/Oelvx4 ) );
  mux2_1 U13386 ( .ip1(\CORTEXM0DS_INST/vis_psp [28]), .ip2(n11602), .s(n11553), .op(\CORTEXM0DS_INST/u_logic/Kjlvx4 ) );
  mux2_1 U13387 ( .ip1(\CORTEXM0DS_INST/vis_psp [29]), .ip2(n11617), .s(n11527), .op(\CORTEXM0DS_INST/u_logic/Mklvx4 ) );
  mux2_1 U13388 ( .ip1(\CORTEXM0DS_INST/vis_psp [26]), .ip2(n11606), .s(n11553), .op(\CORTEXM0DS_INST/u_logic/Tklvx4 ) );
  mux2_1 U13389 ( .ip1(\CORTEXM0DS_INST/vis_psp [5]), .ip2(n11605), .s(n11553), 
        .op(\CORTEXM0DS_INST/u_logic/Allvx4 ) );
  not_ab_or_c_or_d U13390 ( .ip1(n11549), .ip2(n12678), .ip3(n11529), .ip4(
        n11528), .op(n11533) );
  or2_1 U13391 ( .ip1(n12103), .ip2(n11530), .op(n11531) );
  nand3_1 U13392 ( .ip1(n11533), .ip2(n11532), .ip3(n11531), .op(n11619) );
  mux2_1 U13393 ( .ip1(\CORTEXM0DS_INST/vis_psp [21]), .ip2(n11619), .s(n11553), .op(\CORTEXM0DS_INST/u_logic/D8ivx4 ) );
  nand2_1 U13394 ( .ip1(n11535), .ip2(n11534), .op(n11552) );
  inv_1 U13395 ( .ip(n11540), .op(n11546) );
  nor2_1 U13396 ( .ip1(n11537), .ip2(n11536), .op(n11544) );
  or2_1 U13397 ( .ip1(n11538), .ip2(n11539), .op(n11542) );
  or2_1 U13398 ( .ip1(n11540), .ip2(n11539), .op(n11541) );
  nand2_1 U13399 ( .ip1(n11542), .ip2(n11541), .op(n11543) );
  not_ab_or_c_or_d U13400 ( .ip1(n11546), .ip2(n11545), .ip3(n11544), .ip4(
        n11543), .op(n11547) );
  not_ab_or_c_or_d U13401 ( .ip1(n11549), .ip2(n12665), .ip3(n11548), .ip4(
        n11547), .op(n11551) );
  nand3_1 U13402 ( .ip1(n11552), .ip2(n11551), .ip3(n11550), .op(n11620) );
  mux2_1 U13403 ( .ip1(\CORTEXM0DS_INST/vis_psp [13]), .ip2(n11620), .s(n11553), .op(\CORTEXM0DS_INST/u_logic/Scivx4 ) );
  mux2_1 U13404 ( .ip1(\CORTEXM0DS_INST/vis_msp [21]), .ip2(n11619), .s(n11554), .op(\CORTEXM0DS_INST/u_logic/W7ivx4 ) );
  mux2_1 U13405 ( .ip1(\CORTEXM0DS_INST/vis_msp [13]), .ip2(n11620), .s(n11554), .op(\CORTEXM0DS_INST/u_logic/Lcivx4 ) );
  mux2_1 U13406 ( .ip1(\CORTEXM0DS_INST/vis_msp [6]), .ip2(n11622), .s(n11554), 
        .op(\CORTEXM0DS_INST/u_logic/Ahivx4 ) );
  nor2_1 U13407 ( .ip1(n11556), .ip2(n11555), .op(n11562) );
  nand2_1 U13408 ( .ip1(n11557), .ip2(n11562), .op(n11558) );
  mux2_1 U13409 ( .ip1(n11619), .ip2(\CORTEXM0DS_INST/cm0_r14 [23]), .s(n11558), .op(\CORTEXM0DS_INST/u_logic/P7ivx4 ) );
  buf_1 U13410 ( .ip(n11558), .op(n11559) );
  mux2_1 U13411 ( .ip1(n11620), .ip2(\CORTEXM0DS_INST/cm0_r14 [15]), .s(n11559), .op(\CORTEXM0DS_INST/u_logic/Ecivx4 ) );
  mux2_1 U13412 ( .ip1(n11622), .ip2(\CORTEXM0DS_INST/cm0_r14 [8]), .s(n11558), 
        .op(\CORTEXM0DS_INST/u_logic/Tgivx4 ) );
  mux2_1 U13413 ( .ip1(n11577), .ip2(\CORTEXM0DS_INST/cm0_r14 [9]), .s(n11558), 
        .op(\CORTEXM0DS_INST/u_logic/Ilivx4 ) );
  mux2_1 U13414 ( .ip1(n11578), .ip2(\CORTEXM0DS_INST/cm0_r14 [2]), .s(n11558), 
        .op(\CORTEXM0DS_INST/u_logic/Xpivx4 ) );
  mux2_1 U13415 ( .ip1(n11579), .ip2(\CORTEXM0DS_INST/cm0_r14 [10]), .s(n11558), .op(\CORTEXM0DS_INST/u_logic/Muivx4 ) );
  mux2_1 U13416 ( .ip1(n11580), .ip2(\CORTEXM0DS_INST/cm0_r14 [11]), .s(n11558), .op(\CORTEXM0DS_INST/u_logic/Bzivx4 ) );
  mux2_1 U13417 ( .ip1(n11581), .ip2(\CORTEXM0DS_INST/cm0_r14 [12]), .s(n11558), .op(\CORTEXM0DS_INST/u_logic/Q3jvx4 ) );
  mux2_1 U13418 ( .ip1(n11582), .ip2(\CORTEXM0DS_INST/cm0_r14 [13]), .s(n11558), .op(\CORTEXM0DS_INST/u_logic/F8jvx4 ) );
  mux2_1 U13419 ( .ip1(n11583), .ip2(\CORTEXM0DS_INST/cm0_r14 [14]), .s(n11558), .op(\CORTEXM0DS_INST/u_logic/Ucjvx4 ) );
  mux2_1 U13420 ( .ip1(n11584), .ip2(\CORTEXM0DS_INST/cm0_r14 [16]), .s(n11558), .op(\CORTEXM0DS_INST/u_logic/Jhjvx4 ) );
  mux2_1 U13421 ( .ip1(n11585), .ip2(\CORTEXM0DS_INST/cm0_r14 [17]), .s(n11558), .op(\CORTEXM0DS_INST/u_logic/Yljvx4 ) );
  mux2_1 U13422 ( .ip1(n11586), .ip2(\CORTEXM0DS_INST/cm0_r14 [18]), .s(n11558), .op(\CORTEXM0DS_INST/u_logic/Nqjvx4 ) );
  mux2_1 U13423 ( .ip1(n11587), .ip2(\CORTEXM0DS_INST/cm0_r14 [19]), .s(n11558), .op(\CORTEXM0DS_INST/u_logic/Cvjvx4 ) );
  mux2_1 U13424 ( .ip1(n11588), .ip2(\CORTEXM0DS_INST/cm0_r14 [20]), .s(n11558), .op(\CORTEXM0DS_INST/u_logic/Rzjvx4 ) );
  mux2_1 U13425 ( .ip1(n11589), .ip2(\CORTEXM0DS_INST/cm0_r14 [21]), .s(n11558), .op(\CORTEXM0DS_INST/u_logic/G4kvx4 ) );
  mux2_1 U13426 ( .ip1(n11590), .ip2(\CORTEXM0DS_INST/cm0_r14 [22]), .s(n11558), .op(\CORTEXM0DS_INST/u_logic/V8kvx4 ) );
  mux2_1 U13427 ( .ip1(n11591), .ip2(\CORTEXM0DS_INST/cm0_r14 [3]), .s(n11559), 
        .op(\CORTEXM0DS_INST/u_logic/Rdkvx4 ) );
  mux2_1 U13428 ( .ip1(n11592), .ip2(\CORTEXM0DS_INST/cm0_r14 [4]), .s(n11558), 
        .op(\CORTEXM0DS_INST/u_logic/Gikvx4 ) );
  mux2_1 U13429 ( .ip1(n11593), .ip2(\CORTEXM0DS_INST/cm0_r14 [5]), .s(n11558), 
        .op(\CORTEXM0DS_INST/u_logic/Vmkvx4 ) );
  mux2_1 U13430 ( .ip1(n11594), .ip2(\CORTEXM0DS_INST/cm0_r14 [6]), .s(n11559), 
        .op(\CORTEXM0DS_INST/u_logic/Krkvx4 ) );
  mux2_1 U13431 ( .ip1(n11595), .ip2(\CORTEXM0DS_INST/cm0_r14 [24]), .s(n11558), .op(\CORTEXM0DS_INST/u_logic/Zvkvx4 ) );
  mux2_1 U13432 ( .ip1(n11596), .ip2(\CORTEXM0DS_INST/cm0_r14 [25]), .s(n11558), .op(\CORTEXM0DS_INST/u_logic/H0lvx4 ) );
  mux2_1 U13433 ( .ip1(n11597), .ip2(\CORTEXM0DS_INST/cm0_r14 [26]), .s(n11558), .op(\CORTEXM0DS_INST/u_logic/W4lvx4 ) );
  mux2_1 U13434 ( .ip1(n11598), .ip2(\CORTEXM0DS_INST/cm0_r14 [27]), .s(n11559), .op(\CORTEXM0DS_INST/u_logic/L9lvx4 ) );
  mux2_1 U13435 ( .ip1(n11601), .ip2(\CORTEXM0DS_INST/cm0_r14 [29]), .s(n11559), .op(\CORTEXM0DS_INST/u_logic/Aelvx4 ) );
  mux2_1 U13436 ( .ip1(n11602), .ip2(\CORTEXM0DS_INST/cm0_r14 [30]), .s(n11559), .op(\CORTEXM0DS_INST/u_logic/Wilvx4 ) );
  mux2_1 U13437 ( .ip1(n11603), .ip2(\CORTEXM0DS_INST/cm0_r14 [0]), .s(n11559), 
        .op(\CORTEXM0DS_INST/u_logic/Vslvx4 ) );
  mux2_1 U13438 ( .ip1(n11604), .ip2(\CORTEXM0DS_INST/cm0_r14 [1]), .s(n11559), 
        .op(\CORTEXM0DS_INST/u_logic/Ctlvx4 ) );
  mux2_1 U13439 ( .ip1(n11605), .ip2(\CORTEXM0DS_INST/cm0_r14 [7]), .s(n11559), 
        .op(\CORTEXM0DS_INST/u_logic/Jtlvx4 ) );
  mux2_1 U13440 ( .ip1(n11606), .ip2(\CORTEXM0DS_INST/cm0_r14 [28]), .s(n11559), .op(\CORTEXM0DS_INST/u_logic/Qtlvx4 ) );
  mux2_1 U13441 ( .ip1(n11617), .ip2(\CORTEXM0DS_INST/cm0_r14 [31]), .s(n11559), .op(\CORTEXM0DS_INST/u_logic/Xtlvx4 ) );
  mux2_1 U13442 ( .ip1(n11619), .ip2(\CORTEXM0DS_INST/cm0_r12 [23]), .s(n11560), .op(\CORTEXM0DS_INST/u_logic/I7ivx4 ) );
  mux2_1 U13443 ( .ip1(n11620), .ip2(\CORTEXM0DS_INST/cm0_r12 [15]), .s(n11560), .op(\CORTEXM0DS_INST/u_logic/Xbivx4 ) );
  mux2_1 U13444 ( .ip1(n11622), .ip2(\CORTEXM0DS_INST/cm0_r12 [8]), .s(n11560), 
        .op(\CORTEXM0DS_INST/u_logic/Mgivx4 ) );
  mux2_1 U13445 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [23]), .ip2(n11619), .s(n11561), .op(\CORTEXM0DS_INST/u_logic/B7ivx4 ) );
  mux2_1 U13446 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [15]), .ip2(n11620), .s(n11561), .op(\CORTEXM0DS_INST/u_logic/Qbivx4 ) );
  mux2_1 U13447 ( .ip1(\CORTEXM0DS_INST/cm0_r07 [8]), .ip2(n11622), .s(n11561), 
        .op(\CORTEXM0DS_INST/u_logic/Fgivx4 ) );
  inv_1 U13448 ( .ip(n11562), .op(n11575) );
  nor2_1 U13449 ( .ip1(n11563), .ip2(n11575), .op(n11564) );
  buf_1 U13450 ( .ip(n11564), .op(n11565) );
  mux2_1 U13451 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [23]), .ip2(n11619), .s(n11565), .op(\CORTEXM0DS_INST/u_logic/U6ivx4 ) );
  mux2_1 U13452 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [15]), .ip2(n11620), .s(n11564), .op(\CORTEXM0DS_INST/u_logic/Jbivx4 ) );
  mux2_1 U13453 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [8]), .ip2(n11622), .s(n11564), 
        .op(\CORTEXM0DS_INST/u_logic/Yfivx4 ) );
  mux2_1 U13454 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [9]), .ip2(n11577), .s(n11565), 
        .op(\CORTEXM0DS_INST/u_logic/Nkivx4 ) );
  mux2_1 U13455 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [2]), .ip2(n11578), .s(n11565), 
        .op(\CORTEXM0DS_INST/u_logic/Cpivx4 ) );
  mux2_1 U13456 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [10]), .ip2(n11579), .s(n11564), .op(\CORTEXM0DS_INST/u_logic/Rtivx4 ) );
  mux2_1 U13457 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [11]), .ip2(n11580), .s(n11564), .op(\CORTEXM0DS_INST/u_logic/Gyivx4 ) );
  mux2_1 U13458 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [12]), .ip2(n11581), .s(n11564), .op(\CORTEXM0DS_INST/u_logic/V2jvx4 ) );
  mux2_1 U13459 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [13]), .ip2(n11582), .s(n11564), .op(\CORTEXM0DS_INST/u_logic/K7jvx4 ) );
  mux2_1 U13460 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [14]), .ip2(n11583), .s(n11564), .op(\CORTEXM0DS_INST/u_logic/Zbjvx4 ) );
  mux2_1 U13461 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [16]), .ip2(n11584), .s(n11564), .op(\CORTEXM0DS_INST/u_logic/Ogjvx4 ) );
  mux2_1 U13462 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [17]), .ip2(n11585), .s(n11564), .op(\CORTEXM0DS_INST/u_logic/Dljvx4 ) );
  mux2_1 U13463 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [18]), .ip2(n11586), .s(n11564), .op(\CORTEXM0DS_INST/u_logic/Spjvx4 ) );
  mux2_1 U13464 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [19]), .ip2(n11587), .s(n11564), .op(\CORTEXM0DS_INST/u_logic/Hujvx4 ) );
  mux2_1 U13465 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [20]), .ip2(n11588), .s(n11564), .op(\CORTEXM0DS_INST/u_logic/Wyjvx4 ) );
  mux2_1 U13466 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [21]), .ip2(n11589), .s(n11564), .op(\CORTEXM0DS_INST/u_logic/L3kvx4 ) );
  mux2_1 U13467 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [22]), .ip2(n11590), .s(n11564), .op(\CORTEXM0DS_INST/u_logic/A8kvx4 ) );
  mux2_1 U13468 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [3]), .ip2(n11591), .s(n11564), 
        .op(\CORTEXM0DS_INST/u_logic/Wckvx4 ) );
  mux2_1 U13469 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [4]), .ip2(n11592), .s(n11564), 
        .op(\CORTEXM0DS_INST/u_logic/Lhkvx4 ) );
  mux2_1 U13470 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [5]), .ip2(n11593), .s(n11564), 
        .op(\CORTEXM0DS_INST/u_logic/Amkvx4 ) );
  mux2_1 U13471 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [6]), .ip2(n11594), .s(n11565), 
        .op(\CORTEXM0DS_INST/u_logic/Pqkvx4 ) );
  mux2_1 U13472 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [24]), .ip2(n11595), .s(n11564), .op(\CORTEXM0DS_INST/u_logic/Evkvx4 ) );
  mux2_1 U13473 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [25]), .ip2(n11596), .s(n11565), .op(\CORTEXM0DS_INST/u_logic/Mzkvx4 ) );
  mux2_1 U13474 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [26]), .ip2(n11597), .s(n11564), .op(\CORTEXM0DS_INST/u_logic/B4lvx4 ) );
  mux2_1 U13475 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [27]), .ip2(n11598), .s(n11564), .op(\CORTEXM0DS_INST/u_logic/Q8lvx4 ) );
  mux2_1 U13476 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [29]), .ip2(n11601), .s(n11564), .op(\CORTEXM0DS_INST/u_logic/Fdlvx4 ) );
  mux2_1 U13477 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [30]), .ip2(n11602), .s(n11565), .op(\CORTEXM0DS_INST/u_logic/Bilvx4 ) );
  mux2_1 U13478 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [0]), .ip2(n11603), .s(n11565), 
        .op(\CORTEXM0DS_INST/u_logic/Uolvx4 ) );
  mux2_1 U13479 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [1]), .ip2(n11604), .s(n11565), 
        .op(\CORTEXM0DS_INST/u_logic/Bplvx4 ) );
  mux2_1 U13480 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [7]), .ip2(n11605), .s(n11565), 
        .op(\CORTEXM0DS_INST/u_logic/Iplvx4 ) );
  mux2_1 U13481 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [28]), .ip2(n11606), .s(n11565), .op(\CORTEXM0DS_INST/u_logic/Pplvx4 ) );
  mux2_1 U13482 ( .ip1(\CORTEXM0DS_INST/cm0_r06 [31]), .ip2(n11617), .s(n11565), .op(\CORTEXM0DS_INST/u_logic/Wplvx4 ) );
  mux2_1 U13483 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [23]), .ip2(n11619), .s(n11566), .op(\CORTEXM0DS_INST/u_logic/N6ivx4 ) );
  mux2_1 U13484 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [15]), .ip2(n11620), .s(n11566), .op(\CORTEXM0DS_INST/u_logic/Cbivx4 ) );
  mux2_1 U13485 ( .ip1(\CORTEXM0DS_INST/cm0_r05 [8]), .ip2(n11622), .s(n11566), 
        .op(\CORTEXM0DS_INST/u_logic/Rfivx4 ) );
  mux2_1 U13486 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [23]), .ip2(n11619), .s(n11567), .op(\CORTEXM0DS_INST/u_logic/G6ivx4 ) );
  mux2_1 U13487 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [15]), .ip2(n11620), .s(n11567), .op(\CORTEXM0DS_INST/u_logic/Vaivx4 ) );
  mux2_1 U13488 ( .ip1(\CORTEXM0DS_INST/cm0_r04 [8]), .ip2(n11622), .s(n11567), 
        .op(\CORTEXM0DS_INST/u_logic/Kfivx4 ) );
  mux2_1 U13489 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [23]), .ip2(n11619), .s(n11568), .op(\CORTEXM0DS_INST/u_logic/Z5ivx4 ) );
  mux2_1 U13490 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [15]), .ip2(n11620), .s(n11568), .op(\CORTEXM0DS_INST/u_logic/Oaivx4 ) );
  mux2_1 U13491 ( .ip1(\CORTEXM0DS_INST/cm0_r11 [8]), .ip2(n11622), .s(n11568), 
        .op(\CORTEXM0DS_INST/u_logic/Dfivx4 ) );
  nor2_1 U13492 ( .ip1(n11569), .ip2(n11575), .op(n11570) );
  buf_1 U13493 ( .ip(n11570), .op(n11571) );
  mux2_1 U13494 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [23]), .ip2(n11619), .s(n11571), .op(\CORTEXM0DS_INST/u_logic/S5ivx4 ) );
  mux2_1 U13495 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [15]), .ip2(n11620), .s(n11570), .op(\CORTEXM0DS_INST/u_logic/Haivx4 ) );
  mux2_1 U13496 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [8]), .ip2(n11622), .s(n11570), 
        .op(\CORTEXM0DS_INST/u_logic/Weivx4 ) );
  mux2_1 U13497 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [9]), .ip2(n11577), .s(n11570), 
        .op(\CORTEXM0DS_INST/u_logic/Ljivx4 ) );
  mux2_1 U13498 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [2]), .ip2(n11578), .s(n11570), 
        .op(\CORTEXM0DS_INST/u_logic/Aoivx4 ) );
  mux2_1 U13499 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [10]), .ip2(n11579), .s(n11570), .op(\CORTEXM0DS_INST/u_logic/Psivx4 ) );
  mux2_1 U13500 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [11]), .ip2(n11580), .s(n11570), .op(\CORTEXM0DS_INST/u_logic/Exivx4 ) );
  mux2_1 U13501 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [12]), .ip2(n11581), .s(n11570), .op(\CORTEXM0DS_INST/u_logic/T1jvx4 ) );
  mux2_1 U13502 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [13]), .ip2(n11582), .s(n11570), .op(\CORTEXM0DS_INST/u_logic/I6jvx4 ) );
  mux2_1 U13503 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [14]), .ip2(n11583), .s(n11570), .op(\CORTEXM0DS_INST/u_logic/Xajvx4 ) );
  mux2_1 U13504 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [16]), .ip2(n11584), .s(n11570), .op(\CORTEXM0DS_INST/u_logic/Mfjvx4 ) );
  mux2_1 U13505 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [17]), .ip2(n11585), .s(n11570), .op(\CORTEXM0DS_INST/u_logic/Bkjvx4 ) );
  mux2_1 U13506 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [18]), .ip2(n11586), .s(n11570), .op(\CORTEXM0DS_INST/u_logic/Qojvx4 ) );
  mux2_1 U13507 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [19]), .ip2(n11587), .s(n11570), .op(\CORTEXM0DS_INST/u_logic/Ftjvx4 ) );
  mux2_1 U13508 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [20]), .ip2(n11588), .s(n11570), .op(\CORTEXM0DS_INST/u_logic/Uxjvx4 ) );
  mux2_1 U13509 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [21]), .ip2(n11589), .s(n11570), .op(\CORTEXM0DS_INST/u_logic/J2kvx4 ) );
  mux2_1 U13510 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [22]), .ip2(n11590), .s(n11571), .op(\CORTEXM0DS_INST/u_logic/Y6kvx4 ) );
  mux2_1 U13511 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [3]), .ip2(n11591), .s(n11571), 
        .op(\CORTEXM0DS_INST/u_logic/Ubkvx4 ) );
  mux2_1 U13512 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [4]), .ip2(n11592), .s(n11571), 
        .op(\CORTEXM0DS_INST/u_logic/Jgkvx4 ) );
  mux2_1 U13513 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [5]), .ip2(n11593), .s(n11570), 
        .op(\CORTEXM0DS_INST/u_logic/Ykkvx4 ) );
  mux2_1 U13514 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [6]), .ip2(n11594), .s(n11570), 
        .op(\CORTEXM0DS_INST/u_logic/Npkvx4 ) );
  mux2_1 U13515 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [24]), .ip2(n11595), .s(n11571), .op(\CORTEXM0DS_INST/u_logic/Cukvx4 ) );
  mux2_1 U13516 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [25]), .ip2(n11596), .s(n11570), .op(\CORTEXM0DS_INST/u_logic/Kykvx4 ) );
  mux2_1 U13517 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [26]), .ip2(n11597), .s(n11570), .op(\CORTEXM0DS_INST/u_logic/Z2lvx4 ) );
  mux2_1 U13518 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [27]), .ip2(n11598), .s(n11570), .op(\CORTEXM0DS_INST/u_logic/O7lvx4 ) );
  mux2_1 U13519 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [29]), .ip2(n11601), .s(n11570), .op(\CORTEXM0DS_INST/u_logic/Dclvx4 ) );
  mux2_1 U13520 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [30]), .ip2(n11602), .s(n11571), .op(\CORTEXM0DS_INST/u_logic/Zglvx4 ) );
  mux2_1 U13521 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [0]), .ip2(n11603), .s(n11571), 
        .op(\CORTEXM0DS_INST/u_logic/Nvlvx4 ) );
  mux2_1 U13522 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [1]), .ip2(n11604), .s(n11571), 
        .op(\CORTEXM0DS_INST/u_logic/Uvlvx4 ) );
  mux2_1 U13523 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [7]), .ip2(n11605), .s(n11571), 
        .op(\CORTEXM0DS_INST/u_logic/Bwlvx4 ) );
  mux2_1 U13524 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [28]), .ip2(n11606), .s(n11571), .op(\CORTEXM0DS_INST/u_logic/Iwlvx4 ) );
  mux2_1 U13525 ( .ip1(\CORTEXM0DS_INST/cm0_r10 [31]), .ip2(n11617), .s(n11571), .op(\CORTEXM0DS_INST/u_logic/Pwlvx4 ) );
  mux2_1 U13526 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [23]), .ip2(n11619), .s(n11572), .op(\CORTEXM0DS_INST/u_logic/L5ivx4 ) );
  mux2_1 U13527 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [15]), .ip2(n11620), .s(n11572), .op(\CORTEXM0DS_INST/u_logic/Aaivx4 ) );
  mux2_1 U13528 ( .ip1(\CORTEXM0DS_INST/cm0_r09 [8]), .ip2(n11622), .s(n11572), 
        .op(\CORTEXM0DS_INST/u_logic/Peivx4 ) );
  mux2_1 U13529 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [23]), .ip2(n11619), .s(n11573), .op(\CORTEXM0DS_INST/u_logic/E5ivx4 ) );
  mux2_1 U13530 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [15]), .ip2(n11620), .s(n11573), .op(\CORTEXM0DS_INST/u_logic/T9ivx4 ) );
  mux2_1 U13531 ( .ip1(\CORTEXM0DS_INST/cm0_r08 [8]), .ip2(n11622), .s(n11573), 
        .op(\CORTEXM0DS_INST/u_logic/Ieivx4 ) );
  mux2_1 U13532 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [23]), .ip2(n11619), .s(n11574), .op(\CORTEXM0DS_INST/u_logic/X4ivx4 ) );
  mux2_1 U13533 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [15]), .ip2(n11620), .s(n11574), .op(\CORTEXM0DS_INST/u_logic/M9ivx4 ) );
  mux2_1 U13534 ( .ip1(\CORTEXM0DS_INST/cm0_r03 [8]), .ip2(n11622), .s(n11574), 
        .op(\CORTEXM0DS_INST/u_logic/Beivx4 ) );
  nor2_1 U13535 ( .ip1(n11576), .ip2(n11575), .op(n11600) );
  buf_1 U13536 ( .ip(n11600), .op(n11616) );
  mux2_1 U13537 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [23]), .ip2(n11619), .s(n11616), .op(\CORTEXM0DS_INST/u_logic/Q4ivx4 ) );
  mux2_1 U13538 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [15]), .ip2(n11620), .s(n11600), .op(\CORTEXM0DS_INST/u_logic/F9ivx4 ) );
  mux2_1 U13539 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [8]), .ip2(n11622), .s(n11600), 
        .op(\CORTEXM0DS_INST/u_logic/Udivx4 ) );
  mux2_1 U13540 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [9]), .ip2(n11577), .s(n11616), 
        .op(\CORTEXM0DS_INST/u_logic/Jiivx4 ) );
  mux2_1 U13541 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [2]), .ip2(n11578), .s(n11616), 
        .op(\CORTEXM0DS_INST/u_logic/Ymivx4 ) );
  mux2_1 U13542 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [10]), .ip2(n11579), .s(n11600), .op(\CORTEXM0DS_INST/u_logic/Nrivx4 ) );
  mux2_1 U13543 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [11]), .ip2(n11580), .s(n11600), .op(\CORTEXM0DS_INST/u_logic/Cwivx4 ) );
  mux2_1 U13544 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [12]), .ip2(n11581), .s(n11600), .op(\CORTEXM0DS_INST/u_logic/R0jvx4 ) );
  mux2_1 U13545 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [13]), .ip2(n11582), .s(n11600), .op(\CORTEXM0DS_INST/u_logic/G5jvx4 ) );
  mux2_1 U13546 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [14]), .ip2(n11583), .s(n11600), .op(\CORTEXM0DS_INST/u_logic/V9jvx4 ) );
  mux2_1 U13547 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [16]), .ip2(n11584), .s(n11600), .op(\CORTEXM0DS_INST/u_logic/Kejvx4 ) );
  mux2_1 U13548 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [17]), .ip2(n11585), .s(n11600), .op(\CORTEXM0DS_INST/u_logic/Zijvx4 ) );
  mux2_1 U13549 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [18]), .ip2(n11586), .s(n11600), .op(\CORTEXM0DS_INST/u_logic/Onjvx4 ) );
  mux2_1 U13550 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [19]), .ip2(n11587), .s(n11600), .op(\CORTEXM0DS_INST/u_logic/Dsjvx4 ) );
  mux2_1 U13551 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [20]), .ip2(n11588), .s(n11600), .op(\CORTEXM0DS_INST/u_logic/Swjvx4 ) );
  mux2_1 U13552 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [21]), .ip2(n11589), .s(n11600), .op(\CORTEXM0DS_INST/u_logic/H1kvx4 ) );
  mux2_1 U13553 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [22]), .ip2(n11590), .s(n11600), .op(\CORTEXM0DS_INST/u_logic/W5kvx4 ) );
  mux2_1 U13554 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [3]), .ip2(n11591), .s(n11600), 
        .op(\CORTEXM0DS_INST/u_logic/Sakvx4 ) );
  mux2_1 U13555 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [4]), .ip2(n11592), .s(n11600), 
        .op(\CORTEXM0DS_INST/u_logic/Hfkvx4 ) );
  mux2_1 U13556 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [5]), .ip2(n11593), .s(n11600), 
        .op(\CORTEXM0DS_INST/u_logic/Wjkvx4 ) );
  mux2_1 U13557 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [6]), .ip2(n11594), .s(n11616), 
        .op(\CORTEXM0DS_INST/u_logic/Lokvx4 ) );
  mux2_1 U13558 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [24]), .ip2(n11595), .s(n11600), .op(\CORTEXM0DS_INST/u_logic/Atkvx4 ) );
  mux2_1 U13559 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [25]), .ip2(n11596), .s(n11616), .op(\CORTEXM0DS_INST/u_logic/Ixkvx4 ) );
  mux2_1 U13560 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [26]), .ip2(n11597), .s(n11600), .op(\CORTEXM0DS_INST/u_logic/X1lvx4 ) );
  mux2_1 U13561 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [27]), .ip2(n11598), .s(n11600), .op(\CORTEXM0DS_INST/u_logic/M6lvx4 ) );
  nor2_1 U13562 ( .ip1(n11599), .ip2(n11614), .op(n4180) );
  mux2_1 U13563 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [29]), .ip2(n11601), .s(n11600), .op(\CORTEXM0DS_INST/u_logic/Bblvx4 ) );
  mux2_1 U13564 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [30]), .ip2(n11602), .s(n11616), .op(\CORTEXM0DS_INST/u_logic/Xflvx4 ) );
  mux2_1 U13565 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [0]), .ip2(n11603), .s(n11616), 
        .op(\CORTEXM0DS_INST/u_logic/X0mvx4 ) );
  mux2_1 U13566 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [1]), .ip2(n11604), .s(n11616), 
        .op(\CORTEXM0DS_INST/u_logic/E1mvx4 ) );
  mux2_1 U13567 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [7]), .ip2(n11605), .s(n11616), 
        .op(\CORTEXM0DS_INST/u_logic/L1mvx4 ) );
  mux2_1 U13568 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [28]), .ip2(n11606), .s(n11616), .op(\CORTEXM0DS_INST/u_logic/S1mvx4 ) );
  nand2_1 U13569 ( .ip1(n11608), .ip2(n11607), .op(n11613) );
  nand2_1 U13570 ( .ip1(n11609), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [20]), 
        .op(n11612) );
  nand2_1 U13571 ( .ip1(n11610), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [20]), 
        .op(n11611) );
  nand3_1 U13572 ( .ip1(n11613), .ip2(n11612), .ip3(n11611), .op(n4109) );
  nor2_1 U13573 ( .ip1(n11615), .ip2(n11614), .op(n4110) );
  mux2_1 U13574 ( .ip1(\CORTEXM0DS_INST/cm0_r02 [31]), .ip2(n11617), .s(n11616), .op(\CORTEXM0DS_INST/u_logic/Z1mvx4 ) );
  mux2_1 U13575 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [23]), .ip2(n11619), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/J4ivx4 ) );
  mux2_1 U13576 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [15]), .ip2(n11620), .s(n11618), .op(\CORTEXM0DS_INST/u_logic/Y8ivx4 ) );
  mux2_1 U13577 ( .ip1(\CORTEXM0DS_INST/cm0_r01 [8]), .ip2(n11622), .s(n11618), 
        .op(\CORTEXM0DS_INST/u_logic/Ndivx4 ) );
  mux2_1 U13578 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [23]), .ip2(n11619), .s(n11621), .op(\CORTEXM0DS_INST/u_logic/C4ivx4 ) );
  mux2_1 U13579 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [15]), .ip2(n11620), .s(n11621), .op(\CORTEXM0DS_INST/u_logic/R8ivx4 ) );
  mux2_1 U13580 ( .ip1(\CORTEXM0DS_INST/cm0_r00 [8]), .ip2(n11622), .s(n11621), 
        .op(\CORTEXM0DS_INST/u_logic/Gdivx4 ) );
  nor2_1 U13581 ( .ip1(n11623), .ip2(n11811), .op(n3978) );
  nor2_1 U13582 ( .ip1(n11624), .ip2(n11776), .op(n11627) );
  nor2_1 U13583 ( .ip1(n11625), .ip2(n11778), .op(n11626) );
  ab_or_c_or_d U13584 ( .ip1(n11783), .ip2(n11628), .ip3(n11627), .ip4(n11626), 
        .op(n11630) );
  not_ab_or_c_or_d U13585 ( .ip1(n11629), .ip2(n11783), .ip3(1'b0), .ip4(n5938), .op(n11638) );
  mux2_1 U13586 ( .ip1(\CORTEXM0DS_INST/vis_apsr [3]), .ip2(n11630), .s(n11638), .op(\CORTEXM0DS_INST/u_logic/V3ivx4 ) );
  nor2_1 U13587 ( .ip1(n11631), .ip2(n11778), .op(n11637) );
  nor2_1 U13588 ( .ip1(n11632), .ip2(n11776), .op(n11636) );
  nor2_1 U13589 ( .ip1(n11634), .ip2(n11633), .op(n11635) );
  nor4_1 U13590 ( .ip1(n5938), .ip2(n11637), .ip3(n11636), .ip4(n11635), .op(
        n11640) );
  nor2_1 U13591 ( .ip1(\CORTEXM0DS_INST/vis_apsr [2]), .ip2(n11638), .op(
        n11639) );
  nor2_1 U13592 ( .ip1(n11640), .ip2(n11639), .op(
        \CORTEXM0DS_INST/u_logic/Cflvx4 ) );
  inv_1 U13593 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [1]), .op(n11648) );
  inv_1 U13594 ( .ip(n3224), .op(n11641) );
  nor3_1 U13595 ( .ip1(\CORTEXM0DS_INST/u_logic/Qsgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Sx3wx4 ), .ip3(n11641), .op(n11647) );
  nand2_1 U13596 ( .ip1(\CORTEXM0DS_INST/u_logic/R1ivx4 ), .ip2(n11642), .op(
        n11645) );
  nand2_1 U13597 ( .ip1(\CORTEXM0DS_INST/u_logic/K1ivx4 ), .ip2(n11643), .op(
        n11644) );
  nand2_1 U13598 ( .ip1(n11645), .ip2(n11644), .op(n11646) );
  not_ab_or_c_or_d U13599 ( .ip1(\CORTEXM0DS_INST/u_logic/M2ivx4 ), .ip2(
        n11648), .ip3(n11647), .ip4(n11646), .op(n11708) );
  nor2_1 U13600 ( .ip1(\CORTEXM0DS_INST/u_logic/Efgvx4 ), .ip2(n12613), .op(
        n11649) );
  nand4_1 U13601 ( .ip1(n11651), .ip2(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip3(
        n11650), .ip4(n11649), .op(n11657) );
  nand2_1 U13602 ( .ip1(n12405), .ip2(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .op(
        n11656) );
  inv_1 U13603 ( .ip(n11652), .op(n11653) );
  nand3_1 U13604 ( .ip1(n11654), .ip2(n11653), .ip3(n12075), .op(n11655) );
  nand4_1 U13605 ( .ip1(n11658), .ip2(n11657), .ip3(n11656), .ip4(n11655), 
        .op(n11665) );
  nand3_1 U13606 ( .ip1(n11661), .ip2(n11660), .ip3(n11659), .op(n11701) );
  nor2_1 U13607 ( .ip1(n11662), .ip2(n11701), .op(n11664) );
  nor2_1 U13608 ( .ip1(n3217), .ip2(n12646), .op(n12404) );
  nor4_1 U13609 ( .ip1(\CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip2(n12404), .ip3(
        n12686), .ip4(n12096), .op(n11663) );
  not_ab_or_c_or_d U13610 ( .ip1(n12647), .ip2(n11665), .ip3(n11664), .ip4(
        n11663), .op(n11850) );
  nor2_1 U13611 ( .ip1(\CORTEXM0DS_INST/u_logic/Krgvx4 ), .ip2(n11850), .op(
        n11696) );
  inv_1 U13612 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [14]), .op(n11687) );
  nor2_1 U13613 ( .ip1(n3233), .ip2(n11666), .op(n11686) );
  inv_1 U13614 ( .ip(\CORTEXM0DS_INST/u_logic/T2ivx4 ), .op(n11667) );
  nor2_1 U13615 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [0]), .ip2(n11667), 
        .op(n11676) );
  nand2_1 U13616 ( .ip1(\CORTEXM0DS_INST/u_logic/Nzhvx4 ), .ip2(n11668), .op(
        n11674) );
  inv_1 U13617 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [3]), .op(n11669) );
  nand2_1 U13618 ( .ip1(\CORTEXM0DS_INST/u_logic/Y1ivx4 ), .ip2(n11669), .op(
        n11673) );
  inv_1 U13619 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [15]), .op(n11842) );
  nand2_1 U13620 ( .ip1(\CORTEXM0DS_INST/u_logic/Syhvx4 ), .ip2(n11842), .op(
        n11672) );
  inv_1 U13621 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [8]), .op(n11670) );
  nand2_1 U13622 ( .ip1(\CORTEXM0DS_INST/u_logic/P0ivx4 ), .ip2(n11670), .op(
        n11671) );
  nand4_1 U13623 ( .ip1(n11674), .ip2(n11673), .ip3(n11672), .ip4(n11671), 
        .op(n11675) );
  not_ab_or_c_or_d U13624 ( .ip1(\CORTEXM0DS_INST/u_logic/B0ivx4 ), .ip2(
        n11677), .ip3(n11676), .ip4(n11675), .op(n11684) );
  inv_1 U13625 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [9]), .op(n11678) );
  nand2_1 U13626 ( .ip1(\CORTEXM0DS_INST/u_logic/I0ivx4 ), .ip2(n11678), .op(
        n11683) );
  inv_1 U13627 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [13]), .op(n11679) );
  nand2_1 U13628 ( .ip1(\CORTEXM0DS_INST/u_logic/Gzhvx4 ), .ip2(n11679), .op(
        n11682) );
  inv_1 U13629 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [6]), .op(n11680) );
  nand2_1 U13630 ( .ip1(\CORTEXM0DS_INST/u_logic/D1ivx4 ), .ip2(n11680), .op(
        n11681) );
  nand4_1 U13631 ( .ip1(n11684), .ip2(n11683), .ip3(n11682), .ip4(n11681), 
        .op(n11685) );
  not_ab_or_c_or_d U13632 ( .ip1(\CORTEXM0DS_INST/u_logic/Zyhvx4 ), .ip2(
        n11687), .ip3(n11686), .ip4(n11685), .op(n11694) );
  inv_1 U13633 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [11]), .op(n11688) );
  nand2_1 U13634 ( .ip1(\CORTEXM0DS_INST/u_logic/Uzhvx4 ), .ip2(n11688), .op(
        n11693) );
  inv_1 U13635 ( .ip(\CORTEXM0DS_INST/u_logic/Eqgvx4 ), .op(n11826) );
  nand2_1 U13636 ( .ip1(\CORTEXM0DS_INST/u_logic/Owgvx4 ), .ip2(n11826), .op(
        n11692) );
  nor2_1 U13637 ( .ip1(n2326), .ip2(n3224), .op(n11689) );
  nor2_1 U13638 ( .ip1(n12750), .ip2(n11689), .op(n12010) );
  nand2_1 U13639 ( .ip1(n12010), .ip2(n11690), .op(n11691) );
  nand4_1 U13640 ( .ip1(n11694), .ip2(n11693), .ip3(n11692), .ip4(n11691), 
        .op(n11695) );
  not_ab_or_c_or_d U13641 ( .ip1(\CORTEXM0DS_INST/u_logic/W0ivx4 ), .ip2(n3223), .ip3(n11696), .ip4(n11695), .op(n11707) );
  nand3_1 U13642 ( .ip1(n11698), .ip2(n11697), .ip3(n6210), .op(n11699) );
  or2_1 U13643 ( .ip1(n11699), .ip2(n11700), .op(n11703) );
  or2_1 U13644 ( .ip1(n11701), .ip2(n11700), .op(n11702) );
  nand2_1 U13645 ( .ip1(n11703), .ip2(n11702), .op(n11856) );
  nand2_1 U13646 ( .ip1(n11856), .ip2(n11852), .op(n11706) );
  inv_1 U13647 ( .ip(\CORTEXM0DS_INST/u_logic/T1i2z4 [2]), .op(n11704) );
  nand2_1 U13648 ( .ip1(\CORTEXM0DS_INST/u_logic/F2ivx4 ), .ip2(n11704), .op(
        n11705) );
  nand4_1 U13649 ( .ip1(n11708), .ip2(n11707), .ip3(n11706), .ip4(n11705), 
        .op(n11709) );
  nand2_1 U13650 ( .ip1(\CORTEXM0DS_INST/u_logic/Vogvx4 ), .ip2(n11709), .op(
        n11712) );
  not_ab_or_c_or_d U13651 ( .ip1(n11710), .ip2(n10865), .ip3(TXEV_top_out), 
        .ip4(n12687), .op(n11711) );
  nand2_1 U13652 ( .ip1(n11712), .ip2(n11711), .op(n11717) );
  nand4_1 U13653 ( .ip1(n11715), .ip2(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip3(
        n11714), .ip4(n11713), .op(n11716) );
  mux2_1 U13654 ( .ip1(n11717), .ip2(n11716), .s(
        \CORTEXM0DS_INST/u_logic/Ih8vx4 ), .op(
        \CORTEXM0DS_INST/u_logic/H3ivx4 ) );
  inv_1 U13655 ( .ip(n3217), .op(n12396) );
  mux2_1 U13656 ( .ip1(n11719), .ip2(n11718), .s(n12396), .op(n11724) );
  inv_1 U13657 ( .ip(n11720), .op(n11721) );
  not_ab_or_c_or_d U13658 ( .ip1(n11722), .ip2(n11721), .ip3(
        \CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip4(n5938), .op(n11723) );
  mux2_1 U13659 ( .ip1(\CORTEXM0DS_INST/u_logic/Oy8vx4 ), .ip2(n11724), .s(
        n11723), .op(\CORTEXM0DS_INST/u_logic/Sqivx4 ) );
  nand3_1 U13660 ( .ip1(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), .ip2(n11725), .ip3(
        n11730), .op(n11742) );
  or2_1 U13661 ( .ip1(n11726), .ip2(\CORTEXM0DS_INST/cm0_control[1] ), .op(
        n11728) );
  or2_1 U13662 ( .ip1(\CORTEXM0DS_INST/vis_pc [1]), .ip2(
        \CORTEXM0DS_INST/cm0_control[1] ), .op(n11727) );
  nand2_1 U13663 ( .ip1(n11728), .ip2(n11727), .op(n11738) );
  nor2_1 U13664 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n11729), .op(
        n11735) );
  or2_1 U13665 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n11730), .op(
        n11732) );
  or2_1 U13666 ( .ip1(\CORTEXM0DS_INST/u_logic/Uz8vx4 ), .ip2(n11730), .op(
        n11731) );
  nand2_1 U13667 ( .ip1(n11732), .ip2(n11731), .op(n11734) );
  nor2_1 U13668 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6gvx4 ), .ip2(n12550), .op(
        n11739) );
  nor2_1 U13669 ( .ip1(n12334), .ip2(n11739), .op(n11733) );
  nor4_1 U13670 ( .ip1(n11736), .ip2(n11735), .ip3(n11734), .ip4(n11733), .op(
        n11737) );
  or2_1 U13671 ( .ip1(n11738), .ip2(n11737), .op(n11741) );
  nand4_1 U13672 ( .ip1(\CORTEXM0DS_INST/u_logic/B19vx4 ), .ip2(n12034), .ip3(
        n11739), .ip4(n12535), .op(n11740) );
  nand3_1 U13673 ( .ip1(n11742), .ip2(n11741), .ip3(n11740), .op(n11765) );
  nand2_1 U13674 ( .ip1(n11744), .ip2(n11743), .op(n11749) );
  nand2_1 U13675 ( .ip1(n11746), .ip2(n11745), .op(n11747) );
  nand3_1 U13676 ( .ip1(n11749), .ip2(n11748), .ip3(n11747), .op(n11761) );
  nor2_1 U13677 ( .ip1(n11751), .ip2(n11750), .op(n11753) );
  not_ab_or_c_or_d U13678 ( .ip1(n11755), .ip2(n11754), .ip3(n11753), .ip4(
        n11752), .op(n11759) );
  nand2_1 U13679 ( .ip1(\CORTEXM0DS_INST/u_logic/P39vx4 ), .ip2(n11756), .op(
        n11757) );
  nand3_1 U13680 ( .ip1(n11759), .ip2(n11758), .ip3(n11757), .op(n11760) );
  not_ab_or_c_or_d U13681 ( .ip1(n11762), .ip2(n6210), .ip3(n11761), .ip4(
        n11760), .op(n11763) );
  nor2_1 U13682 ( .ip1(n5938), .ip2(n11763), .op(n11764) );
  mux2_1 U13683 ( .ip1(\CORTEXM0DS_INST/u_logic/O7evx4 ), .ip2(n11765), .s(
        n11764), .op(\CORTEXM0DS_INST/u_logic/Hllvx4 ) );
  nand2_1 U13684 ( .ip1(\CORTEXM0DS_INST/vis_pc [1]), .ip2(
        \CORTEXM0DS_INST/u_logic/Hx8vx4 ), .op(n11767) );
  nand2_1 U13685 ( .ip1(n11768), .ip2(n12669), .op(n11766) );
  nand2_1 U13686 ( .ip1(n11767), .ip2(n11766), .op(n11774) );
  nand4_1 U13687 ( .ip1(\CORTEXM0DS_INST/u_logic/Qm9vx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Yo9vx4 ), .ip3(n11769), .ip4(n11768), .op(
        n11770) );
  nand3_1 U13688 ( .ip1(n11771), .ip2(n11770), .ip3(n11862), .op(n11772) );
  nand2_1 U13689 ( .ip1(n11772), .ip2(n12642), .op(n11773) );
  mux2_1 U13690 ( .ip1(n11774), .ip2(\CORTEXM0DS_INST/cm0_control[1] ), .s(
        n11773), .op(\CORTEXM0DS_INST/u_logic/Ollvx4 ) );
  nor3_1 U13691 ( .ip1(n12685), .ip2(n11775), .ip3(n12635), .op(n3128) );
  nor2_1 U13692 ( .ip1(n11777), .ip2(n11776), .op(n11781) );
  nor2_1 U13693 ( .ip1(n11779), .ip2(n11778), .op(n11780) );
  ab_or_c_or_d U13694 ( .ip1(n11783), .ip2(n11782), .ip3(n11781), .ip4(n11780), 
        .op(n11786) );
  not_ab_or_c_or_d U13695 ( .ip1(n11784), .ip2(n11783), .ip3(1'b0), .ip4(n5938), .op(n11785) );
  mux2_1 U13696 ( .ip1(\CORTEXM0DS_INST/vis_apsr [1]), .ip2(n11786), .s(n11785), .op(\CORTEXM0DS_INST/u_logic/Finvx4 ) );
  inv_1 U13697 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [5]), .op(n11905) );
  nor2_1 U13698 ( .ip1(n11810), .ip2(n11905), .op(n3081) );
  and2_1 U13699 ( .ip1(\CORTEXM0DS_INST/u_logic/L0i2z4 [5]), .ip2(n11787), 
        .op(n3082) );
  nand2_1 U13700 ( .ip1(n11788), .ip2(n11821), .op(n11809) );
  nor2_1 U13701 ( .ip1(n11790), .ip2(n11789), .op(n11791) );
  or2_1 U13702 ( .ip1(\CORTEXM0DS_INST/u_logic/Zuh2z4 [9]), .ip2(n11791), .op(
        n11793) );
  or2_1 U13703 ( .ip1(n11833), .ip2(n11791), .op(n11792) );
  nand2_1 U13704 ( .ip1(n11793), .ip2(n11792), .op(n11805) );
  nor2_1 U13705 ( .ip1(n11795), .ip2(n11794), .op(n11798) );
  nor2_1 U13706 ( .ip1(n11814), .ip2(n11796), .op(n11797) );
  not_ab_or_c_or_d U13707 ( .ip1(n11799), .ip2(
        \CORTEXM0DS_INST/u_logic/Czh2z4 [7]), .ip3(n11798), .ip4(n11797), .op(
        n11804) );
  nand2_1 U13708 ( .ip1(n11800), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [7]), 
        .op(n11803) );
  nand2_1 U13709 ( .ip1(\CORTEXM0DS_INST/u_logic/T1i2z4 [7]), .ip2(n11801), 
        .op(n11802) );
  nand4_1 U13710 ( .ip1(n11805), .ip2(n11804), .ip3(n11803), .ip4(n11802), 
        .op(n11806) );
  nand2_1 U13711 ( .ip1(n11807), .ip2(n11806), .op(n11808) );
  nand2_1 U13712 ( .ip1(n11809), .ip2(n11808), .op(n3048) );
  inv_1 U13713 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [7]), .op(n11916) );
  nor2_1 U13714 ( .ip1(n11810), .ip2(n11916), .op(n3049) );
  nor2_1 U13715 ( .ip1(n11812), .ip2(n11811), .op(n3024) );
  nor2_1 U13716 ( .ip1(n11814), .ip2(n11813), .op(n11819) );
  nand2_1 U13717 ( .ip1(n11827), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [21]), 
        .op(n11817) );
  nand2_1 U13718 ( .ip1(n11833), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [13]), 
        .op(n11816) );
  nand2_1 U13719 ( .ip1(n11823), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [29]), 
        .op(n11815) );
  nand3_1 U13720 ( .ip1(n11817), .ip2(n11816), .ip3(n11815), .op(n11818) );
  not_ab_or_c_or_d U13721 ( .ip1(n12637), .ip2(
        \CORTEXM0DS_INST/u_logic/Psh2z4 [1]), .ip3(n11819), .ip4(n11818), .op(
        n11820) );
  nor2_1 U13722 ( .ip1(n11820), .ip2(n11839), .op(n3025) );
  and2_1 U13723 ( .ip1(n11822), .ip2(n11821), .op(n3015) );
  nand2_1 U13724 ( .ip1(n11823), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [31]), 
        .op(n11836) );
  and2_1 U13725 ( .ip1(n11824), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [7]), 
        .op(n11832) );
  nor2_1 U13726 ( .ip1(n11826), .ip2(n11825), .op(n11831) );
  and2_1 U13727 ( .ip1(n11827), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [23]), 
        .op(n11830) );
  nor2_1 U13728 ( .ip1(n11828), .ip2(n12636), .op(n11829) );
  nor4_1 U13729 ( .ip1(n11832), .ip2(n11831), .ip3(n11830), .ip4(n11829), .op(
        n11835) );
  nand2_1 U13730 ( .ip1(n11833), .ip2(\CORTEXM0DS_INST/u_logic/Zuh2z4 [15]), 
        .op(n11834) );
  nand3_1 U13731 ( .ip1(n11836), .ip2(n11835), .ip3(n11834), .op(n11837) );
  not_ab_or_c_or_d U13732 ( .ip1(\CORTEXM0DS_INST/u_logic/Txh2z4 [1]), .ip2(
        n12637), .ip3(n11838), .ip4(n11837), .op(n11840) );
  nor2_1 U13733 ( .ip1(n11840), .ip2(n11839), .op(n3016) );
  nor2_1 U13734 ( .ip1(n11842), .ip2(n11841), .op(n2984) );
  nor2_1 U13735 ( .ip1(n11843), .ip2(n11862), .op(n2791) );
  mux2_1 U13736 ( .ip1(n11865), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [0]), .s(
        n2786), .op(n6192) );
  mux2_1 U13737 ( .ip1(n11865), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [1]), .s(
        n2774), .op(n6189) );
  mux2_1 U13738 ( .ip1(n11865), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [14]), 
        .s(n2757), .op(n6183) );
  nor2_1 U13739 ( .ip1(n11844), .ip2(n11862), .op(n2714) );
  mux2_1 U13740 ( .ip1(n11865), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [6]), .s(
        n2711), .op(n6182) );
  mux2_1 U13741 ( .ip1(n11865), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [5]), .s(
        n2686), .op(n6180) );
  nor2_1 U13742 ( .ip1(n11845), .ip2(n11862), .op(n2648) );
  mux2_1 U13743 ( .ip1(n11865), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [12]), 
        .s(n2645), .op(n6177) );
  mux2_1 U13744 ( .ip1(n11865), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [4]), .s(
        n2644), .op(n6175) );
  nor3_1 U13745 ( .ip1(n11847), .ip2(n11846), .ip3(n11862), .op(n2627) );
  mux2_1 U13746 ( .ip1(n11865), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [3]), .s(
        n2624), .op(n6173) );
  mux2_1 U13747 ( .ip1(n11865), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [2]), .s(
        n2623), .op(n6171) );
  mux2_1 U13748 ( .ip1(n11865), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [7]), .s(
        n2577), .op(n6166) );
  nand2_1 U13749 ( .ip1(n12687), .ip2(n12395), .op(n11848) );
  nand2_1 U13750 ( .ip1(\CORTEXM0DS_INST/u_logic/Krgvx4 ), .ip2(n11848), .op(
        n11849) );
  nand2_1 U13751 ( .ip1(n11850), .ip2(n11849), .op(n6164) );
  or2_1 U13752 ( .ip1(n11851), .ip2(n11852), .op(n11854) );
  or2_1 U13753 ( .ip1(n12687), .ip2(n11852), .op(n11853) );
  nand2_1 U13754 ( .ip1(n11854), .ip2(n11853), .op(n11855) );
  or2_1 U13755 ( .ip1(n11856), .ip2(n11855), .op(n6163) );
  nor2_1 U13756 ( .ip1(n11857), .ip2(n11862), .op(n2544) );
  mux2_1 U13757 ( .ip1(n11865), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [10]), 
        .s(n2541), .op(n6162) );
  mux2_1 U13758 ( .ip1(n11865), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [11]), 
        .s(n2533), .op(n6159) );
  mux2_1 U13759 ( .ip1(n11865), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [9]), .s(
        n2514), .op(n6157) );
  mux2_1 U13760 ( .ip1(n11865), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [8]), .s(
        n2513), .op(n6156) );
  nor2_1 U13761 ( .ip1(n11858), .ip2(n11862), .op(n2512) );
  mux2_1 U13762 ( .ip1(n11865), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [13]), 
        .s(n2500), .op(n6153) );
  nand2_1 U13763 ( .ip1(n11859), .ip2(n12687), .op(n11860) );
  nand3_1 U13764 ( .ip1(n11860), .ip2(n2490), .ip3(
        \CORTEXM0DS_INST/u_logic/Qsgvx4 ), .op(n11861) );
  nand2_1 U13765 ( .ip1(n2492), .ip2(n11861), .op(n6149) );
  nor3_1 U13766 ( .ip1(n11864), .ip2(n11863), .ip3(n11862), .op(n2464) );
  mux2_1 U13767 ( .ip1(n11865), .ip2(\CORTEXM0DS_INST/u_logic/L0i2z4 [15]), 
        .s(n2460), .op(n6147) );
  nand2_1 U13768 ( .ip1(n11866), .ip2(\CORTEXM0DS_INST/u_logic/Mf8vx4 ), .op(
        n11875) );
  nand3_1 U13769 ( .ip1(n11867), .ip2(n12683), .ip3(n12635), .op(n11868) );
  nand3_1 U13770 ( .ip1(n11875), .ip2(\CORTEXM0DS_INST/u_logic/Izgvx4 ), .ip3(
        n11868), .op(n11870) );
  nand3_1 U13771 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [0]), .ip2(
        \CORTEXM0DS_INST/u_logic/F2hvx4 ), .ip3(n11871), .op(n11869) );
  nand2_1 U13772 ( .ip1(n11870), .ip2(n11869), .op(n6145) );
  nand2_1 U13773 ( .ip1(n11875), .ip2(\CORTEXM0DS_INST/u_logic/F2hvx4 ), .op(
        n11872) );
  nand2_1 U13774 ( .ip1(n11871), .ip2(n11879), .op(n11873) );
  nor2_1 U13775 ( .ip1(n11872), .ip2(n11873), .op(n12003) );
  inv_1 U13776 ( .ip(n11872), .op(n11874) );
  nand2_1 U13777 ( .ip1(n11874), .ip2(n11873), .op(n11950) );
  nor2_1 U13778 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [0]), .ip2(n11950), 
        .op(n11877) );
  inv_1 U13779 ( .ip(n11875), .op(n11878) );
  nor3_1 U13780 ( .ip1(\CORTEXM0DS_INST/u_logic/F2hvx4 ), .ip2(n11878), .ip3(
        n11879), .op(n11876) );
  ab_or_c_or_d U13781 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [0]), .ip2(n12003), .ip3(n11877), .ip4(n11876), .op(n6144) );
  or2_1 U13782 ( .ip1(\CORTEXM0DS_INST/u_logic/F2hvx4 ), .ip2(n11878), .op(
        n11881) );
  or2_1 U13783 ( .ip1(n11879), .ip2(n11878), .op(n11880) );
  nand2_1 U13784 ( .ip1(n11881), .ip2(n11880), .op(n11891) );
  nor3_1 U13785 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [0]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [1]), .ip3(n11950), .op(n11883) );
  and2_1 U13786 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [1]), .ip2(n12003), 
        .op(n11882) );
  ab_or_c_or_d U13787 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [1]), .ip2(n11891), .ip3(n11883), .ip4(n11882), .op(n6143) );
  nand2_1 U13788 ( .ip1(n12003), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [2]), 
        .op(n11888) );
  inv_1 U13789 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [2]), .op(n11885) );
  nand2_1 U13790 ( .ip1(n11883), .ip2(n11885), .op(n11889) );
  or2_1 U13791 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [1]), .ip2(n11891), .op(
        n11884) );
  inv_1 U13792 ( .ip(n11950), .op(n12004) );
  or2_1 U13793 ( .ip1(n12004), .ip2(n11891), .op(n11998) );
  nand2_1 U13794 ( .ip1(n11884), .ip2(n11998), .op(n11886) );
  or2_1 U13795 ( .ip1(n11886), .ip2(n11885), .op(n11887) );
  nand3_1 U13796 ( .ip1(n11888), .ip2(n11889), .ip3(n11887), .op(n6142) );
  nor2_1 U13797 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [3]), .ip2(n11889), 
        .op(n11897) );
  inv_1 U13798 ( .ip(n11890), .op(n11892) );
  or2_1 U13799 ( .ip1(n11892), .ip2(n11891), .op(n11893) );
  nand2_1 U13800 ( .ip1(n11998), .ip2(n11893), .op(n11899) );
  nor2_1 U13801 ( .ip1(n11899), .ip2(n11894), .op(n11895) );
  ab_or_c_or_d U13802 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [3]), .ip2(n12003), .ip3(n11897), .ip4(n11895), .op(n6141) );
  nand2_1 U13803 ( .ip1(n12003), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [4]), 
        .op(n11901) );
  nand2_1 U13804 ( .ip1(n11897), .ip2(n11896), .op(n11902) );
  nand2_1 U13805 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [3]), .ip2(n12004), 
        .op(n11898) );
  nand2_1 U13806 ( .ip1(n11899), .ip2(n11898), .op(n11903) );
  nand2_1 U13807 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [4]), .ip2(n11903), 
        .op(n11900) );
  nand3_1 U13808 ( .ip1(n11901), .ip2(n11902), .ip3(n11900), .op(n6140) );
  nor2_1 U13809 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [5]), .ip2(n11902), 
        .op(n11910) );
  or2_1 U13810 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [4]), .ip2(n11903), .op(
        n11904) );
  nand2_1 U13811 ( .ip1(n11904), .ip2(n11998), .op(n11908) );
  nor2_1 U13812 ( .ip1(n11908), .ip2(n11905), .op(n11906) );
  ab_or_c_or_d U13813 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [5]), .ip2(n12003), .ip3(n11910), .ip4(n11906), .op(n6139) );
  nand2_1 U13814 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [5]), .ip2(n12004), 
        .op(n11907) );
  nand2_1 U13815 ( .ip1(n11908), .ip2(n11907), .op(n11914) );
  nand2_1 U13816 ( .ip1(n11914), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [6]), 
        .op(n11912) );
  nand2_1 U13817 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [6]), .ip2(n12003), 
        .op(n11911) );
  inv_1 U13818 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [6]), .op(n11909) );
  nand2_1 U13819 ( .ip1(n11910), .ip2(n11909), .op(n11913) );
  nand3_1 U13820 ( .ip1(n11912), .ip2(n11911), .ip3(n11913), .op(n6138) );
  nor2_1 U13821 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [7]), .ip2(n11913), 
        .op(n11931) );
  or2_1 U13822 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [6]), .ip2(n11914), .op(
        n11915) );
  nand2_1 U13823 ( .ip1(n11915), .ip2(n11998), .op(n11953) );
  nor2_1 U13824 ( .ip1(n11953), .ip2(n11916), .op(n11917) );
  ab_or_c_or_d U13825 ( .ip1(n12003), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [7]), .ip3(n11931), .ip4(n11917), .op(n6137) );
  nand2_1 U13826 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [7]), .ip2(n12004), 
        .op(n11918) );
  nand2_1 U13827 ( .ip1(n11953), .ip2(n11918), .op(n11944) );
  nand2_1 U13828 ( .ip1(n11944), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [8]), 
        .op(n11921) );
  nand2_1 U13829 ( .ip1(n12003), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [8]), 
        .op(n11920) );
  or2_1 U13830 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [8]), .ip2(n11944), .op(
        n11919) );
  nand2_1 U13831 ( .ip1(n11919), .ip2(n11998), .op(n11933) );
  nand2_1 U13832 ( .ip1(n12004), .ip2(n11933), .op(n11924) );
  nand3_1 U13833 ( .ip1(n11921), .ip2(n11920), .ip3(n11924), .op(n6136) );
  mux2_1 U13834 ( .ip1(n11924), .ip2(n11933), .s(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [9]), .op(n11923) );
  nand2_1 U13835 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [9]), .ip2(n12003), 
        .op(n11922) );
  nand2_1 U13836 ( .ip1(n11923), .ip2(n11922), .op(n6135) );
  nor3_1 U13837 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [9]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [10]), .ip3(n11924), .op(n11930) );
  inv_1 U13838 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [10]), .op(n11925) );
  or2_1 U13839 ( .ip1(n11933), .ip2(n11925), .op(n11928) );
  nand2_1 U13840 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [9]), .ip2(n12004), 
        .op(n11926) );
  or2_1 U13841 ( .ip1(n11926), .ip2(n11925), .op(n11927) );
  nand2_1 U13842 ( .ip1(n11928), .ip2(n11927), .op(n11929) );
  ab_or_c_or_d U13843 ( .ip1(n12003), .ip2(
        \CORTEXM0DS_INST/u_logic/Czh2z4 [10]), .ip3(n11930), .ip4(n11929), 
        .op(n6134) );
  nand2_1 U13844 ( .ip1(n12003), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [11]), 
        .op(n11937) );
  nand2_1 U13845 ( .ip1(n11939), .ip2(n11931), .op(n11938) );
  or2_1 U13846 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [9]), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [10]), .op(n11932) );
  nand2_1 U13847 ( .ip1(n11932), .ip2(n12004), .op(n11934) );
  nand2_1 U13848 ( .ip1(n11934), .ip2(n11933), .op(n11935) );
  nand2_1 U13849 ( .ip1(n11935), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [11]), 
        .op(n11936) );
  nand3_1 U13850 ( .ip1(n11937), .ip2(n11938), .ip3(n11936), .op(n6133) );
  nor2_1 U13851 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [12]), .ip2(n11938), 
        .op(n11943) );
  nor2_1 U13852 ( .ip1(n11950), .ip2(n11939), .op(n11951) );
  nor2_1 U13853 ( .ip1(n11951), .ip2(n11944), .op(n11941) );
  inv_1 U13854 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [12]), .op(n11940) );
  nor2_1 U13855 ( .ip1(n11941), .ip2(n11940), .op(n11942) );
  ab_or_c_or_d U13856 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [12]), .ip2(
        n12003), .ip3(n11943), .ip4(n11942), .op(n6132) );
  nand2_1 U13857 ( .ip1(n12003), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [13]), 
        .op(n11948) );
  inv_1 U13858 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [13]), .op(n11945) );
  nand2_1 U13859 ( .ip1(n11943), .ip2(n11945), .op(n11955) );
  not_ab_or_c_or_d U13860 ( .ip1(n12004), .ip2(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [12]), .ip3(n11951), .ip4(n11944), 
        .op(n11946) );
  or2_1 U13861 ( .ip1(n11946), .ip2(n11945), .op(n11947) );
  nand3_1 U13862 ( .ip1(n11948), .ip2(n11955), .ip3(n11947), .op(n6131) );
  or2_1 U13863 ( .ip1(n11950), .ip2(n11949), .op(n11954) );
  inv_1 U13864 ( .ip(n11951), .op(n11952) );
  nand3_1 U13865 ( .ip1(n11954), .ip2(n11953), .ip3(n11952), .op(n11958) );
  nor2_1 U13866 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [14]), .ip2(n11955), 
        .op(n11957) );
  and2_1 U13867 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [14]), .ip2(n12003), 
        .op(n11956) );
  ab_or_c_or_d U13868 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [14]), .ip2(
        n11958), .ip3(n11957), .ip4(n11956), .op(n6130) );
  nand2_1 U13869 ( .ip1(n12003), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [15]), 
        .op(n11962) );
  inv_1 U13870 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [15]), .op(n11960) );
  nand2_1 U13871 ( .ip1(n11957), .ip2(n11960), .op(n11965) );
  or2_1 U13872 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [14]), .ip2(n11958), 
        .op(n11959) );
  nand2_1 U13873 ( .ip1(n11959), .ip2(n11998), .op(n11964) );
  or2_1 U13874 ( .ip1(n11964), .ip2(n11960), .op(n11961) );
  nand3_1 U13875 ( .ip1(n11962), .ip2(n11965), .ip3(n11961), .op(n6129) );
  nand2_1 U13876 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [15]), .ip2(n12004), 
        .op(n11963) );
  nand2_1 U13877 ( .ip1(n11964), .ip2(n11963), .op(n11975) );
  nor2_1 U13878 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [16]), .ip2(n11965), 
        .op(n11967) );
  and2_1 U13879 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [16]), .ip2(n12003), 
        .op(n11966) );
  ab_or_c_or_d U13880 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [16]), .ip2(
        n11975), .ip3(n11967), .ip4(n11966), .op(n6128) );
  nand2_1 U13881 ( .ip1(n12003), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [17]), 
        .op(n11972) );
  inv_1 U13882 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [17]), .op(n11969) );
  nand2_1 U13883 ( .ip1(n11967), .ip2(n11969), .op(n11973) );
  or2_1 U13884 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [16]), .ip2(n11975), 
        .op(n11968) );
  nand2_1 U13885 ( .ip1(n11968), .ip2(n11998), .op(n11970) );
  or2_1 U13886 ( .ip1(n11970), .ip2(n11969), .op(n11971) );
  nand3_1 U13887 ( .ip1(n11972), .ip2(n11973), .ip3(n11971), .op(n6127) );
  nor2_1 U13888 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [18]), .ip2(n11973), 
        .op(n11981) );
  inv_1 U13889 ( .ip(n11974), .op(n11976) );
  or2_1 U13890 ( .ip1(n11976), .ip2(n11975), .op(n11977) );
  nand2_1 U13891 ( .ip1(n11998), .ip2(n11977), .op(n11983) );
  inv_1 U13892 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [18]), .op(n11978) );
  nor2_1 U13893 ( .ip1(n11983), .ip2(n11978), .op(n11979) );
  ab_or_c_or_d U13894 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [18]), .ip2(
        n12003), .ip3(n11981), .ip4(n11979), .op(n6126) );
  nand2_1 U13895 ( .ip1(n12003), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [19]), 
        .op(n11985) );
  inv_1 U13896 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [19]), .op(n11980) );
  nand2_1 U13897 ( .ip1(n11981), .ip2(n11980), .op(n11986) );
  nand2_1 U13898 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [18]), .ip2(n12004), 
        .op(n11982) );
  nand2_1 U13899 ( .ip1(n11983), .ip2(n11982), .op(n11987) );
  nand2_1 U13900 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [19]), .ip2(n11987), 
        .op(n11984) );
  nand3_1 U13901 ( .ip1(n11985), .ip2(n11986), .ip3(n11984), .op(n6125) );
  nor2_1 U13902 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [20]), .ip2(n11986), 
        .op(n11992) );
  or2_1 U13903 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [19]), .ip2(n11987), 
        .op(n11988) );
  nand2_1 U13904 ( .ip1(n11988), .ip2(n11998), .op(n11994) );
  inv_1 U13905 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [20]), .op(n11989) );
  nor2_1 U13906 ( .ip1(n11994), .ip2(n11989), .op(n11990) );
  ab_or_c_or_d U13907 ( .ip1(n12003), .ip2(
        \CORTEXM0DS_INST/u_logic/Czh2z4 [20]), .ip3(n11992), .ip4(n11990), 
        .op(n6124) );
  nand2_1 U13908 ( .ip1(n12003), .ip2(\CORTEXM0DS_INST/u_logic/Czh2z4 [21]), 
        .op(n11996) );
  inv_1 U13909 ( .ip(\CORTEXM0DS_INST/u_logic/Irh2z4 [21]), .op(n11991) );
  nand2_1 U13910 ( .ip1(n11992), .ip2(n11991), .op(n12000) );
  nand2_1 U13911 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [20]), .ip2(n12004), 
        .op(n11993) );
  nand2_1 U13912 ( .ip1(n11994), .ip2(n11993), .op(n11997) );
  nand2_1 U13913 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [21]), .ip2(n11997), 
        .op(n11995) );
  nand3_1 U13914 ( .ip1(n11996), .ip2(n12000), .ip3(n11995), .op(n6123) );
  or2_1 U13915 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [21]), .ip2(n11997), 
        .op(n11999) );
  nand2_1 U13916 ( .ip1(n11999), .ip2(n11998), .op(n12006) );
  mux2_1 U13917 ( .ip1(n12000), .ip2(n12006), .s(
        \CORTEXM0DS_INST/u_logic/Irh2z4 [22]), .op(n12002) );
  nand2_1 U13918 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [22]), .ip2(n12003), 
        .op(n12001) );
  nand2_1 U13919 ( .ip1(n12002), .ip2(n12001), .op(n6122) );
  nand2_1 U13920 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [23]), .ip2(n12003), 
        .op(n12009) );
  nand2_1 U13921 ( .ip1(n12004), .ip2(\CORTEXM0DS_INST/u_logic/Irh2z4 [22]), 
        .op(n12005) );
  nand2_1 U13922 ( .ip1(n12006), .ip2(n12005), .op(n12007) );
  nand2_1 U13923 ( .ip1(\CORTEXM0DS_INST/u_logic/Irh2z4 [23]), .ip2(n12007), 
        .op(n12008) );
  nand2_1 U13924 ( .ip1(n12009), .ip2(n12008), .op(n6121) );
  inv_1 U13925 ( .ip(n12010), .op(n12014) );
  nand2_1 U13926 ( .ip1(n12011), .ip2(n12687), .op(n12012) );
  nand3_1 U13927 ( .ip1(n12012), .ip2(n2328), .ip3(
        \CORTEXM0DS_INST/u_logic/R3hvx4 ), .op(n12013) );
  nand2_1 U13928 ( .ip1(n12014), .ip2(n12013), .op(n6119) );
  nor3_1 U13929 ( .ip1(n3231), .ip2(n2270), .ip3(n2271), .op(n12015) );
  nand4_1 U13930 ( .ip1(\CORTEXM0DS_INST/u_logic/Sx3wx4 ), .ip2(n2267), .ip3(
        n12015), .ip4(\CORTEXM0DS_INST/u_logic/O24wx4 ), .op(n12016) );
  nor2_1 U13931 ( .ip1(n12017), .ip2(n12016), .op(n12018) );
  or2_1 U13932 ( .ip1(SYSRESETREQ_top_out), .ip2(n12018), .op(n6118) );
  nand3_1 U13933 ( .ip1(n2217), .ip2(n2216), .ip3(n2215), .op(n6117) );
  inv_1 U13934 ( .ip(n2213), .op(n2214) );
  or2_1 U13935 ( .ip1(\CORTEXM0DS_INST/u_logic/V2qvx4 ), .ip2(n2209), .op(
        n12021) );
  inv_1 U13936 ( .ip(n2208), .op(n12019) );
  or2_1 U13937 ( .ip1(n12019), .ip2(n2209), .op(n12020) );
  nand2_1 U13938 ( .ip1(n12021), .ip2(n12020), .op(n12022) );
  or2_1 U13939 ( .ip1(n2212), .ip2(n12022), .op(n6116) );
  nor2_1 U13940 ( .ip1(n12472), .ip2(n2205), .op(n12023) );
  nor2_1 U13941 ( .ip1(n12024), .ip2(n12023), .op(n6115) );
  and2_1 U13942 ( .ip1(n12025), .ip2(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .op(
        n12029) );
  not_ab_or_c_or_d U13943 ( .ip1(n3217), .ip2(n12027), .ip3(n5938), .ip4(
        n12026), .op(n12028) );
  or2_1 U13944 ( .ip1(n12029), .ip2(n12028), .op(n6114) );
  nand3_1 U13945 ( .ip1(n12642), .ip2(n2197), .ip3(n2212), .op(n12031) );
  nand2_1 U13946 ( .ip1(\CORTEXM0DS_INST/u_logic/H0gvx4 ), .ip2(n2198), .op(
        n12030) );
  nand2_1 U13947 ( .ip1(n12031), .ip2(n12030), .op(n6113) );
  nand2_1 U13948 ( .ip1(n2212), .ip2(n2197), .op(
        \CORTEXM0DS_INST/u_logic/Xmywx4 ) );
  nor3_1 U13949 ( .ip1(n12034), .ip2(n12033), .ip3(n12032), .op(n12053) );
  nor3_1 U13950 ( .ip1(n12053), .ip2(n12559), .ip3(n12446), .op(n12037) );
  nor2_1 U13951 ( .ip1(n12035), .ip2(n12554), .op(n12036) );
  not_ab_or_c_or_d U13952 ( .ip1(\CORTEXM0DS_INST/u_logic/D69vx4 ), .ip2(
        n12052), .ip3(n12037), .ip4(n12036), .op(n12038) );
  or2_1 U13953 ( .ip1(n12038), .ip2(n5780), .op(n12041) );
  nand2_1 U13954 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n12058), .op(
        n12039) );
  or2_1 U13955 ( .ip1(n12039), .ip2(n5780), .op(n12040) );
  nand2_1 U13956 ( .ip1(n12041), .ip2(n12040), .op(n12045) );
  nor2_1 U13957 ( .ip1(n12043), .ip2(n12042), .op(n12044) );
  ab_or_c_or_d U13958 ( .ip1(n5780), .ip2(\CORTEXM0DS_INST/u_logic/Cq9vx4 ), 
        .ip3(n12045), .ip4(n12044), .op(n6112) );
  nor2_1 U13959 ( .ip1(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip2(n12065), .op(
        n12047) );
  nor2_1 U13960 ( .ip1(n12047), .ip2(n12046), .op(n12048) );
  nor4_1 U13961 ( .ip1(n12051), .ip2(n12050), .ip3(n12049), .ip4(n12048), .op(
        n12063) );
  nand2_1 U13962 ( .ip1(\CORTEXM0DS_INST/u_logic/W49vx4 ), .ip2(n12052), .op(
        n12061) );
  nand2_1 U13963 ( .ip1(\CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Vsevx4 ), .op(n12451) );
  nor2_1 U13964 ( .ip1(n12053), .ip2(n12451), .op(n12057) );
  not_ab_or_c_or_d U13965 ( .ip1(n12055), .ip2(n12054), .ip3(
        \CORTEXM0DS_INST/u_logic/Aj9vx4 ), .ip4(n12584), .op(n12056) );
  not_ab_or_c_or_d U13966 ( .ip1(n12058), .ip2(
        \CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip3(n12057), .ip4(n12056), .op(
        n12060) );
  nand3_1 U13967 ( .ip1(n12061), .ip2(n12060), .ip3(n12059), .op(n12062) );
  not_ab_or_c_or_d U13968 ( .ip1(\CORTEXM0DS_INST/u_logic/P39vx4 ), .ip2(
        n12064), .ip3(n12063), .ip4(n12062), .op(n12066) );
  mux2_1 U13969 ( .ip1(n12066), .ip2(n12065), .s(n5780), .op(n12070) );
  nand2_1 U13970 ( .ip1(n12068), .ip2(n12067), .op(n12069) );
  nand2_1 U13971 ( .ip1(n12070), .ip2(n12069), .op(n6111) );
  nor2_1 U13972 ( .ip1(n12072), .ip2(n12071), .op(n12077) );
  not_ab_or_c_or_d U13973 ( .ip1(\CORTEXM0DS_INST/u_logic/Kg9vx4 ), .ip2(
        n12075), .ip3(n12074), .ip4(n12073), .op(n12076) );
  not_ab_or_c_or_d U13974 ( .ip1(n12079), .ip2(n12078), .ip3(n12077), .ip4(
        n12076), .op(n12087) );
  inv_1 U13975 ( .ip(n12080), .op(n12085) );
  nor2_1 U13976 ( .ip1(n12082), .ip2(n12081), .op(n12084) );
  not_ab_or_c_or_d U13977 ( .ip1(n12085), .ip2(n10865), .ip3(n12084), .ip4(
        n12083), .op(n12086) );
  nand3_1 U13978 ( .ip1(n12088), .ip2(n12087), .ip3(n12086), .op(n2168) );
  nand3_1 U13979 ( .ip1(n12642), .ip2(n12090), .ip3(n12089), .op(n12093) );
  nand2_1 U13980 ( .ip1(\CORTEXM0DS_INST/u_logic/I4gvx4 ), .ip2(n12091), .op(
        n12092) );
  nand2_1 U13981 ( .ip1(n12093), .ip2(n12092), .op(n6110) );
  not_ab_or_c_or_d U13982 ( .ip1(n12095), .ip2(n12686), .ip3(n5938), .ip4(
        n12094), .op(n12097) );
  or2_1 U13983 ( .ip1(n12097), .ip2(n12096), .op(n12098) );
  nand2_1 U13984 ( .ip1(n2136), .ip2(n12098), .op(n6109) );
  inv_1 U13985 ( .ip(n12099), .op(n12106) );
  inv_1 U13986 ( .ip(n12216), .op(n12102) );
  inv_1 U13987 ( .ip(n12308), .op(n12100) );
  not_ab_or_c_or_d U13988 ( .ip1(n12102), .ip2(n12101), .ip3(n12100), .ip4(
        n12305), .op(n12105) );
  nor2_1 U13989 ( .ip1(n12103), .ip2(n12309), .op(n12104) );
  not_ab_or_c_or_d U13990 ( .ip1(n12314), .ip2(n12106), .ip3(n12105), .ip4(
        n12104), .op(\CORTEXM0DS_INST/u_logic/Y92wx4 ) );
  nor2_1 U13991 ( .ip1(\CORTEXM0DS_INST/u_logic/Y92wx4 ), .ip2(n12317), .op(
        n12109) );
  inv_1 U13992 ( .ip(n2120), .op(n12315) );
  nor2_1 U13993 ( .ip1(n12107), .ip2(n12315), .op(n12108) );
  ab_or_c_or_d U13994 ( .ip1(n12321), .ip2(\CORTEXM0DS_INST/vis_pc [22]), 
        .ip3(n12109), .ip4(n12108), .op(n6107) );
  nand2_1 U13995 ( .ip1(\CORTEXM0DS_INST/u_logic/Jjdvx4 ), .ip2(n2120), .op(
        n12111) );
  nand2_1 U13996 ( .ip1(\CORTEXM0DS_INST/vis_pc [14]), .ip2(n12321), .op(
        n12110) );
  nand3_1 U13997 ( .ip1(n12111), .ip2(n2095), .ip3(n12110), .op(n6106) );
  not_ab_or_c_or_d U13998 ( .ip1(n12292), .ip2(n12113), .ip3(n12112), .ip4(
        n12305), .op(n12116) );
  nor2_1 U13999 ( .ip1(n12114), .ip2(n12295), .op(n12115) );
  not_ab_or_c_or_d U14000 ( .ip1(n12300), .ip2(n12117), .ip3(n12116), .ip4(
        n12115), .op(\CORTEXM0DS_INST/u_logic/Z6ovx4 ) );
  nor2_1 U14001 ( .ip1(\CORTEXM0DS_INST/u_logic/Z6ovx4 ), .ip2(n12317), .op(
        n12120) );
  nor2_1 U14002 ( .ip1(n12118), .ip2(n12315), .op(n12119) );
  ab_or_c_or_d U14003 ( .ip1(n12321), .ip2(\CORTEXM0DS_INST/vis_pc [7]), .ip3(
        n12120), .ip4(n12119), .op(n6105) );
  nor2_1 U14004 ( .ip1(n12122), .ip2(n12121), .op(n12130) );
  not_ab_or_c_or_d U14005 ( .ip1(n12122), .ip2(n12121), .ip3(n12130), .ip4(
        n12305), .op(n12125) );
  nor2_1 U14006 ( .ip1(n12123), .ip2(n12295), .op(n12124) );
  not_ab_or_c_or_d U14007 ( .ip1(n12300), .ip2(n12126), .ip3(n12125), .ip4(
        n12124), .op(\CORTEXM0DS_INST/u_logic/Jxovx4 ) );
  inv_1 U14008 ( .ip(\CORTEXM0DS_INST/u_logic/Jxovx4 ), .op(n2069) );
  nand2_1 U14009 ( .ip1(\CORTEXM0DS_INST/u_logic/Gcdvx4 ), .ip2(n2120), .op(
        n12129) );
  nand2_1 U14010 ( .ip1(n12691), .ip2(n2069), .op(n12128) );
  nand2_1 U14011 ( .ip1(\CORTEXM0DS_INST/vis_pc [9]), .ip2(n12321), .op(n12127) );
  nand3_1 U14012 ( .ip1(n12129), .ip2(n12128), .ip3(n12127), .op(n6103) );
  inv_1 U14013 ( .ip(n12130), .op(n12132) );
  nand2_1 U14014 ( .ip1(\CORTEXM0DS_INST/vis_pc [10]), .ip2(n12130), .op(
        n12143) );
  inv_1 U14015 ( .ip(n12143), .op(n12131) );
  not_ab_or_c_or_d U14016 ( .ip1(n12133), .ip2(n12132), .ip3(n12131), .ip4(
        n12305), .op(n12136) );
  nor2_1 U14017 ( .ip1(n12134), .ip2(n12295), .op(n12135) );
  not_ab_or_c_or_d U14018 ( .ip1(n12300), .ip2(n12137), .ip3(n12136), .ip4(
        n12135), .op(\CORTEXM0DS_INST/u_logic/Owovx4 ) );
  inv_1 U14019 ( .ip(\CORTEXM0DS_INST/u_logic/Owovx4 ), .op(n2065) );
  nand2_1 U14020 ( .ip1(\CORTEXM0DS_INST/u_logic/Rddvx4 ), .ip2(n2120), .op(
        n12140) );
  nand2_1 U14021 ( .ip1(n12691), .ip2(n2065), .op(n12139) );
  nand2_1 U14022 ( .ip1(\CORTEXM0DS_INST/vis_pc [10]), .ip2(n12321), .op(
        n12138) );
  nand3_1 U14023 ( .ip1(n12140), .ip2(n12139), .ip3(n12138), .op(n6102) );
  nor2_1 U14024 ( .ip1(n12141), .ip2(n12295), .op(n12146) );
  inv_1 U14025 ( .ip(\CORTEXM0DS_INST/vis_pc [11]), .op(n12144) );
  not_ab_or_c_or_d U14026 ( .ip1(n12144), .ip2(n12143), .ip3(n12142), .ip4(
        n12305), .op(n12145) );
  not_ab_or_c_or_d U14027 ( .ip1(n12300), .ip2(n12147), .ip3(n12146), .ip4(
        n12145), .op(\CORTEXM0DS_INST/u_logic/Cqovx4 ) );
  nor2_1 U14028 ( .ip1(\CORTEXM0DS_INST/u_logic/Cqovx4 ), .ip2(n12317), .op(
        n12150) );
  nor2_1 U14029 ( .ip1(n12148), .ip2(n12315), .op(n12149) );
  ab_or_c_or_d U14030 ( .ip1(n12321), .ip2(\CORTEXM0DS_INST/vis_pc [11]), 
        .ip3(n12150), .ip4(n12149), .op(n6101) );
  nand2_1 U14031 ( .ip1(\CORTEXM0DS_INST/u_logic/Ngdvx4 ), .ip2(n2120), .op(
        n12152) );
  nand2_1 U14032 ( .ip1(\CORTEXM0DS_INST/vis_pc [12]), .ip2(n12321), .op(
        n12151) );
  nand3_1 U14033 ( .ip1(n12152), .ip2(n2060), .ip3(n12151), .op(n6100) );
  nand2_1 U14034 ( .ip1(\CORTEXM0DS_INST/u_logic/Yhdvx4 ), .ip2(n2120), .op(
        n12154) );
  nand2_1 U14035 ( .ip1(\CORTEXM0DS_INST/vis_pc [13]), .ip2(n12321), .op(
        n12153) );
  nand3_1 U14036 ( .ip1(n12154), .ip2(n2057), .ip3(n12153), .op(n6099) );
  inv_1 U14037 ( .ip(n12155), .op(n12158) );
  inv_1 U14038 ( .ip(n12167), .op(n12156) );
  not_ab_or_c_or_d U14039 ( .ip1(n12158), .ip2(n12157), .ip3(n12156), .ip4(
        n12305), .op(n12161) );
  nor2_1 U14040 ( .ip1(n12159), .ip2(n12295), .op(n12160) );
  not_ab_or_c_or_d U14041 ( .ip1(n12300), .ip2(n12162), .ip3(n12161), .ip4(
        n12160), .op(\CORTEXM0DS_INST/u_logic/Vpovx4 ) );
  nor2_1 U14042 ( .ip1(\CORTEXM0DS_INST/u_logic/Vpovx4 ), .ip2(n12317), .op(
        n12165) );
  nor2_1 U14043 ( .ip1(n12163), .ip2(n12315), .op(n12164) );
  ab_or_c_or_d U14044 ( .ip1(n12321), .ip2(\CORTEXM0DS_INST/vis_pc [15]), 
        .ip3(n12165), .ip4(n12164), .op(n6098) );
  not_ab_or_c_or_d U14045 ( .ip1(n12167), .ip2(n12166), .ip3(n12176), .ip4(
        n12305), .op(n12170) );
  nor2_1 U14046 ( .ip1(n12168), .ip2(n12309), .op(n12169) );
  not_ab_or_c_or_d U14047 ( .ip1(n12314), .ip2(n12171), .ip3(n12170), .ip4(
        n12169), .op(\CORTEXM0DS_INST/u_logic/Bv0wx4 ) );
  nor2_1 U14048 ( .ip1(\CORTEXM0DS_INST/u_logic/Bv0wx4 ), .ip2(n12317), .op(
        n12174) );
  nor2_1 U14049 ( .ip1(n12172), .ip2(n12315), .op(n12173) );
  ab_or_c_or_d U14050 ( .ip1(n12321), .ip2(\CORTEXM0DS_INST/vis_pc [16]), 
        .ip3(n12174), .ip4(n12173), .op(n6097) );
  nor2_1 U14051 ( .ip1(n12175), .ip2(n12295), .op(n12181) );
  inv_1 U14052 ( .ip(\CORTEXM0DS_INST/vis_pc [17]), .op(n12179) );
  inv_1 U14053 ( .ip(n12176), .op(n12178) );
  nand2_1 U14054 ( .ip1(\CORTEXM0DS_INST/vis_pc [17]), .ip2(n12176), .op(
        n12187) );
  inv_1 U14055 ( .ip(n12187), .op(n12177) );
  not_ab_or_c_or_d U14056 ( .ip1(n12179), .ip2(n12178), .ip3(n12177), .ip4(
        n12305), .op(n12180) );
  not_ab_or_c_or_d U14057 ( .ip1(n12300), .ip2(n12182), .ip3(n12181), .ip4(
        n12180), .op(\CORTEXM0DS_INST/u_logic/Fq0wx4 ) );
  nor2_1 U14058 ( .ip1(\CORTEXM0DS_INST/u_logic/Fq0wx4 ), .ip2(n12317), .op(
        n12185) );
  nor2_1 U14059 ( .ip1(n12183), .ip2(n12315), .op(n12184) );
  ab_or_c_or_d U14060 ( .ip1(n12321), .ip2(\CORTEXM0DS_INST/vis_pc [17]), 
        .ip3(n12185), .ip4(n12184), .op(n6096) );
  inv_1 U14061 ( .ip(n12197), .op(n12186) );
  not_ab_or_c_or_d U14062 ( .ip1(n12188), .ip2(n12187), .ip3(n12186), .ip4(
        n12305), .op(n12191) );
  nor2_1 U14063 ( .ip1(n12189), .ip2(n12309), .op(n12190) );
  not_ab_or_c_or_d U14064 ( .ip1(n12314), .ip2(n12192), .ip3(n12191), .ip4(
        n12190), .op(\CORTEXM0DS_INST/u_logic/Ql0wx4 ) );
  nor2_1 U14065 ( .ip1(\CORTEXM0DS_INST/u_logic/Ql0wx4 ), .ip2(n12317), .op(
        n12195) );
  nor2_1 U14066 ( .ip1(n12193), .ip2(n12315), .op(n12194) );
  ab_or_c_or_d U14067 ( .ip1(n12321), .ip2(\CORTEXM0DS_INST/vis_pc [18]), 
        .ip3(n12195), .ip4(n12194), .op(n6095) );
  not_ab_or_c_or_d U14068 ( .ip1(n12197), .ip2(n12196), .ip3(n12205), .ip4(
        n12305), .op(n12200) );
  nor2_1 U14069 ( .ip1(n12198), .ip2(n12309), .op(n12199) );
  not_ab_or_c_or_d U14070 ( .ip1(n12314), .ip2(n12201), .ip3(n12200), .ip4(
        n12199), .op(\CORTEXM0DS_INST/u_logic/Ug0wx4 ) );
  nor2_1 U14071 ( .ip1(\CORTEXM0DS_INST/u_logic/Ug0wx4 ), .ip2(n12317), .op(
        n12204) );
  nor2_1 U14072 ( .ip1(n12202), .ip2(n12315), .op(n12203) );
  ab_or_c_or_d U14073 ( .ip1(n12321), .ip2(\CORTEXM0DS_INST/vis_pc [19]), 
        .ip3(n12204), .ip4(n12203), .op(n6094) );
  inv_1 U14074 ( .ip(n12205), .op(n12208) );
  inv_1 U14075 ( .ip(n12218), .op(n12206) );
  not_ab_or_c_or_d U14076 ( .ip1(n12208), .ip2(n12207), .ip3(n12206), .ip4(
        n12305), .op(n12211) );
  nor2_1 U14077 ( .ip1(n12209), .ip2(n12309), .op(n12210) );
  not_ab_or_c_or_d U14078 ( .ip1(n12314), .ip2(n12212), .ip3(n12211), .ip4(
        n12210), .op(\CORTEXM0DS_INST/u_logic/Fc0wx4 ) );
  nor2_1 U14079 ( .ip1(\CORTEXM0DS_INST/u_logic/Fc0wx4 ), .ip2(n12317), .op(
        n12215) );
  nor2_1 U14080 ( .ip1(n12213), .ip2(n12315), .op(n12214) );
  ab_or_c_or_d U14081 ( .ip1(n12321), .ip2(\CORTEXM0DS_INST/vis_pc [20]), 
        .ip3(n12215), .ip4(n12214), .op(n6093) );
  not_ab_or_c_or_d U14082 ( .ip1(n12218), .ip2(n12217), .ip3(n12216), .ip4(
        n12305), .op(n12221) );
  nor2_1 U14083 ( .ip1(n12219), .ip2(n12309), .op(n12220) );
  not_ab_or_c_or_d U14084 ( .ip1(n12314), .ip2(n12222), .ip3(n12221), .ip4(
        n12220), .op(\CORTEXM0DS_INST/u_logic/C70wx4 ) );
  nor2_1 U14085 ( .ip1(\CORTEXM0DS_INST/u_logic/C70wx4 ), .ip2(n12317), .op(
        n12225) );
  nor2_1 U14086 ( .ip1(n12223), .ip2(n12315), .op(n12224) );
  ab_or_c_or_d U14087 ( .ip1(n12321), .ip2(\CORTEXM0DS_INST/vis_pc [21]), 
        .ip3(n12225), .ip4(n12224), .op(n6092) );
  inv_1 U14088 ( .ip(n12226), .op(n12229) );
  inv_1 U14089 ( .ip(\CORTEXM0DS_INST/vis_pc [4]), .op(n12228) );
  inv_1 U14090 ( .ip(n12239), .op(n12227) );
  not_ab_or_c_or_d U14091 ( .ip1(n12229), .ip2(n12228), .ip3(n12227), .ip4(
        n12305), .op(n12232) );
  and2_1 U14092 ( .ip1(n12230), .ip2(n12300), .op(n12231) );
  not_ab_or_c_or_d U14093 ( .ip1(n12314), .ip2(n12233), .ip3(n12232), .ip4(
        n12231), .op(\CORTEXM0DS_INST/u_logic/Rxzvx4 ) );
  nor2_1 U14094 ( .ip1(n12234), .ip2(n12315), .op(n12236) );
  nor2_1 U14095 ( .ip1(\CORTEXM0DS_INST/u_logic/Rxzvx4 ), .ip2(n12317), .op(
        n12235) );
  not_ab_or_c_or_d U14096 ( .ip1(n12320), .ip2(\CORTEXM0DS_INST/vis_ipsr [5]), 
        .ip3(n12236), .ip4(n12235), .op(n12238) );
  nand2_1 U14097 ( .ip1(\CORTEXM0DS_INST/vis_pc [4]), .ip2(n12321), .op(n12237) );
  nand2_1 U14098 ( .ip1(n12238), .ip2(n12237), .op(n6089) );
  not_ab_or_c_or_d U14099 ( .ip1(n12239), .ip2(n12244), .ip3(n12291), .ip4(
        n12305), .op(n12242) );
  nor2_1 U14100 ( .ip1(n12240), .ip2(n12295), .op(n12241) );
  not_ab_or_c_or_d U14101 ( .ip1(n12300), .ip2(n12243), .ip3(n12242), .ip4(
        n12241), .op(\CORTEXM0DS_INST/u_logic/Hszvx4 ) );
  nor2_1 U14102 ( .ip1(\CORTEXM0DS_INST/u_logic/Hszvx4 ), .ip2(n12317), .op(
        n12246) );
  inv_1 U14103 ( .ip(n12321), .op(n12301) );
  nor2_1 U14104 ( .ip1(n12244), .ip2(n12301), .op(n12245) );
  ab_or_c_or_d U14105 ( .ip1(n2120), .ip2(\CORTEXM0DS_INST/u_logic/S6dvx4 ), 
        .ip3(n12246), .ip4(n12245), .op(n6088) );
  inv_1 U14106 ( .ip(n12306), .op(n12249) );
  inv_1 U14107 ( .ip(n12258), .op(n12247) );
  not_ab_or_c_or_d U14108 ( .ip1(n12249), .ip2(n12248), .ip3(n12247), .ip4(
        n12305), .op(n12252) );
  nor2_1 U14109 ( .ip1(n12250), .ip2(n12309), .op(n12251) );
  not_ab_or_c_or_d U14110 ( .ip1(n12314), .ip2(n12253), .ip3(n12252), .ip4(
        n12251), .op(\CORTEXM0DS_INST/u_logic/Rnovx4 ) );
  nor2_1 U14111 ( .ip1(\CORTEXM0DS_INST/u_logic/Rnovx4 ), .ip2(n12317), .op(
        n12256) );
  nor2_1 U14112 ( .ip1(n12254), .ip2(n12315), .op(n12255) );
  ab_or_c_or_d U14113 ( .ip1(n12321), .ip2(\CORTEXM0DS_INST/vis_pc [24]), 
        .ip3(n12256), .ip4(n12255), .op(n6087) );
  not_ab_or_c_or_d U14114 ( .ip1(n12258), .ip2(n12257), .ip3(n12266), .ip4(
        n12305), .op(n12261) );
  nor2_1 U14115 ( .ip1(n12259), .ip2(n12295), .op(n12260) );
  not_ab_or_c_or_d U14116 ( .ip1(n12300), .ip2(n12262), .ip3(n12261), .ip4(
        n12260), .op(\CORTEXM0DS_INST/u_logic/Nhzvx4 ) );
  nor2_1 U14117 ( .ip1(\CORTEXM0DS_INST/u_logic/Nhzvx4 ), .ip2(n12317), .op(
        n12265) );
  nor2_1 U14118 ( .ip1(n12263), .ip2(n12315), .op(n12264) );
  ab_or_c_or_d U14119 ( .ip1(n12321), .ip2(\CORTEXM0DS_INST/vis_pc [25]), 
        .ip3(n12265), .ip4(n12264), .op(n6086) );
  inv_1 U14120 ( .ip(n12266), .op(n12270) );
  inv_1 U14121 ( .ip(\CORTEXM0DS_INST/vis_pc [26]), .op(n12269) );
  inv_1 U14122 ( .ip(n12267), .op(n12268) );
  not_ab_or_c_or_d U14123 ( .ip1(n12270), .ip2(n12269), .ip3(n12268), .ip4(
        n12305), .op(n12273) );
  nor2_1 U14124 ( .ip1(n12271), .ip2(n12309), .op(n12272) );
  not_ab_or_c_or_d U14125 ( .ip1(n12314), .ip2(n12274), .ip3(n12273), .ip4(
        n12272), .op(\CORTEXM0DS_INST/u_logic/Vezvx4 ) );
  nor2_1 U14126 ( .ip1(\CORTEXM0DS_INST/u_logic/Vezvx4 ), .ip2(n12317), .op(
        n12277) );
  nor2_1 U14127 ( .ip1(n12275), .ip2(n12315), .op(n12276) );
  ab_or_c_or_d U14128 ( .ip1(n12321), .ip2(\CORTEXM0DS_INST/vis_pc [26]), 
        .ip3(n12277), .ip4(n12276), .op(n6085) );
  or2_1 U14129 ( .ip1(n12278), .ip2(n12279), .op(n12282) );
  or2_1 U14130 ( .ip1(n12280), .ip2(n12279), .op(n12281) );
  nand2_1 U14131 ( .ip1(n12282), .ip2(n12281), .op(n12283) );
  nor2_1 U14132 ( .ip1(n12284), .ip2(n12283), .op(n12285) );
  nor2_1 U14133 ( .ip1(n12286), .ip2(n12285), .op(n12287) );
  nor2_1 U14134 ( .ip1(n12287), .ip2(n12317), .op(n12290) );
  nor2_1 U14135 ( .ip1(n12288), .ip2(n12315), .op(n12289) );
  ab_or_c_or_d U14136 ( .ip1(n12320), .ip2(\CORTEXM0DS_INST/vis_ipsr [0]), 
        .ip3(n12290), .ip4(n12289), .op(n6082) );
  inv_1 U14137 ( .ip(n12291), .op(n12294) );
  inv_1 U14138 ( .ip(n12292), .op(n12293) );
  not_ab_or_c_or_d U14139 ( .ip1(n12294), .ip2(n12302), .ip3(n12293), .ip4(
        n12305), .op(n12298) );
  nor2_1 U14140 ( .ip1(n12296), .ip2(n12295), .op(n12297) );
  not_ab_or_c_or_d U14141 ( .ip1(n12300), .ip2(n12299), .ip3(n12298), .ip4(
        n12297), .op(\CORTEXM0DS_INST/u_logic/S4qvx4 ) );
  nor2_1 U14142 ( .ip1(\CORTEXM0DS_INST/u_logic/S4qvx4 ), .ip2(n12317), .op(
        n12304) );
  nor2_1 U14143 ( .ip1(n12302), .ip2(n12301), .op(n12303) );
  ab_or_c_or_d U14144 ( .ip1(n2120), .ip2(\CORTEXM0DS_INST/u_logic/C8dvx4 ), 
        .ip3(n12304), .ip4(n12303), .op(n6080) );
  not_ab_or_c_or_d U14145 ( .ip1(n12308), .ip2(n12307), .ip3(n12306), .ip4(
        n12305), .op(n12312) );
  nor2_1 U14146 ( .ip1(n12310), .ip2(n12309), .op(n12311) );
  not_ab_or_c_or_d U14147 ( .ip1(n12314), .ip2(n12313), .ip3(n12312), .ip4(
        n12311), .op(\CORTEXM0DS_INST/u_logic/Y1pvx4 ) );
  nor2_1 U14148 ( .ip1(n12316), .ip2(n12315), .op(n12319) );
  nor2_1 U14149 ( .ip1(\CORTEXM0DS_INST/u_logic/Y1pvx4 ), .ip2(n12317), .op(
        n12318) );
  not_ab_or_c_or_d U14150 ( .ip1(n12320), .ip2(\CORTEXM0DS_INST/cm0_xpsr[24] ), 
        .ip3(n12319), .ip4(n12318), .op(n12323) );
  nand2_1 U14151 ( .ip1(\CORTEXM0DS_INST/vis_pc [23]), .ip2(n12321), .op(
        n12322) );
  nand2_1 U14152 ( .ip1(n12323), .ip2(n12322), .op(n6077) );
  inv_1 U14153 ( .ip(n12324), .op(n12350) );
  nor2_1 U14154 ( .ip1(\CORTEXM0DS_INST/u_logic/Mcgvx4 ), .ip2(n12325), .op(
        n12348) );
  nor2_1 U14155 ( .ip1(n12625), .ip2(n12326), .op(n12346) );
  nand3_1 U14156 ( .ip1(\CORTEXM0DS_INST/u_logic/Cf9vx4 ), .ip2(n12328), .ip3(
        n12327), .op(n12331) );
  not_ab_or_c_or_d U14157 ( .ip1(n12332), .ip2(n12331), .ip3(n12330), .ip4(
        n12329), .op(n12345) );
  not_ab_or_c_or_d U14158 ( .ip1(n12336), .ip2(n12335), .ip3(n12334), .ip4(
        n12333), .op(n12344) );
  nand3_1 U14159 ( .ip1(n12339), .ip2(n12338), .ip3(n12337), .op(n12340) );
  nand3_1 U14160 ( .ip1(n12342), .ip2(n12341), .ip3(n12340), .op(n12343) );
  or4_1 U14161 ( .ip1(n12346), .ip2(n12345), .ip3(n12344), .ip4(n12343), .op(
        n12347) );
  not_ab_or_c_or_d U14162 ( .ip1(n12350), .ip2(n12349), .ip3(n12348), .ip4(
        n12347), .op(n12355) );
  or2_1 U14163 ( .ip1(n12352), .ip2(n12351), .op(n12354) );
  nand3_1 U14164 ( .ip1(n12355), .ip2(n12354), .ip3(n12353), .op(n1789) );
  nand2_1 U14165 ( .ip1(n12356), .ip2(n1770), .op(n12361) );
  nand2_1 U14166 ( .ip1(\CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip2(n12366), .op(
        n12358) );
  nand2_1 U14167 ( .ip1(\CORTEXM0DS_INST/u_logic/I29vx4 ), .ip2(n12367), .op(
        n12357) );
  nand4_1 U14168 ( .ip1(n12384), .ip2(n12359), .ip3(n12358), .ip4(n12357), 
        .op(n12360) );
  nand2_1 U14169 ( .ip1(n12361), .ip2(n12360), .op(n12364) );
  nand3_1 U14170 ( .ip1(n12362), .ip2(n12389), .ip3(n12388), .op(n12363) );
  nand2_1 U14171 ( .ip1(n12364), .ip2(n12363), .op(n6076) );
  nand2_1 U14172 ( .ip1(n12365), .ip2(n1770), .op(n12372) );
  nand2_1 U14173 ( .ip1(\CORTEXM0DS_INST/u_logic/Fb9vx4 ), .ip2(n12366), .op(
        n12370) );
  nand2_1 U14174 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n12381), .op(
        n12369) );
  nand2_1 U14175 ( .ip1(\CORTEXM0DS_INST/u_logic/B19vx4 ), .ip2(n12367), .op(
        n12368) );
  nand4_1 U14176 ( .ip1(n12384), .ip2(n12370), .ip3(n12369), .ip4(n12368), 
        .op(n12371) );
  nand2_1 U14177 ( .ip1(n12372), .ip2(n12371), .op(n12375) );
  nand3_1 U14178 ( .ip1(n12373), .ip2(n12389), .ip3(n12388), .op(n12374) );
  nand2_1 U14179 ( .ip1(n12375), .ip2(n12374), .op(n6075) );
  nand2_1 U14180 ( .ip1(n12376), .ip2(n1770), .op(n12387) );
  nor2_1 U14181 ( .ip1(n12592), .ip2(n12377), .op(n12380) );
  nor2_1 U14182 ( .ip1(n12378), .ip2(n12588), .op(n12379) );
  not_ab_or_c_or_d U14183 ( .ip1(n12381), .ip2(
        \CORTEXM0DS_INST/u_logic/Mc9vx4 ), .ip3(n12380), .ip4(n12379), .op(
        n12385) );
  or2_1 U14184 ( .ip1(n12550), .ip2(n12382), .op(n12383) );
  nand3_1 U14185 ( .ip1(n12385), .ip2(n12384), .ip3(n12383), .op(n12386) );
  nand2_1 U14186 ( .ip1(n12387), .ip2(n12386), .op(n12392) );
  nand3_1 U14187 ( .ip1(n12390), .ip2(n12389), .ip3(n12388), .op(n12391) );
  nand2_1 U14188 ( .ip1(n12392), .ip2(n12391), .op(n6074) );
  nand3_1 U14189 ( .ip1(n12394), .ip2(\CORTEXM0DS_INST/u_logic/Fjgvx4 ), .ip3(
        n12393), .op(n12398) );
  nand3_1 U14190 ( .ip1(n12396), .ip2(n12395), .ip3(n12645), .op(n12397) );
  nand2_1 U14191 ( .ip1(n12398), .ip2(n12397), .op(n12399) );
  nand3_1 U14192 ( .ip1(n12402), .ip2(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip3(
        n12399), .op(n12401) );
  nand2_1 U14193 ( .ip1(\CORTEXM0DS_INST/u_logic/Mk8vx4 ), .ip2(n1709), .op(
        n12400) );
  nand2_1 U14194 ( .ip1(n12401), .ip2(n12400), .op(n6072) );
  nand2_1 U14195 ( .ip1(\CORTEXM0DS_INST/u_logic/Ul8vx4 ), .ip2(n1709), .op(
        n12410) );
  nand3_1 U14196 ( .ip1(\CORTEXM0DS_INST/u_logic/Rkgvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Pp8vx4 ), .ip3(n12405), .op(n12407) );
  nand4_1 U14197 ( .ip1(n12405), .ip2(n12404), .ip3(n12403), .ip4(n12402), 
        .op(n12406) );
  nand2_1 U14198 ( .ip1(n12407), .ip2(n12406), .op(n12408) );
  nand2_1 U14199 ( .ip1(n12642), .ip2(n12408), .op(n12409) );
  nand2_1 U14200 ( .ip1(n12410), .ip2(n12409), .op(n6071) );
  nand2_1 U14201 ( .ip1(n5938), .ip2(\CORTEXM0DS_INST/u_logic/N6hvx4 ), .op(
        n12419) );
  or2_1 U14202 ( .ip1(n1671), .ip2(n1672), .op(n12413) );
  nand3_1 U14203 ( .ip1(n1667), .ip2(n1668), .ip3(
        \CORTEXM0DS_INST/u_logic/Yuovx4 ), .op(n12411) );
  nand2_1 U14204 ( .ip1(n1670), .ip2(n12411), .op(n12412) );
  nand4_1 U14205 ( .ip1(n1675), .ip2(\CORTEXM0DS_INST/u_logic/Ekovx4 ), .ip3(
        n12413), .ip4(n12412), .op(n12415) );
  nand3_1 U14206 ( .ip1(n1672), .ip2(n1664), .ip3(n1663), .op(n12414) );
  not_ab_or_c_or_d U14207 ( .ip1(n12415), .ip2(n12414), .ip3(n1678), .ip4(
        n1677), .op(n12416) );
  nand3_1 U14208 ( .ip1(\CORTEXM0DS_INST/u_logic/Vpovx4 ), .ip2(n12416), .ip3(
        \CORTEXM0DS_INST/u_logic/Rnovx4 ), .op(n12417) );
  nand2_1 U14209 ( .ip1(n3127), .ip2(n12417), .op(n12427) );
  nand2_1 U14210 ( .ip1(\CORTEXM0DS_INST/u_logic/Yuovx4 ), .ip2(n3127), .op(
        n12418) );
  nand3_1 U14211 ( .ip1(n12419), .ip2(n12427), .ip3(n12418), .op(n6070) );
  inv_1 U14212 ( .ip(n12427), .op(n12425) );
  nor2_1 U14213 ( .ip1(\CORTEXM0DS_INST/u_logic/Ekovx4 ), .ip2(n1691), .op(
        n12420) );
  inv_1 U14214 ( .ip(n3127), .op(n12423) );
  not_ab_or_c_or_d U14215 ( .ip1(\CORTEXM0DS_INST/u_logic/Ekovx4 ), .ip2(n1691), .ip3(n12420), .ip4(n12423), .op(n12421) );
  ab_or_c_or_d U14216 ( .ip1(\CORTEXM0DS_INST/u_logic/Z7hvx4 ), .ip2(n5938), 
        .ip3(n12425), .ip4(n12421), .op(n6069) );
  nor2_1 U14217 ( .ip1(n1687), .ip2(n12423), .op(n12422) );
  ab_or_c_or_d U14218 ( .ip1(\CORTEXM0DS_INST/u_logic/L9hvx4 ), .ip2(n5938), 
        .ip3(n12425), .ip4(n12422), .op(n6068) );
  nor2_1 U14219 ( .ip1(n1685), .ip2(n12423), .op(n12424) );
  ab_or_c_or_d U14220 ( .ip1(\CORTEXM0DS_INST/u_logic/Xahvx4 ), .ip2(n5938), 
        .ip3(n12425), .ip4(n12424), .op(n6067) );
  nand2_1 U14221 ( .ip1(n5938), .ip2(\CORTEXM0DS_INST/u_logic/B5hvx4 ), .op(
        n12428) );
  nand2_1 U14222 ( .ip1(n3127), .ip2(\CORTEXM0DS_INST/u_logic/Z6ovx4 ), .op(
        n12426) );
  nand3_1 U14223 ( .ip1(n12428), .ip2(n12427), .ip3(n12426), .op(n6066) );
  inv_1 U14224 ( .ip(n1851), .op(\CORTEXM0DS_INST/u_logic/Fvovx4 ) );
  mux2_1 U14225 ( .ip1(n2212), .ip2(\CORTEXM0DS_INST/u_logic/Xyfvx4 ), .s(
        n5938), .op(n6065) );
  mux2_1 U14226 ( .ip1(n12429), .ip2(\CORTEXM0DS_INST/cm0_primask[0] ), .s(
        n5938), .op(n6064) );
  nand2_1 U14227 ( .ip1(n12457), .ip2(n12472), .op(n12432) );
  nor2_1 U14228 ( .ip1(n12472), .ip2(n12430), .op(n12443) );
  nand2_1 U14229 ( .ip1(\CORTEXM0DS_INST/u_logic/Hnevx4 ), .ip2(n12443), .op(
        n12431) );
  nand3_1 U14230 ( .ip1(n12432), .ip2(n1515), .ip3(n12431), .op(n6063) );
  inv_1 U14231 ( .ip(n12464), .op(n12453) );
  nand2_1 U14232 ( .ip1(n12472), .ip2(n12453), .op(n12434) );
  nand2_1 U14233 ( .ip1(n12443), .ip2(\CORTEXM0DS_INST/u_logic/Roevx4 ), .op(
        n12433) );
  nand3_1 U14234 ( .ip1(n12434), .ip2(n1510), .ip3(n12433), .op(n6062) );
  nand2_1 U14235 ( .ip1(n12466), .ip2(n12472), .op(n12436) );
  nand2_1 U14236 ( .ip1(n12443), .ip2(\CORTEXM0DS_INST/u_logic/Bqevx4 ), .op(
        n12435) );
  nand3_1 U14237 ( .ip1(n12436), .ip2(n1506), .ip3(n12435), .op(n6061) );
  nand2_1 U14238 ( .ip1(n12465), .ip2(n12472), .op(n12438) );
  nand2_1 U14239 ( .ip1(n12443), .ip2(\CORTEXM0DS_INST/u_logic/Lrevx4 ), .op(
        n12437) );
  nand3_1 U14240 ( .ip1(n12438), .ip2(n1505), .ip3(n12437), .op(n6060) );
  nor2_1 U14241 ( .ip1(n12440), .ip2(n12439), .op(n12452) );
  nand2_1 U14242 ( .ip1(n12452), .ip2(n12472), .op(n12442) );
  nand2_1 U14243 ( .ip1(n12443), .ip2(\CORTEXM0DS_INST/u_logic/Vsevx4 ), .op(
        n12441) );
  nand3_1 U14244 ( .ip1(n12442), .ip2(n1501), .ip3(n12441), .op(n6059) );
  nand2_1 U14245 ( .ip1(n12443), .ip2(\CORTEXM0DS_INST/u_logic/Fuevx4 ), .op(
        n12444) );
  nand2_1 U14246 ( .ip1(n1497), .ip2(n12444), .op(n6058) );
  inv_1 U14247 ( .ip(n4814), .op(n12510) );
  nand2_1 U14248 ( .ip1(\CORTEXM0DS_INST/u_logic/Pvevx4 ), .ip2(n12510), .op(
        n12474) );
  nor4_1 U14249 ( .ip1(\CORTEXM0DS_INST/u_logic/O2fvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/D1fvx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Tzevx4 ), .ip4(
        \CORTEXM0DS_INST/u_logic/Jyevx4 ), .op(n12445) );
  or2_1 U14250 ( .ip1(n12445), .ip2(n12446), .op(n12449) );
  nor4_1 U14251 ( .ip1(\CORTEXM0DS_INST/u_logic/Pvevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Zwevx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/K5fvx4 ), .ip4(
        \CORTEXM0DS_INST/u_logic/Z3fvx4 ), .op(n12447) );
  or2_1 U14252 ( .ip1(n12447), .ip2(n12446), .op(n12448) );
  nand2_1 U14253 ( .ip1(n12449), .ip2(n12448), .op(n12644) );
  inv_1 U14254 ( .ip(\CORTEXM0DS_INST/u_logic/Pvevx4 ), .op(n12563) );
  nor2_1 U14255 ( .ip1(n12452), .ip2(n12451), .op(n12450) );
  not_ab_or_c_or_d U14256 ( .ip1(n12452), .ip2(n12451), .ip3(
        \CORTEXM0DS_INST/u_logic/Fuevx4 ), .ip4(n12450), .op(n12470) );
  nor2_1 U14257 ( .ip1(n12457), .ip2(n12454), .op(n12463) );
  or2_1 U14258 ( .ip1(n12457), .ip2(n12453), .op(n12456) );
  or2_1 U14259 ( .ip1(n12454), .ip2(n12453), .op(n12455) );
  nand2_1 U14260 ( .ip1(n12456), .ip2(n12455), .op(n12461) );
  or2_1 U14261 ( .ip1(n12457), .ip2(n12539), .op(n12459) );
  or2_1 U14262 ( .ip1(n12534), .ip2(n12539), .op(n12458) );
  nand2_1 U14263 ( .ip1(n12459), .ip2(n12458), .op(n12460) );
  nor2_1 U14264 ( .ip1(n12461), .ip2(n12460), .op(n12462) );
  not_ab_or_c_or_d U14265 ( .ip1(\CORTEXM0DS_INST/u_logic/Roevx4 ), .ip2(
        n12464), .ip3(n12463), .ip4(n12462), .op(n12469) );
  mux2_1 U14266 ( .ip1(n12549), .ip2(\CORTEXM0DS_INST/u_logic/Lrevx4 ), .s(
        n12465), .op(n12468) );
  mux2_1 U14267 ( .ip1(n12545), .ip2(\CORTEXM0DS_INST/u_logic/Bqevx4 ), .s(
        n12466), .op(n12467) );
  nand4_1 U14268 ( .ip1(n12470), .ip2(n12469), .ip3(n12468), .ip4(n12467), 
        .op(n12471) );
  nand2_1 U14269 ( .ip1(n12472), .ip2(n12471), .op(n12507) );
  nand3_1 U14270 ( .ip1(n12644), .ip2(n12563), .ip3(n12507), .op(n12473) );
  nand3_1 U14271 ( .ip1(n12474), .ip2(n1495), .ip3(n12473), .op(n6057) );
  nand2_1 U14272 ( .ip1(n12510), .ip2(\CORTEXM0DS_INST/u_logic/Zwevx4 ), .op(
        n12478) );
  nand3_1 U14273 ( .ip1(\CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Zwevx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Pvevx4 ), .op(n12475) );
  inv_1 U14274 ( .ip(\CORTEXM0DS_INST/u_logic/Zwevx4 ), .op(n12569) );
  nand3_1 U14275 ( .ip1(n12644), .ip2(n12563), .ip3(n12569), .op(n12479) );
  nand2_1 U14276 ( .ip1(n12475), .ip2(n12479), .op(n12476) );
  nand2_1 U14277 ( .ip1(n12507), .ip2(n12476), .op(n12477) );
  nand3_1 U14278 ( .ip1(n12478), .ip2(n1491), .ip3(n12477), .op(n6056) );
  nand2_1 U14279 ( .ip1(n12510), .ip2(\CORTEXM0DS_INST/u_logic/Jyevx4 ), .op(
        n12483) );
  nand3_1 U14280 ( .ip1(n12479), .ip2(\CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip3(
        \CORTEXM0DS_INST/u_logic/Jyevx4 ), .op(n12480) );
  nor2_1 U14281 ( .ip1(\CORTEXM0DS_INST/u_logic/Jyevx4 ), .ip2(n12479), .op(
        n12497) );
  inv_1 U14282 ( .ip(n12497), .op(n12484) );
  nand2_1 U14283 ( .ip1(n12480), .ip2(n12484), .op(n12481) );
  nand2_1 U14284 ( .ip1(n12507), .ip2(n12481), .op(n12482) );
  nand3_1 U14285 ( .ip1(n12483), .ip2(n1488), .ip3(n12482), .op(n6055) );
  nand2_1 U14286 ( .ip1(n12510), .ip2(\CORTEXM0DS_INST/u_logic/Tzevx4 ), .op(
        n12487) );
  nand2_1 U14287 ( .ip1(\CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Tzevx4 ), .op(n12495) );
  xor2_1 U14288 ( .ip1(n12484), .ip2(n12495), .op(n12485) );
  nand2_1 U14289 ( .ip1(n12507), .ip2(n12485), .op(n12486) );
  nand3_1 U14290 ( .ip1(n12487), .ip2(n1485), .ip3(n12486), .op(n6054) );
  nand2_1 U14291 ( .ip1(n12510), .ip2(\CORTEXM0DS_INST/u_logic/D1fvx4 ), .op(
        n12491) );
  nand2_1 U14292 ( .ip1(n12497), .ip2(n12495), .op(n12488) );
  nand2_1 U14293 ( .ip1(\CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/D1fvx4 ), .op(n12496) );
  xor2_1 U14294 ( .ip1(n12488), .ip2(n12496), .op(n12489) );
  nand2_1 U14295 ( .ip1(n12507), .ip2(n12489), .op(n12490) );
  nand3_1 U14296 ( .ip1(n12491), .ip2(n1482), .ip3(n12490), .op(n6053) );
  nand2_1 U14297 ( .ip1(n12510), .ip2(\CORTEXM0DS_INST/u_logic/O2fvx4 ), .op(
        n12494) );
  nand3_1 U14298 ( .ip1(n12497), .ip2(n12495), .ip3(n12496), .op(n12502) );
  nand2_1 U14299 ( .ip1(\CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/O2fvx4 ), .op(n12504) );
  xor2_1 U14300 ( .ip1(n12502), .ip2(n12504), .op(n12492) );
  nand2_1 U14301 ( .ip1(n12507), .ip2(n12492), .op(n12493) );
  nand3_1 U14302 ( .ip1(n12494), .ip2(n1479), .ip3(n12493), .op(n6052) );
  nand2_1 U14303 ( .ip1(n12510), .ip2(\CORTEXM0DS_INST/u_logic/Z3fvx4 ), .op(
        n12501) );
  nand4_1 U14304 ( .ip1(n12497), .ip2(n12496), .ip3(n12495), .ip4(n12504), 
        .op(n12498) );
  nand2_1 U14305 ( .ip1(\CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Z3fvx4 ), .op(n12503) );
  xor2_1 U14306 ( .ip1(n12498), .ip2(n12503), .op(n12499) );
  nand2_1 U14307 ( .ip1(n12507), .ip2(n12499), .op(n12500) );
  nand3_1 U14308 ( .ip1(n12501), .ip2(n1476), .ip3(n12500), .op(n6051) );
  nand2_1 U14309 ( .ip1(n12510), .ip2(\CORTEXM0DS_INST/u_logic/K5fvx4 ), .op(
        n12509) );
  inv_1 U14310 ( .ip(n12502), .op(n12505) );
  nand3_1 U14311 ( .ip1(n12505), .ip2(n12504), .ip3(n12503), .op(n12506) );
  nand4_1 U14312 ( .ip1(\CORTEXM0DS_INST/u_logic/K5fvx4 ), .ip2(
        \CORTEXM0DS_INST/u_logic/Xlevx4 ), .ip3(n12507), .ip4(n12506), .op(
        n12508) );
  nand3_1 U14313 ( .ip1(n12509), .ip2(n1473), .ip3(n12508), .op(n6050) );
  nand2_1 U14314 ( .ip1(n12510), .ip2(\CORTEXM0DS_INST/u_logic/V6fvx4 ), .op(
        n12511) );
  nand2_1 U14315 ( .ip1(n1403), .ip2(n12511), .op(n6049) );
  nand2_1 U14316 ( .ip1(n1186), .ip2(\CORTEXM0DS_INST/u_logic/Cbfvx4 ), .op(
        n12512) );
  nand2_1 U14317 ( .ip1(n1188), .ip2(n12512), .op(n6047) );
  nand2_1 U14318 ( .ip1(n1186), .ip2(\CORTEXM0DS_INST/u_logic/Mcfvx4 ), .op(
        n12513) );
  nand2_1 U14319 ( .ip1(n1184), .ip2(n12513), .op(n6046) );
  nand2_1 U14320 ( .ip1(n1186), .ip2(\CORTEXM0DS_INST/u_logic/Wdfvx4 ), .op(
        n12514) );
  nand2_1 U14321 ( .ip1(n1182), .ip2(n12514), .op(n6045) );
  nand2_1 U14322 ( .ip1(n1186), .ip2(\CORTEXM0DS_INST/u_logic/Gffvx4 ), .op(
        n12515) );
  nand2_1 U14323 ( .ip1(n1180), .ip2(n12515), .op(n6044) );
  nand2_1 U14324 ( .ip1(n1186), .ip2(\CORTEXM0DS_INST/u_logic/Qgfvx4 ), .op(
        n12516) );
  nand2_1 U14325 ( .ip1(n1178), .ip2(n12516), .op(n6043) );
  nand2_1 U14326 ( .ip1(n1186), .ip2(\CORTEXM0DS_INST/u_logic/Aifvx4 ), .op(
        n12517) );
  nand2_1 U14327 ( .ip1(n1176), .ip2(n12517), .op(n6042) );
  nand2_1 U14328 ( .ip1(n1186), .ip2(\CORTEXM0DS_INST/u_logic/Kjfvx4 ), .op(
        n12518) );
  nand2_1 U14329 ( .ip1(n1174), .ip2(n12518), .op(n6041) );
  nand2_1 U14330 ( .ip1(n1186), .ip2(\CORTEXM0DS_INST/u_logic/Ukfvx4 ), .op(
        n12519) );
  nand2_1 U14331 ( .ip1(n1172), .ip2(n12519), .op(n6040) );
  nor2_1 U14332 ( .ip1(n1169), .ip2(n12527), .op(n12520) );
  mux2_1 U14333 ( .ip1(\CORTEXM0DS_INST/u_logic/Emfvx4 ), .ip2(n12520), .s(
        n12528), .op(n6039) );
  nand2_1 U14334 ( .ip1(n1186), .ip2(\CORTEXM0DS_INST/u_logic/Onfvx4 ), .op(
        n12521) );
  nand2_1 U14335 ( .ip1(n1168), .ip2(n12521), .op(n6038) );
  nand2_1 U14336 ( .ip1(n1186), .ip2(\CORTEXM0DS_INST/u_logic/Yofvx4 ), .op(
        n12522) );
  nand2_1 U14337 ( .ip1(n1166), .ip2(n12522), .op(n6037) );
  nand2_1 U14338 ( .ip1(n1186), .ip2(\CORTEXM0DS_INST/u_logic/Jqfvx4 ), .op(
        n12523) );
  nand2_1 U14339 ( .ip1(n1164), .ip2(n12523), .op(n6036) );
  nand2_1 U14340 ( .ip1(n1186), .ip2(\CORTEXM0DS_INST/u_logic/Urfvx4 ), .op(
        n12524) );
  nand2_1 U14341 ( .ip1(n1162), .ip2(n12524), .op(n6035) );
  nand2_1 U14342 ( .ip1(n1186), .ip2(\CORTEXM0DS_INST/u_logic/Ftfvx4 ), .op(
        n12525) );
  nand2_1 U14343 ( .ip1(n1160), .ip2(n12525), .op(n6034) );
  nor2_1 U14344 ( .ip1(n1157), .ip2(n12527), .op(n12526) );
  mux2_1 U14345 ( .ip1(\CORTEXM0DS_INST/u_logic/Qufvx4 ), .ip2(n12526), .s(
        n12528), .op(n6033) );
  nor2_1 U14346 ( .ip1(n1155), .ip2(n12527), .op(n12529) );
  mux2_1 U14347 ( .ip1(\CORTEXM0DS_INST/u_logic/Bwfvx4 ), .ip2(n12529), .s(
        n12528), .op(n6032) );
  and2_1 U14348 ( .ip1(\CORTEXM0DS_INST/u_logic/K5fvx4 ), .ip2(n12594), .op(
        n12532) );
  nor2_1 U14349 ( .ip1(n12593), .ip2(n12530), .op(n12531) );
  not_ab_or_c_or_d U14350 ( .ip1(n12597), .ip2(
        \CORTEXM0DS_INST/u_logic/Ftfvx4 ), .ip3(n12532), .ip4(n12531), .op(
        n12533) );
  nand3_1 U14351 ( .ip1(n1147), .ip2(n1145), .ip3(n12533), .op(n6030) );
  nor2_1 U14352 ( .ip1(n12534), .ip2(n12568), .op(n12537) );
  nor2_1 U14353 ( .ip1(n12593), .ip2(n12535), .op(n12536) );
  not_ab_or_c_or_d U14354 ( .ip1(n12597), .ip2(
        \CORTEXM0DS_INST/u_logic/Cbfvx4 ), .ip3(n12537), .ip4(n12536), .op(
        n12538) );
  nand3_1 U14355 ( .ip1(n1141), .ip2(n1139), .ip3(n12538), .op(n6029) );
  nor2_1 U14356 ( .ip1(n12539), .ip2(n12568), .op(n12542) );
  nor2_1 U14357 ( .ip1(n12593), .ip2(n12540), .op(n12541) );
  not_ab_or_c_or_d U14358 ( .ip1(n12597), .ip2(
        \CORTEXM0DS_INST/u_logic/Mcfvx4 ), .ip3(n12542), .ip4(n12541), .op(
        n12543) );
  nand3_1 U14359 ( .ip1(n1136), .ip2(n1134), .ip3(n12543), .op(n6028) );
  nor2_1 U14360 ( .ip1(n12593), .ip2(n12544), .op(n12547) );
  nor2_1 U14361 ( .ip1(n12545), .ip2(n12568), .op(n12546) );
  not_ab_or_c_or_d U14362 ( .ip1(n12597), .ip2(
        \CORTEXM0DS_INST/u_logic/Wdfvx4 ), .ip3(n12547), .ip4(n12546), .op(
        n12548) );
  nand3_1 U14363 ( .ip1(n1131), .ip2(n1129), .ip3(n12548), .op(n6027) );
  nor2_1 U14364 ( .ip1(n12549), .ip2(n12568), .op(n12552) );
  nor2_1 U14365 ( .ip1(n12593), .ip2(n12550), .op(n12551) );
  not_ab_or_c_or_d U14366 ( .ip1(n12597), .ip2(
        \CORTEXM0DS_INST/u_logic/Gffvx4 ), .ip3(n12552), .ip4(n12551), .op(
        n12553) );
  nand3_1 U14367 ( .ip1(n1126), .ip2(n1124), .ip3(n12553), .op(n6026) );
  nor2_1 U14368 ( .ip1(n12593), .ip2(n12554), .op(n12556) );
  and2_1 U14369 ( .ip1(\CORTEXM0DS_INST/u_logic/Vsevx4 ), .ip2(n12594), .op(
        n12555) );
  not_ab_or_c_or_d U14370 ( .ip1(n12597), .ip2(
        \CORTEXM0DS_INST/u_logic/Qgfvx4 ), .ip3(n12556), .ip4(n12555), .op(
        n12557) );
  nand3_1 U14371 ( .ip1(n1121), .ip2(n1119), .ip3(n12557), .op(n6025) );
  nor2_1 U14372 ( .ip1(n12593), .ip2(n12558), .op(n12561) );
  nor2_1 U14373 ( .ip1(n12559), .ip2(n12568), .op(n12560) );
  not_ab_or_c_or_d U14374 ( .ip1(n12597), .ip2(
        \CORTEXM0DS_INST/u_logic/Aifvx4 ), .ip3(n12561), .ip4(n12560), .op(
        n12562) );
  nand3_1 U14375 ( .ip1(n1116), .ip2(n1114), .ip3(n12562), .op(n6024) );
  nor2_1 U14376 ( .ip1(n12563), .ip2(n12568), .op(n12566) );
  nor2_1 U14377 ( .ip1(n12593), .ip2(n12564), .op(n12565) );
  not_ab_or_c_or_d U14378 ( .ip1(n12597), .ip2(
        \CORTEXM0DS_INST/u_logic/Kjfvx4 ), .ip3(n12566), .ip4(n12565), .op(
        n12567) );
  nand3_1 U14379 ( .ip1(n1111), .ip2(n1109), .ip3(n12567), .op(n6023) );
  nor2_1 U14380 ( .ip1(n12569), .ip2(n12568), .op(n12572) );
  nor2_1 U14381 ( .ip1(n12593), .ip2(n12570), .op(n12571) );
  not_ab_or_c_or_d U14382 ( .ip1(n12597), .ip2(
        \CORTEXM0DS_INST/u_logic/Ukfvx4 ), .ip3(n12572), .ip4(n12571), .op(
        n12573) );
  nand3_1 U14383 ( .ip1(n1106), .ip2(n1104), .ip3(n12573), .op(n6022) );
  nand2_1 U14384 ( .ip1(\CORTEXM0DS_INST/u_logic/Y99vx4 ), .ip2(n12574), .op(
        n12579) );
  and2_1 U14385 ( .ip1(\CORTEXM0DS_INST/u_logic/Jyevx4 ), .ip2(n12594), .op(
        n12577) );
  nor2_1 U14386 ( .ip1(n1169), .ip2(n12575), .op(n12576) );
  not_ab_or_c_or_d U14387 ( .ip1(\CORTEXM0DS_INST/u_logic/Emfvx4 ), .ip2(
        n12597), .ip3(n12577), .ip4(n12576), .op(n12578) );
  nand3_1 U14388 ( .ip1(n12579), .ip2(n12578), .ip3(n1101), .op(n6021) );
  and2_1 U14389 ( .ip1(\CORTEXM0DS_INST/u_logic/Tzevx4 ), .ip2(n12594), .op(
        n12582) );
  nor2_1 U14390 ( .ip1(n12593), .ip2(n12580), .op(n12581) );
  not_ab_or_c_or_d U14391 ( .ip1(n12597), .ip2(
        \CORTEXM0DS_INST/u_logic/Onfvx4 ), .ip3(n12582), .ip4(n12581), .op(
        n12583) );
  nand3_1 U14392 ( .ip1(n1096), .ip2(n1094), .ip3(n12583), .op(n6020) );
  nor2_1 U14393 ( .ip1(n12593), .ip2(n12584), .op(n12586) );
  and2_1 U14394 ( .ip1(\CORTEXM0DS_INST/u_logic/D1fvx4 ), .ip2(n12594), .op(
        n12585) );
  not_ab_or_c_or_d U14395 ( .ip1(n12597), .ip2(
        \CORTEXM0DS_INST/u_logic/Yofvx4 ), .ip3(n12586), .ip4(n12585), .op(
        n12587) );
  nand3_1 U14396 ( .ip1(n1091), .ip2(n1089), .ip3(n12587), .op(n6019) );
  and2_1 U14397 ( .ip1(\CORTEXM0DS_INST/u_logic/O2fvx4 ), .ip2(n12594), .op(
        n12590) );
  nor2_1 U14398 ( .ip1(n12593), .ip2(n12588), .op(n12589) );
  not_ab_or_c_or_d U14399 ( .ip1(n12597), .ip2(
        \CORTEXM0DS_INST/u_logic/Jqfvx4 ), .ip3(n12590), .ip4(n12589), .op(
        n12591) );
  nand3_1 U14400 ( .ip1(n1086), .ip2(n1084), .ip3(n12591), .op(n6018) );
  nor2_1 U14401 ( .ip1(n12593), .ip2(n12592), .op(n12596) );
  and2_1 U14402 ( .ip1(\CORTEXM0DS_INST/u_logic/Z3fvx4 ), .ip2(n12594), .op(
        n12595) );
  not_ab_or_c_or_d U14403 ( .ip1(n12597), .ip2(
        \CORTEXM0DS_INST/u_logic/Urfvx4 ), .ip3(n12596), .ip4(n12595), .op(
        n12598) );
  nand3_1 U14404 ( .ip1(n1081), .ip2(n1079), .ip3(n12598), .op(n6017) );
  or3_1 U14405 ( .ip1(n4585), .ip2(n12600), .ip3(n12599), .op(n12601) );
  nand2_1 U14406 ( .ip1(n1063), .ip2(n12601), .op(n6015) );
  nor2_1 U14407 ( .ip1(\CORTEXM0DS_INST/u_logic/Dmgvx4 ), .ip2(n12602), .op(
        n1061) );
  nor2_1 U14408 ( .ip1(\CORTEXM0DS_INST/u_logic/Dbgvx4 ), .ip2(n12615), .op(
        n12611) );
  nor2_1 U14409 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n12603), .op(
        n12604) );
  not_ab_or_c_or_d U14410 ( .ip1(n12607), .ip2(n12606), .ip3(n12605), .ip4(
        n12604), .op(n12609) );
  nor2_1 U14411 ( .ip1(n12609), .ip2(n12608), .op(n12610) );
  nor2_1 U14412 ( .ip1(n12611), .ip2(n12610), .op(n12612) );
  nor2_1 U14413 ( .ip1(n12613), .ip2(n12612), .op(n12634) );
  nor3_1 U14414 ( .ip1(\CORTEXM0DS_INST/u_logic/U9gvx4 ), .ip2(n12615), .ip3(
        n12614), .op(n12624) );
  nor2_1 U14415 ( .ip1(\CORTEXM0DS_INST/u_logic/Vdgvx4 ), .ip2(n12616), .op(
        n12620) );
  nor2_1 U14416 ( .ip1(n12618), .ip2(n12617), .op(n12619) );
  nor2_1 U14417 ( .ip1(n12620), .ip2(n12619), .op(n12622) );
  nor2_1 U14418 ( .ip1(n12622), .ip2(n12621), .op(n12623) );
  not_ab_or_c_or_d U14419 ( .ip1(n12626), .ip2(n12625), .ip3(n12624), .ip4(
        n12623), .op(n12632) );
  nand2_1 U14420 ( .ip1(n12628), .ip2(n12627), .op(n12629) );
  nand4_1 U14421 ( .ip1(n12632), .ip2(n12631), .ip3(n12630), .ip4(n12629), 
        .op(n12633) );
  nor2_1 U14422 ( .ip1(n12634), .ip2(n12633), .op(n1062) );
  nor2_1 U14423 ( .ip1(n12636), .ip2(n12635), .op(n489) );
  mux2_1 U14424 ( .ip1(\CORTEXM0DS_INST/u_logic/Uth2z4 [1]), .ip2(n12638), .s(
        n489), .op(n6014) );
  nand2_1 U14425 ( .ip1(n12637), .ip2(\CORTEXM0DS_INST/u_logic/Mf8vx4 ), .op(
        n488) );
  mux2_1 U14426 ( .ip1(n12638), .ip2(\CORTEXM0DS_INST/u_logic/Txh2z4 [1]), .s(
        n488), .op(n6013) );
  mux2_1 U14427 ( .ip1(\CORTEXM0DS_INST/u_logic/Czh2z4 [23]), .ip2(n4711), .s(
        n12695), .op(n6012) );
  mux2_1 U14428 ( .ip1(n4711), .ip2(\CORTEXM0DS_INST/u_logic/Psh2z4 [1]), .s(
        n488), .op(n6011) );
  nor2_1 U14429 ( .ip1(\CORTEXM0DS_INST/u_logic/I4gvx4 ), .ip2(n12639), .op(
        n12640) );
  nor2_1 U14430 ( .ip1(n12641), .ip2(n12640), .op(n12643) );
  mux2_1 U14431 ( .ip1(\CORTEXM0DS_INST/u_logic/A3gvx4 ), .ip2(n12643), .s(
        n12642), .op(n6010) );
  mux2_1 U14432 ( .ip1(\CORTEXM0DS_INST/u_logic/Q5gvx4 ), .ip2(n12644), .s(
        n12645), .op(n6009) );
  mux2_1 U14433 ( .ip1(n12647), .ip2(n12646), .s(n12645), .op(n12648) );
  inv_1 U14434 ( .ip(n12648), .op(n6008) );
  nor3_1 U14435 ( .ip1(n12651), .ip2(n12650), .ip3(n12649), .op(n12655) );
  nor3_1 U14436 ( .ip1(\CORTEXM0DS_INST/u_logic/Mj8vx4 ), .ip2(n12653), .ip3(
        n12652), .op(n12654) );
  or2_1 U14437 ( .ip1(n12655), .ip2(n12654), .op(n12656) );
  mux2_1 U14438 ( .ip1(n12656), .ip2(\CORTEXM0DS_INST/u_logic/Hx8vx4 ), .s(
        n5938), .op(n6007) );
  mux2_1 U14439 ( .ip1(n12657), .ip2(\CORTEXM0DS_INST/u_logic/Mxfvx4 ), .s(
        n1186), .op(n6005) );
  nand2_1 U14440 ( .ip1(n12658), .ip2(n12664), .op(n6003) );
  nand2_1 U14441 ( .ip1(n12659), .ip2(n12664), .op(n6001) );
  nand2_1 U14442 ( .ip1(n12660), .ip2(n12664), .op(n5999) );
  nand2_1 U14443 ( .ip1(n12661), .ip2(n12664), .op(n5997) );
  nand2_1 U14444 ( .ip1(n12662), .ip2(n12664), .op(n5995) );
  nand2_1 U14445 ( .ip1(n12663), .ip2(n12664), .op(n5993) );
  nand2_1 U14446 ( .ip1(n12665), .ip2(n12664), .op(n5991) );
  or2_1 U14447 ( .ip1(n12680), .ip2(n12666), .op(n5989) );
  nand2_1 U14448 ( .ip1(n12667), .ip2(n12680), .op(n5990) );
  nand2_1 U14449 ( .ip1(n12679), .ip2(n12668), .op(n5987) );
  nand2_1 U14450 ( .ip1(n12669), .ip2(n12680), .op(n5988) );
  nand2_1 U14451 ( .ip1(n12679), .ip2(n12670), .op(n5985) );
  nand2_1 U14452 ( .ip1(n12671), .ip2(n12680), .op(n5986) );
  nand2_1 U14453 ( .ip1(n12679), .ip2(n12672), .op(n5983) );
  nand2_1 U14454 ( .ip1(n12673), .ip2(n12680), .op(n5984) );
  nand2_1 U14455 ( .ip1(n12679), .ip2(n12674), .op(n5981) );
  nand2_1 U14456 ( .ip1(n12675), .ip2(n12680), .op(n5982) );
  nand2_1 U14457 ( .ip1(n12679), .ip2(n12676), .op(n5979) );
  nand2_1 U14458 ( .ip1(n12677), .ip2(n12680), .op(n5980) );
  nand2_1 U14459 ( .ip1(n12679), .ip2(n12678), .op(n5977) );
  nand2_1 U14460 ( .ip1(n12681), .ip2(n12680), .op(n5978) );
  and3_1 U14461 ( .ip1(n12683), .ip2(n12682), .ip3(
        \CORTEXM0DS_INST/u_logic/Mf8vx4 ), .op(n2) );
  nor2_1 U14462 ( .ip1(n12685), .ip2(n12684), .op(n1) );
  nor4_1 U14464 ( .ip1(PID_haddr_top[15]), .ip2(PID_haddr_top[16]), .ip3(n6117), .ip4(n5915), .op(n5932) );
  nor4_1 U14465 ( .ip1(PID_haddr_top[31]), .ip2(PID_haddr_top[28]), .ip3(
        PID_haddr_top[25]), .ip4(n2214), .op(n2215) );
  nor4_1 U14466 ( .ip1(PID_haddr_top[29]), .ip2(PID_haddr_top[30]), .ip3(
        PID_haddr_top[24]), .ip4(PID_haddr_top[22]), .op(n2216) );
  nand4_1 U14467 ( .ip1(HREADY_top), .ip2(PID_haddr_top[13]), .ip3(n5932), 
        .ip4(PID_haddr_top[12]), .op(n5931) );
  nor4_1 U14468 ( .ip1(PID_haddr_top[28]), .ip2(n2208), .ip3(n4585), .ip4(
        n2209), .op(n3127) );
  nand4_1 U14469 ( .ip1(PID_haddr_top[13]), .ip2(n2213), .ip3(
        PID_haddr_top[14]), .ip4(n1676), .op(n1678) );
  nor4_1 U14470 ( .ip1(PID_haddr_top[20]), .ip2(PID_haddr_top[19]), .ip3(
        PID_haddr_top[21]), .ip4(PID_haddr_top[18]), .op(n2217) );
  nand4_1 U14471 ( .ip1(\CORTEXM0DS_INST/u_logic/Cqovx4 ), .ip2(n2217), .ip3(
        PID_haddr_top[15]), .ip4(PID_hsize_top[1]), .op(n1677) );
  nor4_1 U14472 ( .ip1(PID_haddr_top[5]), .ip2(PID_haddr_top[10]), .ip3(
        PID_haddr_top[6]), .ip4(PID_haddr_top[11]), .op(n1668) );
  nor4_1 U14473 ( .ip1(PID_hwdata_top[16]), .ip2(PID_hwdata_top[28]), .ip3(
        PID_hwdata_top[24]), .ip4(PID_hwdata_top[17]), .op(n3228) );
  nor4_1 U14474 ( .ip1(PID_hwdata_top[20]), .ip2(PID_hwdata_top[21]), .ip3(
        n3231), .ip4(n3230), .op(n3233) );
  nor4_1 U14475 ( .ip1(PID_hwdata_top[26]), .ip2(PID_hwdata_top[22]), .ip3(
        PID_hwdata_top[18]), .ip4(PID_hwdata_top[19]), .op(n3229) );
  nand4_1 U14476 ( .ip1(PID_hwdata_top[2]), .ip2(PID_hwdata_top[21]), .ip3(
        PID_hwdata_top[20]), .ip4(n3227), .op(n2270) );
  nand4_1 U14477 ( .ip1(HREADY_top), .ip2(n5022), .ip3(n5100), .ip4(n5021), 
        .op(n5428) );
  nor2_1 U14478 ( .ip1(PID_hwdata_top[11]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [11]), .op(n12740) );
  nor2_1 U14479 ( .ip1(PID_hwdata_top[9]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [9]), .op(n12741) );
  nor2_1 U14480 ( .ip1(PID_hwdata_top[10]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [10]), .op(n12742) );
  nor2_1 U14481 ( .ip1(PID_hwdata_top[13]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [13]), .op(n12743) );
  nor2_1 U14482 ( .ip1(PID_hwdata_top[15]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [15]), .op(n12744) );
  nor2_1 U14483 ( .ip1(PID_hwdata_top[8]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [8]), .op(n12745) );
  nor2_1 U14484 ( .ip1(PID_hwdata_top[12]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [12]), .op(n12746) );
  nor2_1 U14485 ( .ip1(PID_hwdata_top[0]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [0]), .op(n12747) );
  nor2_1 U14486 ( .ip1(PID_hwdata_top[3]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [3]), .op(n12748) );
  nor2_1 U14487 ( .ip1(PID_hwdata_top[6]), .ip2(
        \CORTEXM0DS_INST/u_logic/T1i2z4 [6]), .op(n12749) );
  nor2_1 U14488 ( .ip1(PID_hwdata_top[26]), .ip2(n2326), .op(n12750) );
  nor2_1 U14489 ( .ip1(PID_hwdata_top[7]), .ip2(n3223), .op(n12751) );
endmodule

