
module i_i2c_DW_apb_i2c_regfile ( pclk, presetn, wr_en, rd_en, byte_en, 
        reg_addr, ipwdata, iprdata, ic_clr_intr_en, ic_clr_rx_under_en, 
        ic_clr_rx_over_en, ic_clr_tx_over_en, ic_clr_rd_req_en, 
        ic_clr_tx_abrt_en, ic_clr_rx_done_en, ic_clr_activity_en, 
        ic_clr_stop_det_en, ic_clr_start_det_en, ic_clr_gen_call_en, 
        mst_activity, slv_activity, activity, ic_tx_abrt_source, ic_en, 
        slv_rx_aborted_sync, slv_fifo_filled_and_flushed_sync, ic_tar, ic_sar, 
        ic_hs_maddr, ic_fs_hcnt, ic_fs_lcnt, ic_intr_mask, ic_rx_tl_int, 
        ic_enable, ic_hcnt, ic_lcnt, ic_fs_spklen, ic_hs_spklen, ic_intr_stat, 
        ic_raw_intr_stat, ic_hs, ic_fs, ic_ss, ic_master, ic_10bit_mst, 
        ic_10bit_slv, ic_slave_en, p_det_ifaddr, tx_empty_ctrl, rx_pop_data, 
        tx_push_data, fifo_rst_n, tx_fifo_rst_n, tx_pop_sync, rx_push_sync, 
        rx_pop, tx_push, tx_empty, rx_full, tx_full, rx_empty, tx_abrt_flg_edg, 
        abrt_in_rcve_trns, slv_clr_leftover_flg_edg, ic_rstrt_en, ic_sda_setup, 
        ic_sda_hold, ic_ack_general_call, ic_tx_tl_7_, ic_tx_tl_6_, 
        ic_tx_tl_5_, ic_tx_tl_4_, ic_tx_tl_3__BAR, ic_tx_tl_2_, ic_tx_tl_1_, 
        ic_tx_tl_0_ );
  input [3:0] byte_en;
  input [5:0] reg_addr;
  input [31:0] ipwdata;
  output [31:0] iprdata;
  input [16:0] ic_tx_abrt_source;
  output [11:0] ic_tar;
  output [9:0] ic_sar;
  output [2:0] ic_hs_maddr;
  output [15:0] ic_fs_hcnt;
  output [15:0] ic_fs_lcnt;
  output [13:0] ic_intr_mask;
  output [2:0] ic_rx_tl_int;
  output [1:0] ic_enable;
  output [15:0] ic_hcnt;
  output [15:0] ic_lcnt;
  output [7:0] ic_fs_spklen;
  output [7:0] ic_hs_spklen;
  input [13:0] ic_intr_stat;
  input [13:0] ic_raw_intr_stat;
  input [7:0] rx_pop_data;
  output [8:0] tx_push_data;
  output [7:0] ic_sda_setup;
  output [23:0] ic_sda_hold;
  input pclk, presetn, wr_en, rd_en, mst_activity, slv_activity, activity,
         ic_en, slv_rx_aborted_sync, slv_fifo_filled_and_flushed_sync,
         tx_pop_sync, rx_push_sync, tx_empty, rx_full, tx_full, rx_empty,
         tx_abrt_flg_edg, abrt_in_rcve_trns, slv_clr_leftover_flg_edg;
  output ic_clr_intr_en, ic_clr_rx_under_en, ic_clr_rx_over_en,
         ic_clr_tx_over_en, ic_clr_rd_req_en, ic_clr_tx_abrt_en,
         ic_clr_rx_done_en, ic_clr_activity_en, ic_clr_stop_det_en,
         ic_clr_start_det_en, ic_clr_gen_call_en, ic_hs, ic_fs, ic_ss,
         ic_master, ic_10bit_mst, ic_10bit_slv, ic_slave_en, p_det_ifaddr,
         tx_empty_ctrl, fifo_rst_n, tx_fifo_rst_n, rx_pop, tx_push,
         ic_rstrt_en, ic_ack_general_call, ic_tx_tl_7_, ic_tx_tl_6_,
         ic_tx_tl_5_, ic_tx_tl_4_, ic_tx_tl_3__BAR, ic_tx_tl_2_, ic_tx_tl_1_,
         ic_tx_tl_0_;
  wire   activity_r, mst_activity_r, slv_activity_r, ic_con_pre_6_,
         ic_con_pre_2_, ic_con_pre_1_, fifo_rst_n_int, fix_c, n1105, n1107,
         n1109, n1111, n1113, n1115, n1117, n1119, n1121, n1123, n1125, n1127,
         n1129, n1131, n1133, n1135, n1137, n1149, n1151, n1153, n1165, n1167,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n761;
  wire   [3:0] ic_txflr;
  wire   [3:0] ic_txflr_flushed;
  wire   [3:0] ic_rxflr;
  wire   [15:0] hcr_ic_ss_hcnt;
  wire   [15:0] hcr_ic_ss_lcnt;
  wire   [15:0] hcr_ic_hs_hcnt;
  wire   [15:0] hcr_ic_hs_lcnt;

  drp_1 mst_activity_r_reg ( .ip(mst_activity), .ck(pclk), .rb(presetn), .q(
        mst_activity_r) );
  drp_1 slv_activity_r_reg ( .ip(slv_activity), .ck(pclk), .rb(presetn), .q(
        slv_activity_r) );
  drp_1 activity_r_reg ( .ip(activity), .ck(pclk), .rb(presetn), .q(activity_r) );
  drp_1 ic_enable_reg_reg_0_ ( .ip(n1549), .ck(pclk), .rb(presetn), .q(
        ic_enable[0]) );
  drp_1 ic_enable_reg_reg_1_ ( .ip(n1548), .ck(pclk), .rb(presetn), .q(
        ic_enable[1]) );
  drp_1 ic_rxflr_reg_0_ ( .ip(n1546), .ck(pclk), .rb(presetn), .q(ic_rxflr[0])
         );
  drp_1 ic_rxflr_reg_2_ ( .ip(n1544), .ck(pclk), .rb(presetn), .q(ic_rxflr[2])
         );
  drp_1 ic_rxflr_reg_3_ ( .ip(n1547), .ck(pclk), .rb(presetn), .q(ic_rxflr[3])
         );
  drp_1 ic_rxflr_reg_1_ ( .ip(n1545), .ck(pclk), .rb(presetn), .q(ic_rxflr[1])
         );
  drp_1 ic_con_pre_reg_8_ ( .ip(n1543), .ck(pclk), .rb(presetn), .q(
        tx_empty_ctrl) );
  drp_1 ic_con_pre_reg_7_ ( .ip(n1542), .ck(pclk), .rb(presetn), .q(
        p_det_ifaddr) );
  drp_1 ic_tar_reg_reg_11_ ( .ip(n1529), .ck(pclk), .rb(presetn), .q(
        ic_tar[11]) );
  drp_1 ic_tar_reg_reg_10_ ( .ip(n1530), .ck(pclk), .rb(presetn), .q(
        ic_tar[10]) );
  drp_1 ic_tar_reg_reg_9_ ( .ip(n1531), .ck(pclk), .rb(presetn), .q(ic_tar[9])
         );
  drp_1 ic_tar_reg_reg_8_ ( .ip(n1532), .ck(pclk), .rb(presetn), .q(ic_tar[8])
         );
  drp_1 ic_tar_reg_reg_7_ ( .ip(n1513), .ck(pclk), .rb(presetn), .q(ic_tar[7])
         );
  drp_1 ic_tar_reg_reg_5_ ( .ip(n1515), .ck(pclk), .rb(presetn), .q(ic_tar[5])
         );
  drp_1 ic_tar_reg_reg_3_ ( .ip(n1517), .ck(pclk), .rb(presetn), .q(ic_tar[3])
         );
  drp_1 ic_tar_reg_reg_1_ ( .ip(n1519), .ck(pclk), .rb(presetn), .q(ic_tar[1])
         );
  drp_1 ic_sar_reg_9_ ( .ip(n1533), .ck(pclk), .rb(presetn), .q(ic_sar[9]) );
  drp_1 ic_sar_reg_8_ ( .ip(n1534), .ck(pclk), .rb(presetn), .q(ic_sar[8]) );
  drp_1 ic_sar_reg_7_ ( .ip(n1521), .ck(pclk), .rb(presetn), .q(ic_sar[7]) );
  drp_1 ic_sar_reg_5_ ( .ip(n1523), .ck(pclk), .rb(presetn), .q(ic_sar[5]) );
  drp_1 ic_sar_reg_3_ ( .ip(n1525), .ck(pclk), .rb(presetn), .q(ic_sar[3]) );
  drp_1 ic_sar_reg_1_ ( .ip(n1527), .ck(pclk), .rb(presetn), .q(ic_sar[1]) );
  drp_1 r_ic_ss_hcnt_reg_15_ ( .ip(n1504), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[15]) );
  drp_1 r_ic_ss_hcnt_reg_14_ ( .ip(n1497), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[14]) );
  drp_1 r_ic_ss_hcnt_reg_13_ ( .ip(n1498), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[13]) );
  drp_1 r_ic_ss_hcnt_reg_12_ ( .ip(n1499), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[12]) );
  drp_1 r_ic_ss_hcnt_reg_11_ ( .ip(n1500), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[11]) );
  drp_1 r_ic_ss_hcnt_reg_10_ ( .ip(n1501), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[10]) );
  drp_1 r_ic_ss_hcnt_reg_9_ ( .ip(n1502), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[9]) );
  drp_1 r_ic_ss_hcnt_reg_6_ ( .ip(n1506), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[6]) );
  drp_1 r_ic_ss_hcnt_reg_5_ ( .ip(n1507), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[5]) );
  drp_1 r_ic_ss_hcnt_reg_3_ ( .ip(n1509), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[3]) );
  drp_1 r_ic_ss_hcnt_reg_2_ ( .ip(n1510), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[2]) );
  drp_1 r_ic_ss_hcnt_reg_1_ ( .ip(n1511), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[1]) );
  drp_1 r_ic_ss_hcnt_reg_0_ ( .ip(n1512), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_hcnt[0]) );
  drp_1 r_ic_ss_lcnt_reg_3_ ( .ip(n1493), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[3]) );
  drp_1 r_ic_ss_lcnt_reg_5_ ( .ip(n1491), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[5]) );
  drp_1 r_ic_ss_lcnt_reg_15_ ( .ip(n1488), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[15]) );
  drp_1 r_ic_ss_lcnt_reg_9_ ( .ip(n1486), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[9]) );
  drp_1 r_ic_ss_lcnt_reg_10_ ( .ip(n1485), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[10]) );
  drp_1 r_ic_ss_lcnt_reg_11_ ( .ip(n1484), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[11]) );
  drp_1 r_ic_ss_lcnt_reg_12_ ( .ip(n1483), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[12]) );
  drp_1 r_ic_ss_lcnt_reg_13_ ( .ip(n1482), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[13]) );
  drp_1 r_ic_ss_lcnt_reg_14_ ( .ip(n1481), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[14]) );
  drp_1 r_ic_ss_lcnt_reg_0_ ( .ip(n1496), .ck(pclk), .rb(presetn), .q(
        hcr_ic_ss_lcnt[0]) );
  drp_1 r_ic_fs_hcnt_reg_15_ ( .ip(n1472), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[15]) );
  drp_1 r_ic_fs_hcnt_reg_14_ ( .ip(n1465), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[14]) );
  drp_1 r_ic_fs_hcnt_reg_13_ ( .ip(n1466), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[13]) );
  drp_1 r_ic_fs_hcnt_reg_12_ ( .ip(n1467), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[12]) );
  drp_1 r_ic_fs_hcnt_reg_11_ ( .ip(n1468), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[11]) );
  drp_1 r_ic_fs_hcnt_reg_10_ ( .ip(n1469), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[10]) );
  drp_1 r_ic_fs_hcnt_reg_9_ ( .ip(n1470), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[9]) );
  drp_1 r_ic_fs_hcnt_reg_8_ ( .ip(n1471), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[8]) );
  drp_1 r_ic_fs_hcnt_reg_7_ ( .ip(n1473), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[7]) );
  drp_1 r_ic_fs_hcnt_reg_6_ ( .ip(n1474), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[6]) );
  drp_1 r_ic_fs_hcnt_reg_1_ ( .ip(n1479), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[1]) );
  drp_1 r_ic_fs_hcnt_reg_0_ ( .ip(n1480), .ck(pclk), .rb(presetn), .q(
        ic_fs_hcnt[0]) );
  drp_1 r_ic_fs_lcnt_reg_3_ ( .ip(n1461), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[3]) );
  drp_1 r_ic_fs_lcnt_reg_4_ ( .ip(n1460), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[4]) );
  drp_1 r_ic_fs_lcnt_reg_5_ ( .ip(n1459), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[5]) );
  drp_1 r_ic_fs_lcnt_reg_6_ ( .ip(n1458), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[6]) );
  drp_1 r_ic_fs_lcnt_reg_15_ ( .ip(n1456), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[15]) );
  drp_1 r_ic_fs_lcnt_reg_8_ ( .ip(n1455), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[8]) );
  drp_1 r_ic_fs_lcnt_reg_9_ ( .ip(n1454), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[9]) );
  drp_1 r_ic_fs_lcnt_reg_10_ ( .ip(n1453), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[10]) );
  drp_1 r_ic_fs_lcnt_reg_11_ ( .ip(n1452), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[11]) );
  drp_1 r_ic_fs_lcnt_reg_12_ ( .ip(n1451), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[12]) );
  drp_1 r_ic_fs_lcnt_reg_13_ ( .ip(n1450), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[13]) );
  drp_1 r_ic_fs_lcnt_reg_14_ ( .ip(n1449), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[14]) );
  drp_1 r_ic_fs_lcnt_reg_2_ ( .ip(n1462), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[2]) );
  drp_1 r_ic_fs_lcnt_reg_0_ ( .ip(n1464), .ck(pclk), .rb(presetn), .q(
        ic_fs_lcnt[0]) );
  drp_1 r_ic_hs_hcnt_reg_15_ ( .ip(n1440), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[15]) );
  drp_1 r_ic_hs_hcnt_reg_14_ ( .ip(n1433), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[14]) );
  drp_1 r_ic_hs_hcnt_reg_13_ ( .ip(n1434), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[13]) );
  drp_1 r_ic_hs_hcnt_reg_12_ ( .ip(n1435), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[12]) );
  drp_1 r_ic_hs_hcnt_reg_11_ ( .ip(n1436), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[11]) );
  drp_1 r_ic_hs_hcnt_reg_10_ ( .ip(n1437), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[10]) );
  drp_1 r_ic_hs_hcnt_reg_9_ ( .ip(n1438), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[9]) );
  drp_1 r_ic_hs_hcnt_reg_8_ ( .ip(n1439), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[8]) );
  drp_1 r_ic_hs_hcnt_reg_7_ ( .ip(n1441), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[7]) );
  drp_1 r_ic_hs_hcnt_reg_6_ ( .ip(n1442), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[6]) );
  drp_1 r_ic_hs_hcnt_reg_5_ ( .ip(n1443), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[5]) );
  drp_1 r_ic_hs_hcnt_reg_4_ ( .ip(n1444), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[4]) );
  drp_1 r_ic_hs_hcnt_reg_3_ ( .ip(n1445), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[3]) );
  drp_1 r_ic_hs_hcnt_reg_0_ ( .ip(n1448), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_hcnt[0]) );
  drp_1 r_ic_hs_lcnt_reg_3_ ( .ip(n1429), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[3]) );
  drp_1 r_ic_hs_lcnt_reg_5_ ( .ip(n1427), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[5]) );
  drp_1 r_ic_hs_lcnt_reg_6_ ( .ip(n1426), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[6]) );
  drp_1 r_ic_hs_lcnt_reg_7_ ( .ip(n1425), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[7]) );
  drp_1 r_ic_hs_lcnt_reg_15_ ( .ip(n1424), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[15]) );
  drp_1 r_ic_hs_lcnt_reg_8_ ( .ip(n1423), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[8]) );
  drp_1 r_ic_hs_lcnt_reg_9_ ( .ip(n1422), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[9]) );
  drp_1 r_ic_hs_lcnt_reg_10_ ( .ip(n1421), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[10]) );
  drp_1 r_ic_hs_lcnt_reg_11_ ( .ip(n1420), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[11]) );
  drp_1 r_ic_hs_lcnt_reg_12_ ( .ip(n1419), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[12]) );
  drp_1 r_ic_hs_lcnt_reg_13_ ( .ip(n1418), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[13]) );
  drp_1 r_ic_hs_lcnt_reg_14_ ( .ip(n1417), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[14]) );
  drp_1 r_ic_hs_lcnt_reg_2_ ( .ip(n1430), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[2]) );
  drp_1 r_ic_hs_lcnt_reg_1_ ( .ip(n1431), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[1]) );
  drp_1 r_ic_hs_lcnt_reg_0_ ( .ip(n1432), .ck(pclk), .rb(presetn), .q(
        hcr_ic_hs_lcnt[0]) );
  drp_1 r_ic_fs_spklen_reg_7_ ( .ip(n1416), .ck(pclk), .rb(presetn), .q(
        ic_fs_spklen[7]) );
  drp_1 r_ic_fs_spklen_reg_6_ ( .ip(n1415), .ck(pclk), .rb(presetn), .q(
        ic_fs_spklen[6]) );
  drp_1 r_ic_fs_spklen_reg_5_ ( .ip(n1414), .ck(pclk), .rb(presetn), .q(
        ic_fs_spklen[5]) );
  drp_1 r_ic_fs_spklen_reg_4_ ( .ip(n1413), .ck(pclk), .rb(presetn), .q(
        ic_fs_spklen[4]) );
  drp_1 r_ic_fs_spklen_reg_3_ ( .ip(n1412), .ck(pclk), .rb(presetn), .q(
        ic_fs_spklen[3]) );
  drp_1 r_ic_fs_spklen_reg_1_ ( .ip(n1410), .ck(pclk), .rb(presetn), .q(
        ic_fs_spklen[1]) );
  drp_1 r_ic_hs_spklen_reg_7_ ( .ip(n1408), .ck(pclk), .rb(presetn), .q(
        ic_hs_spklen[7]) );
  drp_1 r_ic_hs_spklen_reg_6_ ( .ip(n1407), .ck(pclk), .rb(presetn), .q(
        ic_hs_spklen[6]) );
  drp_1 r_ic_hs_spklen_reg_5_ ( .ip(n1406), .ck(pclk), .rb(presetn), .q(
        ic_hs_spklen[5]) );
  drp_1 r_ic_hs_spklen_reg_4_ ( .ip(n1405), .ck(pclk), .rb(presetn), .q(
        ic_hs_spklen[4]) );
  drp_1 r_ic_hs_spklen_reg_3_ ( .ip(n1404), .ck(pclk), .rb(presetn), .q(
        ic_hs_spklen[3]) );
  drp_1 r_ic_hs_spklen_reg_2_ ( .ip(n1403), .ck(pclk), .rb(presetn), .q(
        ic_hs_spklen[2]) );
  drp_1 r_ic_hs_spklen_reg_1_ ( .ip(n1402), .ck(pclk), .rb(presetn), .q(
        ic_hs_spklen[1]) );
  drp_1 ic_intr_mask_reg_10_ ( .ip(n1398), .ck(pclk), .rb(presetn), .q(
        ic_intr_mask[10]) );
  drp_1 ic_intr_mask_reg_9_ ( .ip(n1399), .ck(pclk), .rb(presetn), .q(
        ic_intr_mask[9]) );
  drp_1 ic_intr_mask_reg_8_ ( .ip(n1400), .ck(pclk), .rb(presetn), .q(
        ic_intr_mask[8]) );
  drp_1 ic_sda_hold_reg_23_ ( .ip(n1388), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[23]) );
  drp_1 ic_sda_hold_reg_22_ ( .ip(n1387), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[22]) );
  drp_1 ic_sda_hold_reg_21_ ( .ip(n1386), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[21]) );
  drp_1 ic_sda_hold_reg_20_ ( .ip(n1385), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[20]) );
  drp_1 ic_sda_hold_reg_19_ ( .ip(n1384), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[19]) );
  drp_1 ic_sda_hold_reg_18_ ( .ip(n1383), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[18]) );
  drp_1 ic_sda_hold_reg_17_ ( .ip(n1382), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[17]) );
  drp_1 ic_sda_hold_reg_16_ ( .ip(n1381), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[16]) );
  drp_1 ic_sda_hold_reg_15_ ( .ip(n1380), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[15]) );
  drp_1 ic_sda_hold_reg_14_ ( .ip(n1379), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[14]) );
  drp_1 ic_sda_hold_reg_13_ ( .ip(n1378), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[13]) );
  drp_1 ic_sda_hold_reg_12_ ( .ip(n1377), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[12]) );
  drp_1 ic_sda_hold_reg_11_ ( .ip(n1376), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[11]) );
  drp_1 ic_sda_hold_reg_10_ ( .ip(n1375), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[10]) );
  drp_1 ic_sda_hold_reg_9_ ( .ip(n1374), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[9]) );
  drp_1 ic_sda_hold_reg_8_ ( .ip(n1373), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[8]) );
  drp_1 ic_sda_hold_reg_7_ ( .ip(n1372), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[7]) );
  drp_1 ic_sda_hold_reg_6_ ( .ip(n1371), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[6]) );
  drp_1 ic_sda_hold_reg_5_ ( .ip(n1370), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[5]) );
  drp_1 ic_sda_hold_reg_4_ ( .ip(n1369), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[4]) );
  drp_1 ic_sda_hold_reg_3_ ( .ip(n1368), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[3]) );
  drp_1 ic_sda_hold_reg_2_ ( .ip(n1367), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[2]) );
  drp_1 ic_sda_hold_reg_1_ ( .ip(n1366), .ck(pclk), .rb(presetn), .q(
        ic_sda_hold[1]) );
  drp_1 fifo_rst_n_int_reg ( .ip(fix_c), .ck(pclk), .rb(presetn), .q(
        fifo_rst_n_int) );
  drp_1 ic_txflr_reg_2_ ( .ip(n1361), .ck(pclk), .rb(presetn), .q(ic_txflr[2])
         );
  drp_1 ic_txflr_reg_3_ ( .ip(n1364), .ck(pclk), .rb(presetn), .q(ic_txflr[3])
         );
  drp_1 ic_txflr_reg_0_ ( .ip(n1363), .ck(pclk), .rb(presetn), .q(ic_txflr[0])
         );
  drp_1 ic_txflr_reg_1_ ( .ip(n1362), .ck(pclk), .rb(presetn), .q(ic_txflr[1])
         );
  drp_1 ic_hs_maddr_reg_2_ ( .ip(n1167), .ck(pclk), .rb(presetn), .q(
        ic_hs_maddr[2]) );
  drp_1 ic_hs_maddr_reg_1_ ( .ip(n1165), .ck(pclk), .rb(presetn), .q(
        ic_hs_maddr[1]) );
  drp_1 ic_rx_tl_reg_2_ ( .ip(n1153), .ck(pclk), .rb(presetn), .q(
        ic_rx_tl_int[2]) );
  drp_1 ic_rx_tl_reg_1_ ( .ip(n1151), .ck(pclk), .rb(presetn), .q(
        ic_rx_tl_int[1]) );
  drp_1 ic_rx_tl_reg_0_ ( .ip(n1149), .ck(pclk), .rb(presetn), .q(
        ic_rx_tl_int[0]) );
  drp_1 ic_tx_tl_reg_2_ ( .ip(n1137), .ck(pclk), .rb(presetn), .q(ic_tx_tl_2_)
         );
  drp_1 ic_tx_tl_reg_1_ ( .ip(n1135), .ck(pclk), .rb(presetn), .q(ic_tx_tl_1_)
         );
  drp_1 ic_tx_tl_reg_0_ ( .ip(n1133), .ck(pclk), .rb(presetn), .q(ic_tx_tl_0_)
         );
  drp_1 ic_sda_setup_reg_7_ ( .ip(n1131), .ck(pclk), .rb(presetn), .q(
        ic_sda_setup[7]) );
  drp_1 ic_sda_setup_reg_4_ ( .ip(n1129), .ck(pclk), .rb(presetn), .q(
        ic_sda_setup[4]) );
  drp_1 ic_sda_setup_reg_3_ ( .ip(n1127), .ck(pclk), .rb(presetn), .q(
        ic_sda_setup[3]) );
  drp_1 ic_sda_setup_reg_1_ ( .ip(n1125), .ck(pclk), .rb(presetn), .q(
        ic_sda_setup[1]) );
  drp_1 ic_sda_setup_reg_0_ ( .ip(n1123), .ck(pclk), .rb(presetn), .q(
        ic_sda_setup[0]) );
  drp_1 ic_txflr_flushed_reg_0_ ( .ip(n1121), .ck(pclk), .rb(presetn), .q(
        ic_txflr_flushed[0]) );
  drp_1 ic_txflr_flushed_reg_1_ ( .ip(n1119), .ck(pclk), .rb(presetn), .q(
        ic_txflr_flushed[1]) );
  drp_1 ic_txflr_flushed_reg_3_ ( .ip(n1117), .ck(pclk), .rb(presetn), .q(
        ic_txflr_flushed[3]) );
  drp_1 ic_txflr_flushed_reg_2_ ( .ip(n1115), .ck(pclk), .rb(presetn), .q(
        ic_txflr_flushed[2]) );
  drsp_1 ic_ack_general_call_reg ( .ip(n1105), .ck(pclk), .rb(1'b1), .s(n3), 
        .q(ic_ack_general_call) );
  drsp_1 ic_intr_mask_reg_4_ ( .ip(n1392), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_intr_mask[4]) );
  drsp_1 ic_intr_mask_reg_11_ ( .ip(n1397), .ck(pclk), .rb(1'b1), .s(n761), 
        .q(ic_intr_mask[11]) );
  drsp_1 ic_intr_mask_reg_3_ ( .ip(n1393), .ck(pclk), .rb(1'b1), .s(n4), .q(
        ic_intr_mask[3]) );
  drsp_1 ic_intr_mask_reg_6_ ( .ip(n1390), .ck(pclk), .rb(1'b1), .s(n3), .q(
        ic_intr_mask[6]) );
  drsp_1 ic_intr_mask_reg_1_ ( .ip(n1395), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_intr_mask[1]) );
  drsp_1 ic_intr_mask_reg_0_ ( .ip(n1396), .ck(pclk), .rb(1'b1), .s(n761), .q(
        ic_intr_mask[0]) );
  drsp_1 ic_intr_mask_reg_7_ ( .ip(n1389), .ck(pclk), .rb(1'b1), .s(n4), .q(
        ic_intr_mask[7]) );
  drsp_1 ic_intr_mask_reg_2_ ( .ip(n1394), .ck(pclk), .rb(1'b1), .s(n3), .q(
        ic_intr_mask[2]) );
  drsp_1 ic_intr_mask_reg_5_ ( .ip(n1391), .ck(pclk), .rb(1'b1), .s(n761), .q(
        ic_intr_mask[5]) );
  drsp_1 ic_hs_maddr_reg_0_ ( .ip(n1113), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_hs_maddr[0]) );
  drsp_1 r_ic_hs_spklen_reg_0_ ( .ip(n1401), .ck(pclk), .rb(1'b1), .s(n761), 
        .q(ic_hs_spklen[0]) );
  drsp_1 r_ic_fs_spklen_reg_0_ ( .ip(n1409), .ck(pclk), .rb(1'b1), .s(n4), .q(
        ic_fs_spklen[0]) );
  drsp_1 r_ic_fs_spklen_reg_2_ ( .ip(n1411), .ck(pclk), .rb(1'b1), .s(n3), .q(
        ic_fs_spklen[2]) );
  drsp_1 ic_sda_setup_reg_6_ ( .ip(n1111), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_sda_setup[6]) );
  drsp_1 ic_sda_setup_reg_2_ ( .ip(n1107), .ck(pclk), .rb(1'b1), .s(n761), .q(
        ic_sda_setup[2]) );
  drsp_1 ic_sda_setup_reg_5_ ( .ip(n1109), .ck(pclk), .rb(1'b1), .s(n4), .q(
        ic_sda_setup[5]) );
  drsp_1 ic_con_pre_reg_4_ ( .ip(n1539), .ck(pclk), .rb(1'b1), .s(n3), .q(
        ic_10bit_mst) );
  drsp_1 ic_con_pre_reg_2_ ( .ip(n1537), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_con_pre_2_) );
  drsp_1 ic_con_pre_reg_1_ ( .ip(n1536), .ck(pclk), .rb(1'b1), .s(n761), .q(
        ic_con_pre_1_) );
  drsp_1 ic_con_pre_reg_3_ ( .ip(n1538), .ck(pclk), .rb(1'b1), .s(n4), .q(
        ic_10bit_slv) );
  drsp_1 ic_con_pre_reg_6_ ( .ip(n1541), .ck(pclk), .rb(1'b1), .s(n3), .q(
        ic_con_pre_6_) );
  drsp_1 ic_con_pre_reg_0_ ( .ip(n1535), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_master) );
  drsp_1 ic_con_pre_reg_5_ ( .ip(n1540), .ck(pclk), .rb(1'b1), .s(n761), .q(
        ic_rstrt_en) );
  drsp_1 ic_sar_reg_4_ ( .ip(n1524), .ck(pclk), .rb(1'b1), .s(n4), .q(
        ic_sar[4]) );
  drsp_1 ic_sar_reg_6_ ( .ip(n1522), .ck(pclk), .rb(1'b1), .s(n3), .q(
        ic_sar[6]) );
  drsp_1 ic_sar_reg_0_ ( .ip(n1528), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_sar[0]) );
  drsp_1 ic_sar_reg_2_ ( .ip(n1526), .ck(pclk), .rb(1'b1), .s(n761), .q(
        ic_sar[2]) );
  drsp_1 r_ic_hs_hcnt_reg_2_ ( .ip(n1446), .ck(pclk), .rb(1'b1), .s(n4), .q(
        hcr_ic_hs_hcnt[2]) );
  drsp_1 r_ic_hs_hcnt_reg_1_ ( .ip(n1447), .ck(pclk), .rb(1'b1), .s(n3), .q(
        hcr_ic_hs_hcnt[1]) );
  drsp_1 r_ic_fs_hcnt_reg_2_ ( .ip(n1478), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_fs_hcnt[2]) );
  drsp_1 r_ic_fs_hcnt_reg_5_ ( .ip(n1475), .ck(pclk), .rb(1'b1), .s(n761), .q(
        ic_fs_hcnt[5]) );
  drsp_1 ic_tar_reg_reg_4_ ( .ip(n1516), .ck(pclk), .rb(1'b1), .s(n4), .q(
        ic_tar[4]) );
  drsp_1 ic_tar_reg_reg_6_ ( .ip(n1514), .ck(pclk), .rb(1'b1), .s(n3), .q(
        ic_tar[6]) );
  drsp_1 ic_tar_reg_reg_0_ ( .ip(n1520), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_tar[0]) );
  drsp_1 ic_tar_reg_reg_2_ ( .ip(n1518), .ck(pclk), .rb(1'b1), .s(n761), .q(
        ic_tar[2]) );
  drsp_1 r_ic_fs_lcnt_reg_7_ ( .ip(n1457), .ck(pclk), .rb(1'b1), .s(n4), .q(
        ic_fs_lcnt[7]) );
  drsp_1 r_ic_hs_lcnt_reg_4_ ( .ip(n1428), .ck(pclk), .rb(1'b1), .s(n3), .q(
        hcr_ic_hs_lcnt[4]) );
  drsp_1 r_ic_ss_lcnt_reg_8_ ( .ip(n1487), .ck(pclk), .rb(1'b1), .s(n2), .q(
        hcr_ic_ss_lcnt[8]) );
  drsp_1 r_ic_ss_lcnt_reg_6_ ( .ip(n1490), .ck(pclk), .rb(1'b1), .s(n761), .q(
        hcr_ic_ss_lcnt[6]) );
  drsp_1 r_ic_ss_lcnt_reg_4_ ( .ip(n1492), .ck(pclk), .rb(1'b1), .s(n4), .q(
        hcr_ic_ss_lcnt[4]) );
  drsp_1 r_ic_ss_lcnt_reg_2_ ( .ip(n1494), .ck(pclk), .rb(1'b1), .s(n3), .q(
        hcr_ic_ss_lcnt[2]) );
  drsp_1 r_ic_ss_lcnt_reg_1_ ( .ip(n1495), .ck(pclk), .rb(1'b1), .s(n2), .q(
        hcr_ic_ss_lcnt[1]) );
  drsp_1 r_ic_ss_lcnt_reg_7_ ( .ip(n1489), .ck(pclk), .rb(1'b1), .s(n761), .q(
        hcr_ic_ss_lcnt[7]) );
  drsp_1 r_ic_fs_lcnt_reg_1_ ( .ip(n1463), .ck(pclk), .rb(1'b1), .s(n4), .q(
        ic_fs_lcnt[1]) );
  drsp_1 ic_sda_hold_reg_0_ ( .ip(n1365), .ck(pclk), .rb(1'b1), .s(n3), .q(
        ic_sda_hold[0]) );
  drsp_1 r_ic_ss_hcnt_reg_8_ ( .ip(n1503), .ck(pclk), .rb(1'b1), .s(n2), .q(
        hcr_ic_ss_hcnt[8]) );
  drsp_1 r_ic_ss_hcnt_reg_4_ ( .ip(n1508), .ck(pclk), .rb(1'b1), .s(n761), .q(
        hcr_ic_ss_hcnt[4]) );
  drsp_1 r_ic_ss_hcnt_reg_7_ ( .ip(n1505), .ck(pclk), .rb(1'b1), .s(n4), .q(
        hcr_ic_ss_hcnt[7]) );
  drsp_1 r_ic_fs_hcnt_reg_4_ ( .ip(n1476), .ck(pclk), .rb(1'b1), .s(n3), .q(
        ic_fs_hcnt[4]) );
  drsp_1 r_ic_fs_hcnt_reg_3_ ( .ip(n1477), .ck(pclk), .rb(1'b1), .s(n2), .q(
        ic_fs_hcnt[3]) );
  nand3_1 U3 ( .ip1(n7), .ip2(n6), .ip3(n5), .op(ic_hcnt[1]) );
  nor4_1 U4 ( .ip1(ipwdata[14]), .ip2(ipwdata[12]), .ip3(ipwdata[13]), .ip4(
        ipwdata[15]), .op(n328) );
  buf_1 U5 ( .ip(n647), .op(n648) );
  inv_1 U6 ( .ip(presetn), .op(n2) );
  inv_1 U7 ( .ip(presetn), .op(n3) );
  inv_1 U8 ( .ip(presetn), .op(n4) );
  inv_1 U60 ( .ip(ic_con_pre_1_), .op(n477) );
  nand2_1 U61 ( .ip1(n477), .ip2(ic_fs_hcnt[1]), .op(n7) );
  inv_1 U62 ( .ip(ic_con_pre_2_), .op(n552) );
  nor2_1 U63 ( .ip1(n477), .ip2(n552), .op(ic_hs) );
  nand2_1 U64 ( .ip1(hcr_ic_hs_hcnt[1]), .ip2(ic_hs), .op(n6) );
  nor2_1 U65 ( .ip1(ic_con_pre_2_), .ip2(n477), .op(ic_ss) );
  nand2_1 U66 ( .ip1(hcr_ic_ss_hcnt[1]), .ip2(ic_ss), .op(n5) );
  nor2_1 U67 ( .ip1(reg_addr[0]), .ip2(reg_addr[5]), .op(n20) );
  nand2_1 U68 ( .ip1(reg_addr[1]), .ip2(n20), .op(n269) );
  inv_1 U69 ( .ip(reg_addr[4]), .op(n21) );
  inv_1 U70 ( .ip(reg_addr[2]), .op(n233) );
  nand3_1 U71 ( .ip1(n21), .ip2(n233), .ip3(reg_addr[3]), .op(n19) );
  nor2_1 U72 ( .ip1(n269), .ip2(n19), .op(n522) );
  inv_1 U73 ( .ip(reg_addr[0]), .op(n14) );
  nor2_1 U74 ( .ip1(reg_addr[5]), .ip2(n14), .op(n15) );
  nand2_1 U75 ( .ip1(reg_addr[1]), .ip2(n15), .op(n273) );
  inv_1 U76 ( .ip(reg_addr[3]), .op(n251) );
  nand3_1 U77 ( .ip1(reg_addr[2]), .ip2(n251), .ip3(n21), .op(n236) );
  nor2_1 U78 ( .ip1(n273), .ip2(n236), .op(n523) );
  and2_1 U79 ( .ip1(n523), .ip2(ic_fs_hcnt[13]), .op(n13) );
  nor2_1 U80 ( .ip1(n269), .ip2(n236), .op(n532) );
  nand2_1 U81 ( .ip1(n532), .ip2(hcr_ic_ss_lcnt[13]), .op(n11) );
  nand3_1 U82 ( .ip1(reg_addr[3]), .ip2(reg_addr[4]), .ip3(reg_addr[2]), .op(
        n294) );
  nor2_1 U83 ( .ip1(n273), .ip2(n294), .op(n646) );
  nand2_1 U84 ( .ip1(n646), .ip2(ic_sda_hold[13]), .op(n10) );
  inv_1 U85 ( .ip(n20), .op(n84) );
  or2_1 U86 ( .ip1(n19), .ip2(reg_addr[1]), .op(n111) );
  nor2_1 U87 ( .ip1(n84), .ip2(n111), .op(n524) );
  nand2_1 U88 ( .ip1(n524), .ip2(ic_fs_lcnt[13]), .op(n9) );
  nand3_1 U89 ( .ip1(n251), .ip2(n21), .ip3(n233), .op(n112) );
  or2_1 U90 ( .ip1(n112), .ip2(reg_addr[1]), .op(n83) );
  nand2_1 U91 ( .ip1(reg_addr[5]), .ip2(n14), .op(n101) );
  nor2_1 U92 ( .ip1(n83), .ip2(n101), .op(n549) );
  nand2_1 U93 ( .ip1(n549), .ip2(ic_tx_abrt_source[13]), .op(n8) );
  nand4_1 U94 ( .ip1(n11), .ip2(n10), .ip3(n9), .ip4(n8), .op(n12) );
  not_ab_or_c_or_d U95 ( .ip1(hcr_ic_hs_lcnt[13]), .ip2(n522), .ip3(n13), 
        .ip4(n12), .op(n18) );
  nand3_1 U96 ( .ip1(reg_addr[1]), .ip2(reg_addr[5]), .ip3(n14), .op(n235) );
  nor2_1 U97 ( .ip1(n235), .ip2(n294), .op(iprdata[29]) );
  inv_1 U98 ( .ip(iprdata[29]), .op(n548) );
  inv_1 U99 ( .ip(reg_addr[1]), .op(n296) );
  nand2_1 U100 ( .ip1(n15), .ip2(n296), .op(n267) );
  nor2_1 U101 ( .ip1(n267), .ip2(n236), .op(n533) );
  nand2_1 U102 ( .ip1(n533), .ip2(hcr_ic_ss_hcnt[13]), .op(n17) );
  inv_1 U103 ( .ip(n15), .op(n26) );
  nor2_1 U104 ( .ip1(n26), .ip2(n111), .op(n525) );
  nand2_1 U105 ( .ip1(n525), .ip2(hcr_ic_hs_hcnt[13]), .op(n16) );
  nand4_1 U106 ( .ip1(n18), .ip2(n548), .ip3(n17), .ip4(n16), .op(iprdata[13])
         );
  nor2_1 U107 ( .ip1(n273), .ip2(n19), .op(n499) );
  nand2_1 U108 ( .ip1(n499), .ip2(ic_intr_stat[11]), .op(n25) );
  nand2_1 U109 ( .ip1(n20), .ip2(n296), .op(n278) );
  nand3_1 U110 ( .ip1(reg_addr[3]), .ip2(reg_addr[2]), .ip3(n21), .op(n105) );
  nor2_1 U111 ( .ip1(n278), .ip2(n105), .op(n644) );
  nand2_1 U112 ( .ip1(n644), .ip2(ic_intr_mask[11]), .op(n24) );
  nor2_1 U113 ( .ip1(n267), .ip2(n105), .op(n485) );
  nand2_1 U114 ( .ip1(n485), .ip2(ic_raw_intr_stat[11]), .op(n23) );
  nand2_1 U115 ( .ip1(n533), .ip2(hcr_ic_ss_hcnt[11]), .op(n22) );
  and4_1 U116 ( .ip1(n25), .ip2(n24), .ip3(n23), .ip4(n22), .op(n36) );
  nor2_1 U117 ( .ip1(n26), .ip2(n83), .op(n587) );
  and2_1 U118 ( .ip1(n524), .ip2(ic_fs_lcnt[11]), .op(n32) );
  nand2_1 U119 ( .ip1(n522), .ip2(hcr_ic_hs_lcnt[11]), .op(n30) );
  nand2_1 U120 ( .ip1(n532), .ip2(hcr_ic_ss_lcnt[11]), .op(n29) );
  nand2_1 U121 ( .ip1(n523), .ip2(ic_fs_hcnt[11]), .op(n28) );
  nand2_1 U122 ( .ip1(n646), .ip2(ic_sda_hold[11]), .op(n27) );
  nand4_1 U123 ( .ip1(n30), .ip2(n29), .ip3(n28), .ip4(n27), .op(n31) );
  not_ab_or_c_or_d U124 ( .ip1(ic_tar[11]), .ip2(n587), .ip3(n32), .ip4(n31), 
        .op(n35) );
  nand2_1 U125 ( .ip1(n525), .ip2(hcr_ic_hs_hcnt[11]), .op(n34) );
  nand2_1 U126 ( .ip1(n549), .ip2(ic_tx_abrt_source[11]), .op(n33) );
  nand4_1 U127 ( .ip1(n36), .ip2(n35), .ip3(n34), .ip4(n33), .op(iprdata[11])
         );
  and2_1 U128 ( .ip1(n523), .ip2(ic_fs_hcnt[12]), .op(n42) );
  nand2_1 U129 ( .ip1(n532), .ip2(hcr_ic_ss_lcnt[12]), .op(n40) );
  nand2_1 U130 ( .ip1(n646), .ip2(ic_sda_hold[12]), .op(n39) );
  nand2_1 U131 ( .ip1(n524), .ip2(ic_fs_lcnt[12]), .op(n38) );
  nand2_1 U132 ( .ip1(n549), .ip2(ic_tx_abrt_source[12]), .op(n37) );
  nand4_1 U133 ( .ip1(n40), .ip2(n39), .ip3(n38), .ip4(n37), .op(n41) );
  not_ab_or_c_or_d U134 ( .ip1(hcr_ic_hs_lcnt[12]), .ip2(n522), .ip3(n42), 
        .ip4(n41), .op(n45) );
  nand2_1 U135 ( .ip1(n533), .ip2(hcr_ic_ss_hcnt[12]), .op(n44) );
  nand2_1 U136 ( .ip1(n525), .ip2(hcr_ic_hs_hcnt[12]), .op(n43) );
  nand4_1 U137 ( .ip1(n45), .ip2(n548), .ip3(n44), .ip4(n43), .op(iprdata[12])
         );
  and2_1 U138 ( .ip1(n499), .ip2(ic_intr_stat[10]), .op(n46) );
  nand2_1 U139 ( .ip1(reg_addr[0]), .ip2(reg_addr[5]), .op(n295) );
  nor3_1 U140 ( .ip1(reg_addr[1]), .ip2(n295), .ip3(n294), .op(n498) );
  not_ab_or_c_or_d U141 ( .ip1(n549), .ip2(ic_tx_abrt_source[10]), .ip3(n46), 
        .ip4(n498), .op(n59) );
  nand2_1 U142 ( .ip1(n644), .ip2(ic_intr_mask[10]), .op(n50) );
  nand2_1 U143 ( .ip1(ic_raw_intr_stat[10]), .ip2(n485), .op(n49) );
  nand2_1 U144 ( .ip1(n533), .ip2(hcr_ic_ss_hcnt[10]), .op(n48) );
  nand2_1 U145 ( .ip1(n522), .ip2(hcr_ic_hs_lcnt[10]), .op(n47) );
  nand4_1 U146 ( .ip1(n50), .ip2(n49), .ip3(n48), .ip4(n47), .op(n55) );
  nand2_1 U147 ( .ip1(ic_fs_hcnt[10]), .ip2(n523), .op(n53) );
  nand2_1 U148 ( .ip1(n532), .ip2(hcr_ic_ss_lcnt[10]), .op(n52) );
  nand2_1 U149 ( .ip1(n646), .ip2(ic_sda_hold[10]), .op(n51) );
  nand3_1 U150 ( .ip1(n53), .ip2(n52), .ip3(n51), .op(n54) );
  not_ab_or_c_or_d U151 ( .ip1(n587), .ip2(ic_tar[10]), .ip3(n55), .ip4(n54), 
        .op(n58) );
  nand2_1 U152 ( .ip1(n524), .ip2(ic_fs_lcnt[10]), .op(n57) );
  nand2_1 U153 ( .ip1(n525), .ip2(hcr_ic_hs_hcnt[10]), .op(n56) );
  nand4_1 U154 ( .ip1(n59), .ip2(n58), .ip3(n57), .ip4(n56), .op(iprdata[10])
         );
  nor2_1 U155 ( .ip1(n269), .ip2(n112), .op(n586) );
  not_ab_or_c_or_d U156 ( .ip1(n586), .ip2(ic_sar[9]), .ip3(iprdata[29]), 
        .ip4(n498), .op(n74) );
  nand2_1 U157 ( .ip1(n524), .ip2(ic_fs_lcnt[9]), .op(n62) );
  nand2_1 U158 ( .ip1(n532), .ip2(hcr_ic_ss_lcnt[9]), .op(n61) );
  nand2_1 U159 ( .ip1(n646), .ip2(ic_sda_hold[9]), .op(n60) );
  nand3_1 U160 ( .ip1(n62), .ip2(n61), .ip3(n60), .op(n70) );
  and2_1 U161 ( .ip1(n533), .ip2(hcr_ic_ss_hcnt[9]), .op(n64) );
  and2_1 U162 ( .ip1(n523), .ip2(ic_fs_hcnt[9]), .op(n63) );
  not_ab_or_c_or_d U163 ( .ip1(n522), .ip2(hcr_ic_hs_lcnt[9]), .ip3(n64), 
        .ip4(n63), .op(n68) );
  nand2_1 U164 ( .ip1(n525), .ip2(hcr_ic_hs_hcnt[9]), .op(n67) );
  nand2_1 U165 ( .ip1(n549), .ip2(ic_tx_abrt_source[9]), .op(n66) );
  nand2_1 U166 ( .ip1(ic_raw_intr_stat[9]), .ip2(n485), .op(n65) );
  nand4_1 U167 ( .ip1(n68), .ip2(n67), .ip3(n66), .ip4(n65), .op(n69) );
  not_ab_or_c_or_d U168 ( .ip1(n587), .ip2(ic_tar[9]), .ip3(n70), .ip4(n69), 
        .op(n73) );
  nand2_1 U169 ( .ip1(n499), .ip2(ic_intr_stat[9]), .op(n72) );
  nand2_1 U170 ( .ip1(n644), .ip2(ic_intr_mask[9]), .op(n71) );
  nand4_1 U171 ( .ip1(n74), .ip2(n73), .ip3(n72), .ip4(n71), .op(iprdata[9])
         );
  nand2_1 U172 ( .ip1(n644), .ip2(ic_intr_mask[8]), .op(n78) );
  nand2_1 U173 ( .ip1(n586), .ip2(ic_sar[8]), .op(n77) );
  nand2_1 U174 ( .ip1(n485), .ip2(ic_raw_intr_stat[8]), .op(n76) );
  nand2_1 U175 ( .ip1(n522), .ip2(hcr_ic_hs_lcnt[8]), .op(n75) );
  nand4_1 U176 ( .ip1(n78), .ip2(n77), .ip3(n76), .ip4(n75), .op(n91) );
  nand2_1 U177 ( .ip1(n533), .ip2(hcr_ic_ss_hcnt[8]), .op(n82) );
  nand2_1 U178 ( .ip1(n523), .ip2(ic_fs_hcnt[8]), .op(n81) );
  nand2_1 U179 ( .ip1(n532), .ip2(hcr_ic_ss_lcnt[8]), .op(n80) );
  nand2_1 U180 ( .ip1(n646), .ip2(ic_sda_hold[8]), .op(n79) );
  nand4_1 U181 ( .ip1(n82), .ip2(n81), .ip3(n80), .ip4(n79), .op(n90) );
  nor2_1 U182 ( .ip1(n84), .ip2(n83), .op(n582) );
  nand2_1 U183 ( .ip1(n582), .ip2(tx_empty_ctrl), .op(n88) );
  nand2_1 U184 ( .ip1(n587), .ip2(ic_tar[8]), .op(n87) );
  nand2_1 U185 ( .ip1(n524), .ip2(ic_fs_lcnt[8]), .op(n86) );
  nand2_1 U186 ( .ip1(n525), .ip2(hcr_ic_hs_hcnt[8]), .op(n85) );
  nand4_1 U187 ( .ip1(n88), .ip2(n87), .ip3(n86), .ip4(n85), .op(n89) );
  nor3_1 U188 ( .ip1(n91), .ip2(n90), .ip3(n89), .op(n94) );
  or2_1 U189 ( .ip1(n295), .ip2(n294), .op(n541) );
  nand2_1 U190 ( .ip1(n499), .ip2(ic_intr_stat[8]), .op(n93) );
  nand2_1 U191 ( .ip1(n549), .ip2(ic_tx_abrt_source[8]), .op(n92) );
  nand4_1 U192 ( .ip1(n94), .ip2(n541), .ip3(n93), .ip4(n92), .op(iprdata[8])
         );
  and2_1 U193 ( .ip1(n644), .ip2(ic_intr_mask[2]), .op(n100) );
  nor2_1 U194 ( .ip1(n278), .ip2(n236), .op(n506) );
  nand2_1 U195 ( .ip1(n506), .ip2(rx_pop_data[2]), .op(n98) );
  nand2_1 U196 ( .ip1(n485), .ip2(ic_raw_intr_stat[2]), .op(n97) );
  nor2_1 U197 ( .ip1(n269), .ip2(n294), .op(n486) );
  nand2_1 U198 ( .ip1(n486), .ip2(ic_rxflr[2]), .op(n96) );
  nor2_1 U199 ( .ip1(n278), .ip2(n294), .op(n302) );
  nand2_1 U200 ( .ip1(n302), .ip2(tx_empty), .op(n95) );
  nand4_1 U201 ( .ip1(n98), .ip2(n97), .ip3(n96), .ip4(n95), .op(n99) );
  not_ab_or_c_or_d U202 ( .ip1(n586), .ip2(ic_sar[2]), .ip3(n100), .ip4(n99), 
        .op(n128) );
  nor2_1 U203 ( .ip1(n111), .ip2(n101), .op(n638) );
  nand2_1 U204 ( .ip1(n638), .ip2(ic_fs_spklen[2]), .op(n104) );
  nand2_1 U205 ( .ip1(n582), .ip2(ic_con_pre_2_), .op(n103) );
  nand2_1 U206 ( .ip1(n524), .ip2(ic_fs_lcnt[2]), .op(n102) );
  nand3_1 U207 ( .ip1(n104), .ip2(n103), .ip3(n102), .op(n124) );
  nor2_1 U208 ( .ip1(n269), .ip2(n105), .op(n679) );
  nand2_1 U209 ( .ip1(n549), .ip2(ic_tx_abrt_source[2]), .op(n109) );
  nand2_1 U210 ( .ip1(n525), .ip2(hcr_ic_hs_hcnt[2]), .op(n108) );
  nor3_1 U211 ( .ip1(n296), .ip2(n295), .ip3(n236), .op(n276) );
  nand2_1 U212 ( .ip1(n276), .ip2(slv_fifo_filled_and_flushed_sync), .op(n107)
         );
  nor2_1 U213 ( .ip1(n273), .ip2(n105), .op(n684) );
  nand2_1 U214 ( .ip1(n684), .ip2(ic_tx_tl_2_), .op(n106) );
  nand4_1 U215 ( .ip1(n109), .ip2(n108), .ip3(n107), .ip4(n106), .op(n110) );
  not_ab_or_c_or_d U216 ( .ip1(n679), .ip2(ic_rx_tl_int[2]), .ip3(n498), .ip4(
        n110), .op(n122) );
  and2_1 U217 ( .ip1(n523), .ip2(ic_fs_hcnt[2]), .op(n118) );
  nand2_1 U218 ( .ip1(n532), .ip2(hcr_ic_ss_lcnt[2]), .op(n116) );
  nand2_1 U219 ( .ip1(n646), .ip2(ic_sda_hold[2]), .op(n115) );
  nor2_1 U220 ( .ip1(n295), .ip2(n111), .op(n641) );
  nand2_1 U221 ( .ip1(n641), .ip2(ic_hs_spklen[2]), .op(n114) );
  nor2_1 U222 ( .ip1(n273), .ip2(n112), .op(n677) );
  nand2_1 U223 ( .ip1(n677), .ip2(ic_hs_maddr[2]), .op(n113) );
  nand4_1 U224 ( .ip1(n116), .ip2(n115), .ip3(n114), .ip4(n113), .op(n117) );
  not_ab_or_c_or_d U225 ( .ip1(hcr_ic_ss_hcnt[2]), .ip2(n533), .ip3(n118), 
        .ip4(n117), .op(n121) );
  nand2_1 U226 ( .ip1(n522), .ip2(hcr_ic_hs_lcnt[2]), .op(n120) );
  nor2_1 U227 ( .ip1(n267), .ip2(n294), .op(n487) );
  nand2_1 U228 ( .ip1(n487), .ip2(ic_txflr[2]), .op(n119) );
  nand4_1 U229 ( .ip1(n122), .ip2(n121), .ip3(n120), .ip4(n119), .op(n123) );
  not_ab_or_c_or_d U230 ( .ip1(n587), .ip2(ic_tar[2]), .ip3(n124), .ip4(n123), 
        .op(n127) );
  nor3_1 U231 ( .ip1(reg_addr[1]), .ip2(n295), .ip3(n236), .op(n690) );
  nand2_1 U232 ( .ip1(n690), .ip2(ic_sda_setup[2]), .op(n126) );
  nand2_1 U233 ( .ip1(n499), .ip2(ic_intr_stat[2]), .op(n125) );
  nand4_1 U234 ( .ip1(n128), .ip2(n127), .ip3(n126), .ip4(n125), .op(
        iprdata[2]) );
  nand2_1 U235 ( .ip1(n533), .ip2(hcr_ic_ss_hcnt[4]), .op(n132) );
  nand2_1 U236 ( .ip1(n302), .ip2(rx_full), .op(n131) );
  nand2_1 U237 ( .ip1(n522), .ip2(hcr_ic_hs_lcnt[4]), .op(n130) );
  nand2_1 U238 ( .ip1(n523), .ip2(ic_fs_hcnt[4]), .op(n129) );
  and4_1 U239 ( .ip1(n132), .ip2(n131), .ip3(n130), .ip4(n129), .op(n151) );
  and2_1 U240 ( .ip1(n644), .ip2(ic_intr_mask[4]), .op(n138) );
  nand2_1 U241 ( .ip1(n499), .ip2(ic_intr_stat[4]), .op(n136) );
  nand2_1 U242 ( .ip1(n690), .ip2(ic_sda_setup[4]), .op(n135) );
  nand2_1 U243 ( .ip1(n506), .ip2(rx_pop_data[4]), .op(n134) );
  nand2_1 U244 ( .ip1(n485), .ip2(ic_raw_intr_stat[4]), .op(n133) );
  nand4_1 U245 ( .ip1(n136), .ip2(n135), .ip3(n134), .ip4(n133), .op(n137) );
  not_ab_or_c_or_d U246 ( .ip1(n586), .ip2(ic_sar[4]), .ip3(n138), .ip4(n137), 
        .op(n150) );
  nand2_1 U247 ( .ip1(n638), .ip2(ic_fs_spklen[4]), .op(n141) );
  nand2_1 U248 ( .ip1(n532), .ip2(hcr_ic_ss_lcnt[4]), .op(n140) );
  nand2_1 U249 ( .ip1(n646), .ip2(ic_sda_hold[4]), .op(n139) );
  nand3_1 U250 ( .ip1(n141), .ip2(n140), .ip3(n139), .op(n147) );
  nand2_1 U251 ( .ip1(n582), .ip2(ic_10bit_mst), .op(n145) );
  nand2_1 U252 ( .ip1(n587), .ip2(ic_tar[4]), .op(n144) );
  nand2_1 U253 ( .ip1(n524), .ip2(ic_fs_lcnt[4]), .op(n143) );
  nand2_1 U254 ( .ip1(n549), .ip2(ic_tx_abrt_source[4]), .op(n142) );
  nand4_1 U255 ( .ip1(n145), .ip2(n144), .ip3(n143), .ip4(n142), .op(n146) );
  not_ab_or_c_or_d U256 ( .ip1(n641), .ip2(ic_hs_spklen[4]), .ip3(n147), .ip4(
        n146), .op(n149) );
  nand2_1 U257 ( .ip1(n525), .ip2(hcr_ic_hs_hcnt[4]), .op(n148) );
  nand4_1 U258 ( .ip1(n151), .ip2(n150), .ip3(n149), .ip4(n148), .op(
        iprdata[4]) );
  nand2_1 U259 ( .ip1(ic_raw_intr_stat[7]), .ip2(n485), .op(n155) );
  nand2_1 U260 ( .ip1(n533), .ip2(hcr_ic_ss_hcnt[7]), .op(n154) );
  nand2_1 U261 ( .ip1(n522), .ip2(hcr_ic_hs_lcnt[7]), .op(n153) );
  nand2_1 U262 ( .ip1(n523), .ip2(ic_fs_hcnt[7]), .op(n152) );
  and4_1 U263 ( .ip1(n155), .ip2(n154), .ip3(n153), .ip4(n152), .op(n173) );
  nand2_1 U264 ( .ip1(n690), .ip2(ic_sda_setup[7]), .op(n159) );
  nand2_1 U265 ( .ip1(n644), .ip2(ic_intr_mask[7]), .op(n158) );
  nand2_1 U266 ( .ip1(n586), .ip2(ic_sar[7]), .op(n157) );
  nand2_1 U267 ( .ip1(n506), .ip2(rx_pop_data[7]), .op(n156) );
  nand4_1 U268 ( .ip1(n159), .ip2(n158), .ip3(n157), .ip4(n156), .op(n160) );
  not_ab_or_c_or_d U269 ( .ip1(n499), .ip2(ic_intr_stat[7]), .ip3(n498), .ip4(
        n160), .op(n172) );
  nand2_1 U270 ( .ip1(n638), .ip2(ic_fs_spklen[7]), .op(n163) );
  nand2_1 U271 ( .ip1(n532), .ip2(hcr_ic_ss_lcnt[7]), .op(n162) );
  nand2_1 U272 ( .ip1(n646), .ip2(ic_sda_hold[7]), .op(n161) );
  nand3_1 U273 ( .ip1(n163), .ip2(n162), .ip3(n161), .op(n169) );
  nand2_1 U274 ( .ip1(n582), .ip2(p_det_ifaddr), .op(n167) );
  nand2_1 U275 ( .ip1(n587), .ip2(ic_tar[7]), .op(n166) );
  nand2_1 U276 ( .ip1(n524), .ip2(ic_fs_lcnt[7]), .op(n165) );
  nand2_1 U277 ( .ip1(n549), .ip2(ic_tx_abrt_source[7]), .op(n164) );
  nand4_1 U278 ( .ip1(n167), .ip2(n166), .ip3(n165), .ip4(n164), .op(n168) );
  not_ab_or_c_or_d U279 ( .ip1(n641), .ip2(ic_hs_spklen[7]), .ip3(n169), .ip4(
        n168), .op(n171) );
  nand2_1 U280 ( .ip1(n525), .ip2(hcr_ic_hs_hcnt[7]), .op(n170) );
  nand4_1 U281 ( .ip1(n173), .ip2(n172), .ip3(n171), .ip4(n170), .op(
        iprdata[7]) );
  inv_1 U282 ( .ip(n302), .op(n484) );
  nor2_1 U283 ( .ip1(tx_full), .ip2(n484), .op(n179) );
  nand2_1 U284 ( .ip1(n506), .ip2(rx_pop_data[1]), .op(n177) );
  nand2_1 U285 ( .ip1(ic_raw_intr_stat[1]), .ip2(n485), .op(n176) );
  nand2_1 U286 ( .ip1(n487), .ip2(ic_txflr[1]), .op(n175) );
  nand2_1 U287 ( .ip1(n522), .ip2(hcr_ic_hs_lcnt[1]), .op(n174) );
  nand4_1 U288 ( .ip1(n177), .ip2(n176), .ip3(n175), .ip4(n174), .op(n178) );
  not_ab_or_c_or_d U289 ( .ip1(ic_rxflr[1]), .ip2(n486), .ip3(n179), .ip4(n178), .op(n204) );
  nand2_1 U290 ( .ip1(n582), .ip2(ic_con_pre_1_), .op(n182) );
  nand2_1 U291 ( .ip1(n524), .ip2(ic_fs_lcnt[1]), .op(n181) );
  nand2_1 U292 ( .ip1(n549), .ip2(ic_tx_abrt_source[1]), .op(n180) );
  nand3_1 U293 ( .ip1(n182), .ip2(n181), .ip3(n180), .op(n200) );
  and2_1 U294 ( .ip1(n684), .ip2(ic_tx_tl_1_), .op(n188) );
  nand2_1 U295 ( .ip1(n679), .ip2(ic_rx_tl_int[1]), .op(n186) );
  nand3_1 U296 ( .ip1(reg_addr[4]), .ip2(reg_addr[3]), .ip3(n233), .op(n272)
         );
  nor2_1 U297 ( .ip1(n273), .ip2(n272), .op(n322) );
  nand2_1 U298 ( .ip1(n322), .ip2(ic_enable[1]), .op(n185) );
  nand2_1 U299 ( .ip1(n499), .ip2(ic_intr_stat[1]), .op(n184) );
  nand2_1 U300 ( .ip1(n690), .ip2(ic_sda_setup[1]), .op(n183) );
  nand4_1 U301 ( .ip1(n186), .ip2(n185), .ip3(n184), .ip4(n183), .op(n187) );
  not_ab_or_c_or_d U302 ( .ip1(slv_rx_aborted_sync), .ip2(n276), .ip3(n188), 
        .ip4(n187), .op(n198) );
  not_ab_or_c_or_d U303 ( .ip1(n677), .ip2(ic_hs_maddr[1]), .ip3(iprdata[29]), 
        .ip4(n498), .op(n197) );
  and2_1 U304 ( .ip1(n523), .ip2(ic_fs_hcnt[1]), .op(n194) );
  nand2_1 U305 ( .ip1(n532), .ip2(hcr_ic_ss_lcnt[1]), .op(n192) );
  nand2_1 U306 ( .ip1(n646), .ip2(ic_sda_hold[1]), .op(n191) );
  nand2_1 U307 ( .ip1(n641), .ip2(ic_hs_spklen[1]), .op(n190) );
  nand2_1 U308 ( .ip1(n638), .ip2(ic_fs_spklen[1]), .op(n189) );
  nand4_1 U309 ( .ip1(n192), .ip2(n191), .ip3(n190), .ip4(n189), .op(n193) );
  not_ab_or_c_or_d U310 ( .ip1(hcr_ic_ss_hcnt[1]), .ip2(n533), .ip3(n194), 
        .ip4(n193), .op(n196) );
  nand2_1 U311 ( .ip1(n525), .ip2(hcr_ic_hs_hcnt[1]), .op(n195) );
  nand4_1 U312 ( .ip1(n198), .ip2(n197), .ip3(n196), .ip4(n195), .op(n199) );
  not_ab_or_c_or_d U313 ( .ip1(n587), .ip2(ic_tar[1]), .ip3(n200), .ip4(n199), 
        .op(n203) );
  nand2_1 U314 ( .ip1(n644), .ip2(ic_intr_mask[1]), .op(n202) );
  nand2_1 U315 ( .ip1(n586), .ip2(ic_sar[1]), .op(n201) );
  nand4_1 U316 ( .ip1(n204), .ip2(n203), .ip3(n202), .ip4(n201), .op(
        iprdata[1]) );
  nand2_1 U317 ( .ip1(n586), .ip2(ic_sar[5]), .op(n208) );
  nand2_1 U318 ( .ip1(n506), .ip2(rx_pop_data[5]), .op(n207) );
  nand2_1 U319 ( .ip1(ic_raw_intr_stat[5]), .ip2(n485), .op(n206) );
  nand2_1 U320 ( .ip1(n522), .ip2(hcr_ic_hs_lcnt[5]), .op(n205) );
  nand4_1 U321 ( .ip1(n208), .ip2(n207), .ip3(n206), .ip4(n205), .op(n209) );
  not_ab_or_c_or_d U322 ( .ip1(n499), .ip2(ic_intr_stat[5]), .ip3(iprdata[29]), 
        .ip4(n209), .op(n228) );
  nand2_1 U323 ( .ip1(n302), .ip2(mst_activity_r), .op(n213) );
  nand2_1 U324 ( .ip1(n533), .ip2(hcr_ic_ss_hcnt[5]), .op(n212) );
  nand2_1 U325 ( .ip1(n646), .ip2(ic_sda_hold[5]), .op(n211) );
  nand2_1 U326 ( .ip1(n523), .ip2(ic_fs_hcnt[5]), .op(n210) );
  nand4_1 U327 ( .ip1(n213), .ip2(n212), .ip3(n211), .ip4(n210), .op(n224) );
  nand2_1 U328 ( .ip1(n641), .ip2(ic_hs_spklen[5]), .op(n217) );
  nand2_1 U329 ( .ip1(n638), .ip2(ic_fs_spklen[5]), .op(n216) );
  nand2_1 U330 ( .ip1(n582), .ip2(ic_rstrt_en), .op(n215) );
  nand2_1 U331 ( .ip1(n532), .ip2(hcr_ic_ss_lcnt[5]), .op(n214) );
  nand4_1 U332 ( .ip1(n217), .ip2(n216), .ip3(n215), .ip4(n214), .op(n223) );
  nand2_1 U333 ( .ip1(n587), .ip2(ic_tar[5]), .op(n221) );
  nand2_1 U334 ( .ip1(n524), .ip2(ic_fs_lcnt[5]), .op(n220) );
  nand2_1 U335 ( .ip1(n549), .ip2(ic_tx_abrt_source[5]), .op(n219) );
  nand2_1 U336 ( .ip1(n525), .ip2(hcr_ic_hs_hcnt[5]), .op(n218) );
  nand4_1 U337 ( .ip1(n221), .ip2(n220), .ip3(n219), .ip4(n218), .op(n222) );
  nor3_1 U338 ( .ip1(n224), .ip2(n223), .ip3(n222), .op(n227) );
  nand2_1 U339 ( .ip1(n690), .ip2(ic_sda_setup[5]), .op(n226) );
  nand2_1 U340 ( .ip1(n644), .ip2(ic_intr_mask[5]), .op(n225) );
  nand4_1 U341 ( .ip1(n228), .ip2(n227), .ip3(n226), .ip4(n225), .op(
        iprdata[5]) );
  nor2_1 U342 ( .ip1(n278), .ip2(n272), .op(ic_clr_stop_det_en) );
  nand2_1 U343 ( .ip1(ic_clr_stop_det_en), .ip2(ic_raw_intr_stat[9]), .op(n232) );
  nor2_1 U344 ( .ip1(n267), .ip2(n272), .op(ic_clr_start_det_en) );
  inv_1 U345 ( .ip(ic_clr_start_det_en), .op(n230) );
  nor2_1 U346 ( .ip1(ic_raw_intr_stat[10]), .ip2(n230), .op(n229) );
  or2_1 U347 ( .ip1(n230), .ip2(n229), .op(n231) );
  nand2_1 U348 ( .ip1(n232), .ip2(n231), .op(n241) );
  nand2_1 U349 ( .ip1(n587), .ip2(ic_tar[0]), .op(n239) );
  nand3_1 U350 ( .ip1(reg_addr[4]), .ip2(n251), .ip3(n233), .op(n277) );
  nor2_1 U351 ( .ip1(n267), .ip2(n277), .op(ic_clr_rx_under_en) );
  or2_1 U352 ( .ip1(n485), .ip2(ic_clr_rx_under_en), .op(n234) );
  nand2_1 U353 ( .ip1(ic_raw_intr_stat[0]), .ip2(n234), .op(n238) );
  nor2_1 U354 ( .ip1(n236), .ip2(n235), .op(n708) );
  nand2_1 U355 ( .ip1(ic_ack_general_call), .ip2(n708), .op(n237) );
  nand3_1 U356 ( .ip1(n239), .ip2(n238), .ip3(n237), .op(n240) );
  not_ab_or_c_or_d U357 ( .ip1(n641), .ip2(ic_hs_spklen[0]), .ip3(n241), .ip4(
        n240), .op(n293) );
  nor2_1 U358 ( .ip1(n269), .ip2(n272), .op(ic_clr_gen_call_en) );
  nand2_1 U359 ( .ip1(ic_txflr[0]), .ip2(n487), .op(n245) );
  nand2_1 U360 ( .ip1(n522), .ip2(hcr_ic_hs_lcnt[0]), .op(n244) );
  nand2_1 U361 ( .ip1(n533), .ip2(hcr_ic_ss_hcnt[0]), .op(n243) );
  nand2_1 U362 ( .ip1(n523), .ip2(ic_fs_hcnt[0]), .op(n242) );
  nand4_1 U363 ( .ip1(n245), .ip2(n244), .ip3(n243), .ip4(n242), .op(n250) );
  nand2_1 U364 ( .ip1(n532), .ip2(hcr_ic_ss_lcnt[0]), .op(n248) );
  nand2_1 U365 ( .ip1(ic_sda_hold[0]), .ip2(n646), .op(n247) );
  nand2_1 U366 ( .ip1(ic_hs_maddr[0]), .ip2(n677), .op(n246) );
  nand3_1 U367 ( .ip1(n248), .ip2(n247), .ip3(n246), .op(n249) );
  not_ab_or_c_or_d U368 ( .ip1(ic_clr_gen_call_en), .ip2(ic_raw_intr_stat[11]), 
        .ip3(n250), .ip4(n249), .op(n292) );
  nand3_1 U369 ( .ip1(reg_addr[4]), .ip2(reg_addr[2]), .ip3(n251), .op(n270)
         );
  nor2_1 U370 ( .ip1(n273), .ip2(n270), .op(ic_clr_activity_en) );
  nand2_1 U371 ( .ip1(n690), .ip2(ic_sda_setup[0]), .op(n255) );
  nand2_1 U372 ( .ip1(n499), .ip2(ic_intr_stat[0]), .op(n254) );
  nand2_1 U373 ( .ip1(n644), .ip2(ic_intr_mask[0]), .op(n253) );
  nand2_1 U374 ( .ip1(n586), .ip2(ic_sar[0]), .op(n252) );
  nand4_1 U375 ( .ip1(n255), .ip2(n254), .ip3(n253), .ip4(n252), .op(n260) );
  nand2_1 U376 ( .ip1(n506), .ip2(rx_pop_data[0]), .op(n258) );
  nand2_1 U377 ( .ip1(ic_rxflr[0]), .ip2(n486), .op(n257) );
  nand2_1 U378 ( .ip1(n302), .ip2(activity_r), .op(n256) );
  nand3_1 U379 ( .ip1(n258), .ip2(n257), .ip3(n256), .op(n259) );
  not_ab_or_c_or_d U380 ( .ip1(ic_clr_activity_en), .ip2(ic_raw_intr_stat[8]), 
        .ip3(n260), .ip4(n259), .op(n291) );
  nand2_1 U381 ( .ip1(ic_fs_spklen[0]), .ip2(n638), .op(n264) );
  nand2_1 U382 ( .ip1(ic_master), .ip2(n582), .op(n263) );
  nand2_1 U383 ( .ip1(n524), .ip2(ic_fs_lcnt[0]), .op(n262) );
  nand2_1 U384 ( .ip1(n549), .ip2(ic_tx_abrt_source[0]), .op(n261) );
  nand4_1 U385 ( .ip1(n264), .ip2(n263), .ip3(n262), .ip4(n261), .op(n289) );
  nor2_1 U386 ( .ip1(n269), .ip2(n277), .op(ic_clr_rx_over_en) );
  and2_1 U387 ( .ip1(ic_clr_rx_over_en), .ip2(ic_raw_intr_stat[1]), .op(n265)
         );
  nor2_1 U388 ( .ip1(n273), .ip2(n277), .op(ic_clr_tx_over_en) );
  mux2_1 U389 ( .ip1(n265), .ip2(ic_raw_intr_stat[3]), .s(ic_clr_tx_over_en), 
        .op(n266) );
  nor2_1 U390 ( .ip1(n270), .ip2(n278), .op(ic_clr_rd_req_en) );
  mux2_1 U391 ( .ip1(n266), .ip2(ic_raw_intr_stat[5]), .s(ic_clr_rd_req_en), 
        .op(n268) );
  nor2_1 U392 ( .ip1(n270), .ip2(n267), .op(ic_clr_tx_abrt_en) );
  inv_1 U393 ( .ip(ic_clr_tx_abrt_en), .op(n383) );
  mux2_1 U394 ( .ip1(ic_raw_intr_stat[6]), .ip2(n268), .s(n383), .op(n271) );
  nor2_1 U395 ( .ip1(n270), .ip2(n269), .op(ic_clr_rx_done_en) );
  mux2_1 U396 ( .ip1(n271), .ip2(ic_raw_intr_stat[7]), .s(ic_clr_rx_done_en), 
        .op(n288) );
  inv_1 U397 ( .ip(ic_enable[0]), .op(n703) );
  nor3_1 U398 ( .ip1(n273), .ip2(n272), .ip3(n703), .op(n275) );
  and2_1 U399 ( .ip1(ic_tx_tl_0_), .ip2(n684), .op(n274) );
  not_ab_or_c_or_d U400 ( .ip1(n276), .ip2(ic_en), .ip3(n275), .ip4(n274), 
        .op(n286) );
  nand2_1 U401 ( .ip1(n525), .ip2(hcr_ic_hs_hcnt[0]), .op(n285) );
  nor2_1 U402 ( .ip1(n278), .ip2(n277), .op(ic_clr_intr_en) );
  nor4_1 U403 ( .ip1(ic_raw_intr_stat[1]), .ip2(ic_raw_intr_stat[3]), .ip3(
        ic_raw_intr_stat[0]), .ip4(ic_raw_intr_stat[2]), .op(n281) );
  nor4_1 U404 ( .ip1(ic_raw_intr_stat[9]), .ip2(ic_raw_intr_stat[10]), .ip3(
        ic_raw_intr_stat[11]), .ip4(ic_raw_intr_stat[4]), .op(n280) );
  nor4_1 U405 ( .ip1(ic_raw_intr_stat[5]), .ip2(ic_raw_intr_stat[6]), .ip3(
        ic_raw_intr_stat[7]), .ip4(ic_raw_intr_stat[8]), .op(n279) );
  nand3_1 U406 ( .ip1(n281), .ip2(n280), .ip3(n279), .op(n282) );
  nand2_1 U407 ( .ip1(ic_clr_intr_en), .ip2(n282), .op(n284) );
  nand2_1 U408 ( .ip1(ic_rx_tl_int[0]), .ip2(n679), .op(n283) );
  nand4_1 U409 ( .ip1(n286), .ip2(n285), .ip3(n284), .ip4(n283), .op(n287) );
  nor3_1 U410 ( .ip1(n289), .ip2(n288), .ip3(n287), .op(n290) );
  nand4_1 U411 ( .ip1(n293), .ip2(n292), .ip3(n291), .ip4(n290), .op(
        iprdata[0]) );
  nor3_1 U412 ( .ip1(n296), .ip2(n295), .ip3(n294), .op(iprdata[30]) );
  nand2_1 U413 ( .ip1(n586), .ip2(ic_sar[6]), .op(n300) );
  nand2_1 U414 ( .ip1(n506), .ip2(rx_pop_data[6]), .op(n299) );
  nand2_1 U415 ( .ip1(ic_raw_intr_stat[6]), .ip2(n485), .op(n298) );
  nand2_1 U416 ( .ip1(n522), .ip2(hcr_ic_hs_lcnt[6]), .op(n297) );
  nand4_1 U417 ( .ip1(n300), .ip2(n299), .ip3(n298), .ip4(n297), .op(n301) );
  not_ab_or_c_or_d U418 ( .ip1(n499), .ip2(ic_intr_stat[6]), .ip3(iprdata[30]), 
        .ip4(n301), .op(n321) );
  nand2_1 U419 ( .ip1(n302), .ip2(slv_activity_r), .op(n306) );
  nand2_1 U420 ( .ip1(n533), .ip2(hcr_ic_ss_hcnt[6]), .op(n305) );
  nand2_1 U421 ( .ip1(n646), .ip2(ic_sda_hold[6]), .op(n304) );
  nand2_1 U422 ( .ip1(n523), .ip2(ic_fs_hcnt[6]), .op(n303) );
  nand4_1 U423 ( .ip1(n306), .ip2(n305), .ip3(n304), .ip4(n303), .op(n317) );
  nand2_1 U424 ( .ip1(n641), .ip2(ic_hs_spklen[6]), .op(n310) );
  nand2_1 U425 ( .ip1(n638), .ip2(ic_fs_spklen[6]), .op(n309) );
  nand2_1 U426 ( .ip1(n582), .ip2(ic_con_pre_6_), .op(n308) );
  nand2_1 U427 ( .ip1(n532), .ip2(hcr_ic_ss_lcnt[6]), .op(n307) );
  nand4_1 U428 ( .ip1(n310), .ip2(n309), .ip3(n308), .ip4(n307), .op(n316) );
  nand2_1 U429 ( .ip1(n587), .ip2(ic_tar[6]), .op(n314) );
  nand2_1 U430 ( .ip1(n524), .ip2(ic_fs_lcnt[6]), .op(n313) );
  nand2_1 U431 ( .ip1(n549), .ip2(ic_tx_abrt_source[6]), .op(n312) );
  nand2_1 U432 ( .ip1(n525), .ip2(hcr_ic_hs_hcnt[6]), .op(n311) );
  nand4_1 U433 ( .ip1(n314), .ip2(n313), .ip3(n312), .ip4(n311), .op(n315) );
  nor3_1 U434 ( .ip1(n317), .ip2(n316), .ip3(n315), .op(n320) );
  nand2_1 U435 ( .ip1(n690), .ip2(ic_sda_setup[6]), .op(n319) );
  nand2_1 U436 ( .ip1(n644), .ip2(ic_intr_mask[6]), .op(n318) );
  nand4_1 U437 ( .ip1(n321), .ip2(n320), .ip3(n319), .ip4(n318), .op(
        iprdata[6]) );
  nand2_1 U438 ( .ip1(n506), .ip2(rd_en), .op(n558) );
  inv_1 U439 ( .ip(n558), .op(rx_pop) );
  nand2_1 U440 ( .ip1(n322), .ip2(wr_en), .op(n553) );
  nor2_1 U441 ( .ip1(ipwdata[0]), .ip2(n553), .op(n382) );
  or2_1 U442 ( .ip1(n703), .ip2(n382), .op(n324) );
  or2_1 U443 ( .ip1(n553), .ip2(n382), .op(n323) );
  nand2_1 U444 ( .ip1(n324), .ip2(n323), .op(n1549) );
  inv_1 U445 ( .ip(presetn), .op(n761) );
  and2_1 U446 ( .ip1(n703), .ip2(wr_en), .op(n689) );
  nand2_1 U447 ( .ip1(n524), .ip2(n689), .op(n620) );
  mux2_1 U448 ( .ip1(ipwdata[14]), .ip2(ic_fs_lcnt[14]), .s(n620), .op(n1449)
         );
  mux2_1 U449 ( .ip1(ipwdata[13]), .ip2(ic_fs_lcnt[13]), .s(n620), .op(n1450)
         );
  mux2_1 U450 ( .ip1(ipwdata[12]), .ip2(ic_fs_lcnt[12]), .s(n620), .op(n1451)
         );
  mux2_1 U451 ( .ip1(ipwdata[11]), .ip2(ic_fs_lcnt[11]), .s(n620), .op(n1452)
         );
  mux2_1 U452 ( .ip1(ipwdata[10]), .ip2(ic_fs_lcnt[10]), .s(n620), .op(n1453)
         );
  mux2_1 U453 ( .ip1(ipwdata[9]), .ip2(ic_fs_lcnt[9]), .s(n620), .op(n1454) );
  mux2_1 U454 ( .ip1(ipwdata[8]), .ip2(ic_fs_lcnt[8]), .s(n620), .op(n1455) );
  mux2_1 U455 ( .ip1(ipwdata[15]), .ip2(ic_fs_lcnt[15]), .s(n620), .op(n1456)
         );
  inv_1 U456 ( .ip(ipwdata[5]), .op(n326) );
  inv_1 U457 ( .ip(ipwdata[6]), .op(n325) );
  nand2_1 U458 ( .ip1(n326), .ip2(n325), .op(n327) );
  nor4_1 U459 ( .ip1(ipwdata[3]), .ip2(ipwdata[4]), .ip3(ipwdata[7]), .ip4(
        n327), .op(n682) );
  nor4_1 U460 ( .ip1(ipwdata[8]), .ip2(ipwdata[9]), .ip3(ipwdata[10]), .ip4(
        ipwdata[11]), .op(n329) );
  nand3_1 U461 ( .ip1(n682), .ip2(n329), .ip3(n328), .op(n600) );
  or2_1 U462 ( .ip1(ipwdata[2]), .ip2(n600), .op(n331) );
  or2_1 U463 ( .ip1(ipwdata[1]), .ip2(n600), .op(n330) );
  nand2_1 U464 ( .ip1(n331), .ip2(n330), .op(n364) );
  nand2_1 U465 ( .ip1(n533), .ip2(n689), .op(n597) );
  nor2_1 U466 ( .ip1(n364), .ip2(n597), .op(n596) );
  nand2_1 U467 ( .ip1(ipwdata[14]), .ip2(n596), .op(n333) );
  nand2_1 U468 ( .ip1(hcr_ic_ss_hcnt[14]), .ip2(n597), .op(n332) );
  nand2_1 U469 ( .ip1(n333), .ip2(n332), .op(n1497) );
  nand2_1 U470 ( .ip1(ipwdata[13]), .ip2(n596), .op(n335) );
  nand2_1 U471 ( .ip1(hcr_ic_ss_hcnt[13]), .ip2(n597), .op(n334) );
  nand2_1 U472 ( .ip1(n335), .ip2(n334), .op(n1498) );
  nand2_1 U473 ( .ip1(ipwdata[12]), .ip2(n596), .op(n337) );
  nand2_1 U474 ( .ip1(hcr_ic_ss_hcnt[12]), .ip2(n597), .op(n336) );
  nand2_1 U475 ( .ip1(n337), .ip2(n336), .op(n1499) );
  nand2_1 U476 ( .ip1(ipwdata[11]), .ip2(n596), .op(n339) );
  nand2_1 U477 ( .ip1(hcr_ic_ss_hcnt[11]), .ip2(n597), .op(n338) );
  nand2_1 U478 ( .ip1(n339), .ip2(n338), .op(n1500) );
  nand2_1 U479 ( .ip1(ipwdata[10]), .ip2(n596), .op(n341) );
  nand2_1 U480 ( .ip1(hcr_ic_ss_hcnt[10]), .ip2(n597), .op(n340) );
  nand2_1 U481 ( .ip1(n341), .ip2(n340), .op(n1501) );
  nand2_1 U482 ( .ip1(ipwdata[9]), .ip2(n596), .op(n343) );
  nand2_1 U483 ( .ip1(hcr_ic_ss_hcnt[9]), .ip2(n597), .op(n342) );
  nand2_1 U484 ( .ip1(n343), .ip2(n342), .op(n1502) );
  nand2_1 U485 ( .ip1(ipwdata[8]), .ip2(n596), .op(n345) );
  nand2_1 U486 ( .ip1(hcr_ic_ss_hcnt[8]), .ip2(n597), .op(n344) );
  nand2_1 U487 ( .ip1(n345), .ip2(n344), .op(n1503) );
  nand2_1 U488 ( .ip1(ipwdata[15]), .ip2(n596), .op(n347) );
  nand2_1 U489 ( .ip1(hcr_ic_ss_hcnt[15]), .ip2(n597), .op(n346) );
  nand2_1 U490 ( .ip1(n347), .ip2(n346), .op(n1504) );
  nand2_1 U491 ( .ip1(n522), .ip2(n689), .op(n637) );
  mux2_1 U492 ( .ip1(ipwdata[14]), .ip2(hcr_ic_hs_lcnt[14]), .s(n637), .op(
        n1417) );
  mux2_1 U493 ( .ip1(ipwdata[13]), .ip2(hcr_ic_hs_lcnt[13]), .s(n637), .op(
        n1418) );
  mux2_1 U494 ( .ip1(ipwdata[12]), .ip2(hcr_ic_hs_lcnt[12]), .s(n637), .op(
        n1419) );
  mux2_1 U495 ( .ip1(ipwdata[11]), .ip2(hcr_ic_hs_lcnt[11]), .s(n637), .op(
        n1420) );
  mux2_1 U496 ( .ip1(ipwdata[10]), .ip2(hcr_ic_hs_lcnt[10]), .s(n637), .op(
        n1421) );
  mux2_1 U497 ( .ip1(ipwdata[9]), .ip2(hcr_ic_hs_lcnt[9]), .s(n637), .op(n1422) );
  mux2_1 U498 ( .ip1(ipwdata[8]), .ip2(hcr_ic_hs_lcnt[8]), .s(n637), .op(n1423) );
  mux2_1 U499 ( .ip1(ipwdata[15]), .ip2(hcr_ic_hs_lcnt[15]), .s(n637), .op(
        n1424) );
  nand2_1 U500 ( .ip1(n525), .ip2(n689), .op(n630) );
  nor2_1 U501 ( .ip1(n364), .ip2(n630), .op(n629) );
  nand2_1 U502 ( .ip1(ipwdata[14]), .ip2(n629), .op(n349) );
  nand2_1 U503 ( .ip1(hcr_ic_hs_hcnt[14]), .ip2(n630), .op(n348) );
  nand2_1 U504 ( .ip1(n349), .ip2(n348), .op(n1433) );
  nand2_1 U505 ( .ip1(ipwdata[13]), .ip2(n629), .op(n351) );
  nand2_1 U506 ( .ip1(hcr_ic_hs_hcnt[13]), .ip2(n630), .op(n350) );
  nand2_1 U507 ( .ip1(n351), .ip2(n350), .op(n1434) );
  nand2_1 U508 ( .ip1(ipwdata[12]), .ip2(n629), .op(n353) );
  nand2_1 U509 ( .ip1(hcr_ic_hs_hcnt[12]), .ip2(n630), .op(n352) );
  nand2_1 U510 ( .ip1(n353), .ip2(n352), .op(n1435) );
  nand2_1 U511 ( .ip1(ipwdata[11]), .ip2(n629), .op(n355) );
  nand2_1 U512 ( .ip1(hcr_ic_hs_hcnt[11]), .ip2(n630), .op(n354) );
  nand2_1 U513 ( .ip1(n355), .ip2(n354), .op(n1436) );
  nand2_1 U514 ( .ip1(ipwdata[10]), .ip2(n629), .op(n357) );
  nand2_1 U515 ( .ip1(hcr_ic_hs_hcnt[10]), .ip2(n630), .op(n356) );
  nand2_1 U516 ( .ip1(n357), .ip2(n356), .op(n1437) );
  nand2_1 U517 ( .ip1(ipwdata[9]), .ip2(n629), .op(n359) );
  nand2_1 U518 ( .ip1(hcr_ic_hs_hcnt[9]), .ip2(n630), .op(n358) );
  nand2_1 U519 ( .ip1(n359), .ip2(n358), .op(n1438) );
  nand2_1 U520 ( .ip1(ipwdata[8]), .ip2(n629), .op(n361) );
  nand2_1 U521 ( .ip1(hcr_ic_hs_hcnt[8]), .ip2(n630), .op(n360) );
  nand2_1 U522 ( .ip1(n361), .ip2(n360), .op(n1439) );
  nand2_1 U523 ( .ip1(ipwdata[15]), .ip2(n629), .op(n363) );
  nand2_1 U524 ( .ip1(hcr_ic_hs_hcnt[15]), .ip2(n630), .op(n362) );
  nand2_1 U525 ( .ip1(n363), .ip2(n362), .op(n1440) );
  nand2_1 U526 ( .ip1(n523), .ip2(n689), .op(n609) );
  nor2_1 U527 ( .ip1(n364), .ip2(n609), .op(n608) );
  nand2_1 U528 ( .ip1(ipwdata[12]), .ip2(n608), .op(n366) );
  nand2_1 U529 ( .ip1(ic_fs_hcnt[12]), .ip2(n609), .op(n365) );
  nand2_1 U530 ( .ip1(n366), .ip2(n365), .op(n1467) );
  nand2_1 U531 ( .ip1(ipwdata[13]), .ip2(n608), .op(n368) );
  nand2_1 U532 ( .ip1(ic_fs_hcnt[13]), .ip2(n609), .op(n367) );
  nand2_1 U533 ( .ip1(n368), .ip2(n367), .op(n1466) );
  nand2_1 U534 ( .ip1(ipwdata[14]), .ip2(n608), .op(n370) );
  nand2_1 U535 ( .ip1(ic_fs_hcnt[14]), .ip2(n609), .op(n369) );
  nand2_1 U536 ( .ip1(n370), .ip2(n369), .op(n1465) );
  nand2_1 U537 ( .ip1(ipwdata[11]), .ip2(n608), .op(n372) );
  nand2_1 U538 ( .ip1(ic_fs_hcnt[11]), .ip2(n609), .op(n371) );
  nand2_1 U539 ( .ip1(n372), .ip2(n371), .op(n1468) );
  nand2_1 U540 ( .ip1(ipwdata[10]), .ip2(n608), .op(n374) );
  nand2_1 U541 ( .ip1(ic_fs_hcnt[10]), .ip2(n609), .op(n373) );
  nand2_1 U542 ( .ip1(n374), .ip2(n373), .op(n1469) );
  nand2_1 U543 ( .ip1(ipwdata[9]), .ip2(n608), .op(n376) );
  nand2_1 U544 ( .ip1(ic_fs_hcnt[9]), .ip2(n609), .op(n375) );
  nand2_1 U545 ( .ip1(n376), .ip2(n375), .op(n1470) );
  nand2_1 U546 ( .ip1(ipwdata[8]), .ip2(n608), .op(n378) );
  nand2_1 U547 ( .ip1(ic_fs_hcnt[8]), .ip2(n609), .op(n377) );
  nand2_1 U548 ( .ip1(n378), .ip2(n377), .op(n1471) );
  nand2_1 U549 ( .ip1(ipwdata[15]), .ip2(n608), .op(n380) );
  nand2_1 U550 ( .ip1(ic_fs_hcnt[15]), .ip2(n609), .op(n379) );
  nand2_1 U551 ( .ip1(n380), .ip2(n379), .op(n1472) );
  nand2_1 U552 ( .ip1(n532), .ip2(n689), .op(n601) );
  mux2_1 U553 ( .ip1(ipwdata[14]), .ip2(hcr_ic_ss_lcnt[14]), .s(n601), .op(
        n1481) );
  mux2_1 U554 ( .ip1(ipwdata[13]), .ip2(hcr_ic_ss_lcnt[13]), .s(n601), .op(
        n1482) );
  mux2_1 U555 ( .ip1(ipwdata[12]), .ip2(hcr_ic_ss_lcnt[12]), .s(n601), .op(
        n1483) );
  mux2_1 U556 ( .ip1(ipwdata[11]), .ip2(hcr_ic_ss_lcnt[11]), .s(n601), .op(
        n1484) );
  mux2_1 U557 ( .ip1(ipwdata[10]), .ip2(hcr_ic_ss_lcnt[10]), .s(n601), .op(
        n1485) );
  mux2_1 U558 ( .ip1(ipwdata[9]), .ip2(hcr_ic_ss_lcnt[9]), .s(n601), .op(n1486) );
  mux2_1 U559 ( .ip1(ipwdata[8]), .ip2(hcr_ic_ss_lcnt[8]), .s(n601), .op(n1487) );
  mux2_1 U560 ( .ip1(ipwdata[15]), .ip2(hcr_ic_ss_lcnt[15]), .s(n601), .op(
        n1488) );
  nand2_1 U561 ( .ip1(n506), .ip2(wr_en), .op(n651) );
  inv_1 U562 ( .ip(n651), .op(tx_push) );
  inv_1 U563 ( .ip(tx_abrt_flg_edg), .op(n554) );
  nand2_1 U564 ( .ip1(n554), .ip2(ic_enable[0]), .op(n381) );
  nor2_1 U565 ( .ip1(n382), .ip2(n381), .op(fifo_rst_n) );
  inv_1 U566 ( .ip(fifo_rst_n), .op(n559) );
  or2_1 U567 ( .ip1(n383), .ip2(n559), .op(n385) );
  inv_1 U568 ( .ip(fifo_rst_n_int), .op(n649) );
  or2_1 U569 ( .ip1(n649), .ip2(n559), .op(n384) );
  nand2_1 U570 ( .ip1(n385), .ip2(n384), .op(n386) );
  or2_1 U571 ( .ip1(n386), .ip2(n703), .op(fix_c) );
  nand2_1 U572 ( .ip1(n477), .ip2(ic_fs_lcnt[0]), .op(n389) );
  nand2_1 U573 ( .ip1(hcr_ic_ss_lcnt[0]), .ip2(ic_ss), .op(n388) );
  nand2_1 U574 ( .ip1(hcr_ic_hs_lcnt[0]), .ip2(ic_hs), .op(n387) );
  nand3_1 U575 ( .ip1(n389), .ip2(n388), .ip3(n387), .op(ic_lcnt[0]) );
  nand2_1 U576 ( .ip1(n477), .ip2(ic_fs_lcnt[1]), .op(n392) );
  nand2_1 U577 ( .ip1(hcr_ic_hs_lcnt[1]), .ip2(ic_hs), .op(n391) );
  nand2_1 U578 ( .ip1(hcr_ic_ss_lcnt[1]), .ip2(ic_ss), .op(n390) );
  nand3_1 U579 ( .ip1(n392), .ip2(n391), .ip3(n390), .op(ic_lcnt[1]) );
  nand2_1 U580 ( .ip1(n477), .ip2(ic_fs_lcnt[2]), .op(n395) );
  nand2_1 U581 ( .ip1(hcr_ic_hs_lcnt[2]), .ip2(ic_hs), .op(n394) );
  nand2_1 U582 ( .ip1(hcr_ic_ss_lcnt[2]), .ip2(ic_ss), .op(n393) );
  nand3_1 U583 ( .ip1(n395), .ip2(n394), .ip3(n393), .op(ic_lcnt[2]) );
  nand2_1 U584 ( .ip1(n477), .ip2(ic_fs_lcnt[3]), .op(n398) );
  nand2_1 U585 ( .ip1(hcr_ic_hs_lcnt[3]), .ip2(ic_hs), .op(n397) );
  nand2_1 U586 ( .ip1(hcr_ic_ss_lcnt[3]), .ip2(ic_ss), .op(n396) );
  nand3_1 U587 ( .ip1(n398), .ip2(n397), .ip3(n396), .op(ic_lcnt[3]) );
  nand2_1 U588 ( .ip1(n477), .ip2(ic_fs_lcnt[4]), .op(n401) );
  nand2_1 U589 ( .ip1(hcr_ic_hs_lcnt[4]), .ip2(ic_hs), .op(n400) );
  nand2_1 U590 ( .ip1(hcr_ic_ss_lcnt[4]), .ip2(ic_ss), .op(n399) );
  nand3_1 U591 ( .ip1(n401), .ip2(n400), .ip3(n399), .op(ic_lcnt[4]) );
  nand2_1 U592 ( .ip1(n477), .ip2(ic_fs_lcnt[5]), .op(n404) );
  nand2_1 U593 ( .ip1(hcr_ic_hs_lcnt[5]), .ip2(ic_hs), .op(n403) );
  nand2_1 U594 ( .ip1(hcr_ic_ss_lcnt[5]), .ip2(ic_ss), .op(n402) );
  nand3_1 U595 ( .ip1(n404), .ip2(n403), .ip3(n402), .op(ic_lcnt[5]) );
  nand2_1 U596 ( .ip1(n477), .ip2(ic_fs_lcnt[6]), .op(n407) );
  nand2_1 U597 ( .ip1(hcr_ic_hs_lcnt[6]), .ip2(ic_hs), .op(n406) );
  nand2_1 U598 ( .ip1(hcr_ic_ss_lcnt[6]), .ip2(ic_ss), .op(n405) );
  nand3_1 U599 ( .ip1(n407), .ip2(n406), .ip3(n405), .op(ic_lcnt[6]) );
  nand2_1 U600 ( .ip1(n477), .ip2(ic_fs_lcnt[7]), .op(n410) );
  nand2_1 U601 ( .ip1(hcr_ic_hs_lcnt[7]), .ip2(ic_hs), .op(n409) );
  nand2_1 U602 ( .ip1(hcr_ic_ss_lcnt[7]), .ip2(ic_ss), .op(n408) );
  nand3_1 U603 ( .ip1(n410), .ip2(n409), .ip3(n408), .op(ic_lcnt[7]) );
  nand2_1 U604 ( .ip1(n477), .ip2(ic_fs_lcnt[8]), .op(n413) );
  nand2_1 U605 ( .ip1(hcr_ic_hs_lcnt[8]), .ip2(ic_hs), .op(n412) );
  nand2_1 U606 ( .ip1(hcr_ic_ss_lcnt[8]), .ip2(ic_ss), .op(n411) );
  nand3_1 U607 ( .ip1(n413), .ip2(n412), .ip3(n411), .op(ic_lcnt[8]) );
  nand2_1 U608 ( .ip1(n477), .ip2(ic_fs_lcnt[9]), .op(n416) );
  nand2_1 U609 ( .ip1(hcr_ic_hs_lcnt[9]), .ip2(ic_hs), .op(n415) );
  nand2_1 U610 ( .ip1(hcr_ic_ss_lcnt[9]), .ip2(ic_ss), .op(n414) );
  nand3_1 U611 ( .ip1(n416), .ip2(n415), .ip3(n414), .op(ic_lcnt[9]) );
  nand2_1 U612 ( .ip1(n477), .ip2(ic_fs_lcnt[10]), .op(n419) );
  nand2_1 U613 ( .ip1(hcr_ic_hs_lcnt[10]), .ip2(ic_hs), .op(n418) );
  nand2_1 U614 ( .ip1(hcr_ic_ss_lcnt[10]), .ip2(ic_ss), .op(n417) );
  nand3_1 U615 ( .ip1(n419), .ip2(n418), .ip3(n417), .op(ic_lcnt[10]) );
  nand2_1 U616 ( .ip1(n477), .ip2(ic_fs_lcnt[11]), .op(n422) );
  nand2_1 U617 ( .ip1(hcr_ic_hs_lcnt[11]), .ip2(ic_hs), .op(n421) );
  nand2_1 U618 ( .ip1(hcr_ic_ss_lcnt[11]), .ip2(ic_ss), .op(n420) );
  nand3_1 U619 ( .ip1(n422), .ip2(n421), .ip3(n420), .op(ic_lcnt[11]) );
  nand2_1 U620 ( .ip1(n477), .ip2(ic_fs_lcnt[12]), .op(n425) );
  nand2_1 U621 ( .ip1(hcr_ic_hs_lcnt[12]), .ip2(ic_hs), .op(n424) );
  nand2_1 U622 ( .ip1(hcr_ic_ss_lcnt[12]), .ip2(ic_ss), .op(n423) );
  nand3_1 U623 ( .ip1(n425), .ip2(n424), .ip3(n423), .op(ic_lcnt[12]) );
  nand2_1 U624 ( .ip1(n477), .ip2(ic_fs_lcnt[13]), .op(n428) );
  nand2_1 U625 ( .ip1(hcr_ic_hs_lcnt[13]), .ip2(ic_hs), .op(n427) );
  nand2_1 U626 ( .ip1(hcr_ic_ss_lcnt[13]), .ip2(ic_ss), .op(n426) );
  nand3_1 U627 ( .ip1(n428), .ip2(n427), .ip3(n426), .op(ic_lcnt[13]) );
  nand2_1 U628 ( .ip1(n477), .ip2(ic_fs_lcnt[14]), .op(n431) );
  nand2_1 U629 ( .ip1(hcr_ic_hs_lcnt[14]), .ip2(ic_hs), .op(n430) );
  nand2_1 U630 ( .ip1(hcr_ic_ss_lcnt[14]), .ip2(ic_ss), .op(n429) );
  nand3_1 U631 ( .ip1(n431), .ip2(n430), .ip3(n429), .op(ic_lcnt[14]) );
  nand2_1 U632 ( .ip1(n477), .ip2(ic_fs_lcnt[15]), .op(n434) );
  nand2_1 U633 ( .ip1(hcr_ic_hs_lcnt[15]), .ip2(ic_hs), .op(n433) );
  nand2_1 U634 ( .ip1(hcr_ic_ss_lcnt[15]), .ip2(ic_ss), .op(n432) );
  nand3_1 U635 ( .ip1(n434), .ip2(n433), .ip3(n432), .op(ic_lcnt[15]) );
  nand2_1 U636 ( .ip1(hcr_ic_hs_hcnt[0]), .ip2(ic_hs), .op(n437) );
  nand2_1 U637 ( .ip1(ic_fs_hcnt[0]), .ip2(n477), .op(n436) );
  nand2_1 U638 ( .ip1(hcr_ic_ss_hcnt[0]), .ip2(ic_ss), .op(n435) );
  nand3_1 U639 ( .ip1(n437), .ip2(n436), .ip3(n435), .op(ic_hcnt[0]) );
  nand2_1 U640 ( .ip1(n477), .ip2(ic_fs_hcnt[2]), .op(n440) );
  nand2_1 U641 ( .ip1(hcr_ic_hs_hcnt[2]), .ip2(ic_hs), .op(n439) );
  nand2_1 U642 ( .ip1(hcr_ic_ss_hcnt[2]), .ip2(ic_ss), .op(n438) );
  nand3_1 U643 ( .ip1(n440), .ip2(n439), .ip3(n438), .op(ic_hcnt[2]) );
  nand2_1 U644 ( .ip1(n477), .ip2(ic_fs_hcnt[3]), .op(n443) );
  nand2_1 U645 ( .ip1(hcr_ic_hs_hcnt[3]), .ip2(ic_hs), .op(n442) );
  nand2_1 U646 ( .ip1(hcr_ic_ss_hcnt[3]), .ip2(ic_ss), .op(n441) );
  nand3_1 U647 ( .ip1(n443), .ip2(n442), .ip3(n441), .op(ic_hcnt[3]) );
  nand2_1 U648 ( .ip1(n477), .ip2(ic_fs_hcnt[4]), .op(n446) );
  nand2_1 U649 ( .ip1(hcr_ic_hs_hcnt[4]), .ip2(ic_hs), .op(n445) );
  nand2_1 U650 ( .ip1(hcr_ic_ss_hcnt[4]), .ip2(ic_ss), .op(n444) );
  nand3_1 U651 ( .ip1(n446), .ip2(n445), .ip3(n444), .op(ic_hcnt[4]) );
  nand2_1 U652 ( .ip1(n477), .ip2(ic_fs_hcnt[5]), .op(n449) );
  nand2_1 U653 ( .ip1(hcr_ic_hs_hcnt[5]), .ip2(ic_hs), .op(n448) );
  nand2_1 U654 ( .ip1(hcr_ic_ss_hcnt[5]), .ip2(ic_ss), .op(n447) );
  nand3_1 U655 ( .ip1(n449), .ip2(n448), .ip3(n447), .op(ic_hcnt[5]) );
  nand2_1 U656 ( .ip1(n477), .ip2(ic_fs_hcnt[6]), .op(n452) );
  nand2_1 U657 ( .ip1(hcr_ic_hs_hcnt[6]), .ip2(ic_hs), .op(n451) );
  nand2_1 U658 ( .ip1(hcr_ic_ss_hcnt[6]), .ip2(ic_ss), .op(n450) );
  nand3_1 U659 ( .ip1(n452), .ip2(n451), .ip3(n450), .op(ic_hcnt[6]) );
  nand2_1 U660 ( .ip1(n477), .ip2(ic_fs_hcnt[7]), .op(n455) );
  nand2_1 U661 ( .ip1(hcr_ic_hs_hcnt[7]), .ip2(ic_hs), .op(n454) );
  nand2_1 U662 ( .ip1(hcr_ic_ss_hcnt[7]), .ip2(ic_ss), .op(n453) );
  nand3_1 U663 ( .ip1(n455), .ip2(n454), .ip3(n453), .op(ic_hcnt[7]) );
  nand2_1 U664 ( .ip1(n477), .ip2(ic_fs_hcnt[8]), .op(n458) );
  nand2_1 U665 ( .ip1(hcr_ic_hs_hcnt[8]), .ip2(ic_hs), .op(n457) );
  nand2_1 U666 ( .ip1(hcr_ic_ss_hcnt[8]), .ip2(ic_ss), .op(n456) );
  nand3_1 U667 ( .ip1(n458), .ip2(n457), .ip3(n456), .op(ic_hcnt[8]) );
  nand2_1 U668 ( .ip1(n477), .ip2(ic_fs_hcnt[9]), .op(n461) );
  nand2_1 U669 ( .ip1(hcr_ic_hs_hcnt[9]), .ip2(ic_hs), .op(n460) );
  nand2_1 U670 ( .ip1(hcr_ic_ss_hcnt[9]), .ip2(ic_ss), .op(n459) );
  nand3_1 U671 ( .ip1(n461), .ip2(n460), .ip3(n459), .op(ic_hcnt[9]) );
  nand2_1 U672 ( .ip1(n477), .ip2(ic_fs_hcnt[10]), .op(n464) );
  nand2_1 U673 ( .ip1(hcr_ic_hs_hcnt[10]), .ip2(ic_hs), .op(n463) );
  nand2_1 U674 ( .ip1(hcr_ic_ss_hcnt[10]), .ip2(ic_ss), .op(n462) );
  nand3_1 U675 ( .ip1(n464), .ip2(n463), .ip3(n462), .op(ic_hcnt[10]) );
  nand2_1 U676 ( .ip1(n477), .ip2(ic_fs_hcnt[11]), .op(n467) );
  nand2_1 U677 ( .ip1(hcr_ic_hs_hcnt[11]), .ip2(ic_hs), .op(n466) );
  nand2_1 U678 ( .ip1(hcr_ic_ss_hcnt[11]), .ip2(ic_ss), .op(n465) );
  nand3_1 U679 ( .ip1(n467), .ip2(n466), .ip3(n465), .op(ic_hcnt[11]) );
  nand2_1 U680 ( .ip1(n477), .ip2(ic_fs_hcnt[12]), .op(n470) );
  nand2_1 U681 ( .ip1(hcr_ic_hs_hcnt[12]), .ip2(ic_hs), .op(n469) );
  nand2_1 U682 ( .ip1(hcr_ic_ss_hcnt[12]), .ip2(ic_ss), .op(n468) );
  nand3_1 U683 ( .ip1(n470), .ip2(n469), .ip3(n468), .op(ic_hcnt[12]) );
  nand2_1 U684 ( .ip1(n477), .ip2(ic_fs_hcnt[13]), .op(n473) );
  nand2_1 U685 ( .ip1(hcr_ic_hs_hcnt[13]), .ip2(ic_hs), .op(n472) );
  nand2_1 U686 ( .ip1(hcr_ic_ss_hcnt[13]), .ip2(ic_ss), .op(n471) );
  nand3_1 U687 ( .ip1(n473), .ip2(n472), .ip3(n471), .op(ic_hcnt[13]) );
  nand2_1 U688 ( .ip1(n477), .ip2(ic_fs_hcnt[14]), .op(n476) );
  nand2_1 U689 ( .ip1(hcr_ic_hs_hcnt[14]), .ip2(ic_hs), .op(n475) );
  nand2_1 U690 ( .ip1(hcr_ic_ss_hcnt[14]), .ip2(ic_ss), .op(n474) );
  nand3_1 U691 ( .ip1(n476), .ip2(n475), .ip3(n474), .op(ic_hcnt[14]) );
  nand2_1 U692 ( .ip1(n477), .ip2(ic_fs_hcnt[15]), .op(n480) );
  nand2_1 U693 ( .ip1(hcr_ic_hs_hcnt[15]), .ip2(ic_hs), .op(n479) );
  nand2_1 U694 ( .ip1(hcr_ic_ss_hcnt[15]), .ip2(ic_ss), .op(n478) );
  nand3_1 U695 ( .ip1(n480), .ip2(n479), .ip3(n478), .op(ic_hcnt[15]) );
  nand2_1 U696 ( .ip1(n523), .ip2(ic_fs_hcnt[3]), .op(n483) );
  nand2_1 U697 ( .ip1(n532), .ip2(hcr_ic_ss_lcnt[3]), .op(n482) );
  nand2_1 U698 ( .ip1(n646), .ip2(ic_sda_hold[3]), .op(n481) );
  nand3_1 U699 ( .ip1(n483), .ip2(n482), .ip3(n481), .op(n512) );
  nor2_1 U700 ( .ip1(rx_empty), .ip2(n484), .op(n493) );
  nand2_1 U701 ( .ip1(ic_raw_intr_stat[3]), .ip2(n485), .op(n491) );
  nand2_1 U702 ( .ip1(n486), .ip2(ic_rxflr[3]), .op(n490) );
  nand2_1 U703 ( .ip1(n487), .ip2(ic_txflr[3]), .op(n489) );
  nand2_1 U704 ( .ip1(n533), .ip2(hcr_ic_ss_hcnt[3]), .op(n488) );
  nand4_1 U705 ( .ip1(n491), .ip2(n490), .ip3(n489), .ip4(n488), .op(n492) );
  not_ab_or_c_or_d U706 ( .ip1(hcr_ic_hs_lcnt[3]), .ip2(n522), .ip3(n493), 
        .ip4(n492), .op(n510) );
  nand2_1 U707 ( .ip1(n587), .ip2(ic_tar[3]), .op(n497) );
  nand2_1 U708 ( .ip1(n638), .ip2(ic_fs_spklen[3]), .op(n496) );
  nand2_1 U709 ( .ip1(n582), .ip2(ic_10bit_slv), .op(n495) );
  nand2_1 U710 ( .ip1(n524), .ip2(ic_fs_lcnt[3]), .op(n494) );
  nand4_1 U711 ( .ip1(n497), .ip2(n496), .ip3(n495), .ip4(n494), .op(n505) );
  not_ab_or_c_or_d U712 ( .ip1(n499), .ip2(ic_intr_stat[3]), .ip3(iprdata[29]), 
        .ip4(n498), .op(n503) );
  nand2_1 U713 ( .ip1(n525), .ip2(hcr_ic_hs_hcnt[3]), .op(n502) );
  nand2_1 U714 ( .ip1(n690), .ip2(ic_sda_setup[3]), .op(n501) );
  nand2_1 U715 ( .ip1(n644), .ip2(ic_intr_mask[3]), .op(n500) );
  nand4_1 U716 ( .ip1(n503), .ip2(n502), .ip3(n501), .ip4(n500), .op(n504) );
  not_ab_or_c_or_d U717 ( .ip1(n549), .ip2(ic_tx_abrt_source[3]), .ip3(n505), 
        .ip4(n504), .op(n509) );
  nand2_1 U718 ( .ip1(n506), .ip2(rx_pop_data[3]), .op(n508) );
  nand2_1 U719 ( .ip1(n586), .ip2(ic_sar[3]), .op(n507) );
  nand4_1 U720 ( .ip1(n510), .ip2(n509), .ip3(n508), .ip4(n507), .op(n511) );
  ab_or_c_or_d U721 ( .ip1(n641), .ip2(ic_hs_spklen[3]), .ip3(n512), .ip4(n511), .op(iprdata[3]) );
  inv_1 U722 ( .ip(ic_con_pre_6_), .op(ic_slave_en) );
  nand2_1 U723 ( .ip1(n522), .ip2(hcr_ic_hs_lcnt[14]), .op(n521) );
  and2_1 U724 ( .ip1(n523), .ip2(ic_fs_hcnt[14]), .op(n518) );
  nand2_1 U725 ( .ip1(n524), .ip2(ic_fs_lcnt[14]), .op(n516) );
  nand2_1 U726 ( .ip1(n646), .ip2(ic_sda_hold[14]), .op(n515) );
  nand2_1 U727 ( .ip1(n549), .ip2(ic_tx_abrt_source[14]), .op(n514) );
  nand2_1 U728 ( .ip1(n525), .ip2(hcr_ic_hs_hcnt[14]), .op(n513) );
  nand4_1 U729 ( .ip1(n516), .ip2(n515), .ip3(n514), .ip4(n513), .op(n517) );
  not_ab_or_c_or_d U730 ( .ip1(n532), .ip2(hcr_ic_ss_lcnt[14]), .ip3(n518), 
        .ip4(n517), .op(n520) );
  nand2_1 U731 ( .ip1(n533), .ip2(hcr_ic_ss_hcnt[14]), .op(n519) );
  nand3_1 U732 ( .ip1(n521), .ip2(n520), .ip3(n519), .op(iprdata[14]) );
  nand2_1 U733 ( .ip1(n522), .ip2(hcr_ic_hs_lcnt[15]), .op(n536) );
  and2_1 U734 ( .ip1(n523), .ip2(ic_fs_hcnt[15]), .op(n531) );
  nand2_1 U735 ( .ip1(n524), .ip2(ic_fs_lcnt[15]), .op(n529) );
  nand2_1 U736 ( .ip1(n646), .ip2(ic_sda_hold[15]), .op(n528) );
  nand2_1 U737 ( .ip1(n549), .ip2(ic_tx_abrt_source[15]), .op(n527) );
  nand2_1 U738 ( .ip1(n525), .ip2(hcr_ic_hs_hcnt[15]), .op(n526) );
  nand4_1 U739 ( .ip1(n529), .ip2(n528), .ip3(n527), .ip4(n526), .op(n530) );
  not_ab_or_c_or_d U740 ( .ip1(n532), .ip2(hcr_ic_ss_lcnt[15]), .ip3(n531), 
        .ip4(n530), .op(n535) );
  nand2_1 U741 ( .ip1(n533), .ip2(hcr_ic_ss_hcnt[15]), .op(n534) );
  nand3_1 U742 ( .ip1(n536), .ip2(n535), .ip3(n534), .op(iprdata[15]) );
  nand2_1 U743 ( .ip1(ic_tx_abrt_source[16]), .ip2(n549), .op(n538) );
  nand2_1 U744 ( .ip1(n646), .ip2(ic_sda_hold[16]), .op(n537) );
  nand3_1 U745 ( .ip1(n538), .ip2(n541), .ip3(n537), .op(iprdata[16]) );
  nand2_1 U746 ( .ip1(ic_sda_hold[17]), .ip2(n646), .op(n539) );
  nand3_1 U747 ( .ip1(n539), .ip2(n541), .ip3(n548), .op(iprdata[17]) );
  nand2_1 U748 ( .ip1(n646), .ip2(ic_sda_hold[18]), .op(n540) );
  nand2_1 U749 ( .ip1(n541), .ip2(n540), .op(iprdata[18]) );
  and2_1 U750 ( .ip1(n646), .ip2(ic_sda_hold[19]), .op(iprdata[19]) );
  nand2_1 U751 ( .ip1(ic_sda_hold[20]), .ip2(n646), .op(n542) );
  inv_1 U752 ( .ip(iprdata[30]), .op(n551) );
  nand3_1 U753 ( .ip1(n542), .ip2(n551), .ip3(n548), .op(iprdata[20]) );
  nand2_1 U754 ( .ip1(n646), .ip2(ic_sda_hold[21]), .op(n543) );
  nand2_1 U755 ( .ip1(n548), .ip2(n543), .op(iprdata[21]) );
  nand2_1 U756 ( .ip1(n646), .ip2(ic_sda_hold[22]), .op(n544) );
  nand2_1 U757 ( .ip1(n551), .ip2(n544), .op(iprdata[22]) );
  nand2_1 U758 ( .ip1(ic_sda_hold[23]), .ip2(n646), .op(n546) );
  nand2_1 U759 ( .ip1(ic_txflr_flushed[0]), .ip2(n549), .op(n545) );
  nand2_1 U760 ( .ip1(n546), .ip2(n545), .op(iprdata[23]) );
  nand2_1 U761 ( .ip1(n549), .ip2(ic_txflr_flushed[1]), .op(n547) );
  nand2_1 U762 ( .ip1(n548), .ip2(n547), .op(iprdata[24]) );
  and2_1 U763 ( .ip1(n549), .ip2(ic_txflr_flushed[2]), .op(iprdata[25]) );
  nand2_1 U764 ( .ip1(n549), .ip2(ic_txflr_flushed[3]), .op(n550) );
  nand2_1 U765 ( .ip1(n551), .ip2(n550), .op(iprdata[26]) );
  nor2_1 U766 ( .ip1(ic_con_pre_1_), .ip2(n552), .op(ic_fs) );
  nor3_1 U767 ( .ip1(n703), .ip2(n553), .ip3(n680), .op(n555) );
  mux2_1 U768 ( .ip1(n555), .ip2(n554), .s(ic_enable[1]), .op(n1548) );
  inv_1 U769 ( .ip(ic_rxflr[1]), .op(n557) );
  inv_1 U770 ( .ip(rx_push_sync), .op(n556) );
  nor4_1 U771 ( .ip1(n559), .ip2(n556), .ip3(ic_rxflr[3]), .ip4(rx_pop), .op(
        n562) );
  nand2_1 U772 ( .ip1(ic_rxflr[0]), .ip2(n562), .op(n574) );
  nor2_1 U773 ( .ip1(n557), .ip2(n574), .op(n578) );
  nand2_1 U774 ( .ip1(ic_rxflr[2]), .ip2(n578), .op(n569) );
  nor4_1 U775 ( .ip1(ic_rxflr[0]), .ip2(ic_rxflr[3]), .ip3(ic_rxflr[1]), .ip4(
        ic_rxflr[2]), .op(n560) );
  nor4_1 U776 ( .ip1(rx_push_sync), .ip2(n560), .ip3(n559), .ip4(n558), .op(
        n565) );
  inv_1 U777 ( .ip(n562), .op(n561) );
  nor2_1 U778 ( .ip1(n561), .ip2(ic_rxflr[1]), .op(n564) );
  inv_1 U779 ( .ip(n565), .op(n573) );
  mux2_1 U780 ( .ip1(n561), .ip2(n573), .s(ic_rxflr[0]), .op(n563) );
  nor2_1 U781 ( .ip1(n565), .ip2(n562), .op(n571) );
  nand2_1 U782 ( .ip1(fifo_rst_n), .ip2(n571), .op(n570) );
  nand2_1 U783 ( .ip1(n563), .ip2(n570), .op(n576) );
  not_ab_or_c_or_d U784 ( .ip1(ic_rxflr[1]), .ip2(n565), .ip3(n564), .ip4(n576), .op(n579) );
  nand2_1 U785 ( .ip1(ic_rxflr[2]), .ip2(n565), .op(n566) );
  nand2_1 U786 ( .ip1(n579), .ip2(n566), .op(n567) );
  nand2_1 U787 ( .ip1(ic_rxflr[3]), .ip2(n567), .op(n568) );
  nand2_1 U788 ( .ip1(n569), .ip2(n568), .op(n1547) );
  mux2_1 U789 ( .ip1(n571), .ip2(n570), .s(ic_rxflr[0]), .op(n572) );
  inv_1 U790 ( .ip(n572), .op(n1546) );
  nor3_1 U791 ( .ip1(ic_rxflr[0]), .ip2(ic_rxflr[1]), .ip3(n573), .op(n577) );
  nor2_1 U792 ( .ip1(ic_rxflr[1]), .ip2(n574), .op(n575) );
  ab_or_c_or_d U793 ( .ip1(ic_rxflr[1]), .ip2(n576), .ip3(n577), .ip4(n575), 
        .op(n1545) );
  or2_1 U794 ( .ip1(n578), .ip2(n577), .op(n581) );
  inv_1 U795 ( .ip(n579), .op(n580) );
  mux2_1 U796 ( .ip1(n581), .ip2(n580), .s(ic_rxflr[2]), .op(n1544) );
  nand2_1 U797 ( .ip1(n582), .ip2(n689), .op(n585) );
  mux2_1 U798 ( .ip1(ipwdata[8]), .ip2(tx_empty_ctrl), .s(n585), .op(n1543) );
  mux2_1 U799 ( .ip1(ipwdata[7]), .ip2(p_det_ifaddr), .s(n585), .op(n1542) );
  mux2_1 U800 ( .ip1(ipwdata[6]), .ip2(ic_con_pre_6_), .s(n585), .op(n1541) );
  mux2_1 U801 ( .ip1(ipwdata[5]), .ip2(ic_rstrt_en), .s(n585), .op(n1540) );
  mux2_1 U802 ( .ip1(ipwdata[4]), .ip2(ic_10bit_mst), .s(n585), .op(n1539) );
  mux2_1 U803 ( .ip1(ipwdata[3]), .ip2(ic_10bit_slv), .s(n585), .op(n1538) );
  inv_1 U804 ( .ip(ipwdata[2]), .op(n678) );
  nand2_1 U805 ( .ip1(ipwdata[1]), .ip2(n678), .op(n583) );
  mux2_1 U806 ( .ip1(n583), .ip2(ic_con_pre_2_), .s(n585), .op(n1537) );
  nand2_1 U807 ( .ip1(ipwdata[2]), .ip2(n680), .op(n584) );
  mux2_1 U808 ( .ip1(n584), .ip2(ic_con_pre_1_), .s(n585), .op(n1536) );
  mux2_1 U809 ( .ip1(ipwdata[0]), .ip2(ic_master), .s(n585), .op(n1535) );
  nand2_1 U810 ( .ip1(n586), .ip2(n689), .op(n588) );
  mux2_1 U811 ( .ip1(ipwdata[8]), .ip2(ic_sar[8]), .s(n588), .op(n1534) );
  mux2_1 U812 ( .ip1(ipwdata[9]), .ip2(ic_sar[9]), .s(n588), .op(n1533) );
  nand2_1 U813 ( .ip1(n587), .ip2(n689), .op(n589) );
  mux2_1 U814 ( .ip1(ipwdata[8]), .ip2(ic_tar[8]), .s(n589), .op(n1532) );
  mux2_1 U815 ( .ip1(ipwdata[9]), .ip2(ic_tar[9]), .s(n589), .op(n1531) );
  mux2_1 U816 ( .ip1(ipwdata[10]), .ip2(ic_tar[10]), .s(n589), .op(n1530) );
  mux2_1 U817 ( .ip1(ipwdata[11]), .ip2(ic_tar[11]), .s(n589), .op(n1529) );
  mux2_1 U818 ( .ip1(ipwdata[0]), .ip2(ic_sar[0]), .s(n588), .op(n1528) );
  mux2_1 U819 ( .ip1(ipwdata[1]), .ip2(ic_sar[1]), .s(n588), .op(n1527) );
  mux2_1 U820 ( .ip1(ipwdata[2]), .ip2(ic_sar[2]), .s(n588), .op(n1526) );
  mux2_1 U821 ( .ip1(ipwdata[3]), .ip2(ic_sar[3]), .s(n588), .op(n1525) );
  mux2_1 U822 ( .ip1(ipwdata[4]), .ip2(ic_sar[4]), .s(n588), .op(n1524) );
  mux2_1 U823 ( .ip1(ipwdata[5]), .ip2(ic_sar[5]), .s(n588), .op(n1523) );
  mux2_1 U824 ( .ip1(ipwdata[6]), .ip2(ic_sar[6]), .s(n588), .op(n1522) );
  mux2_1 U825 ( .ip1(ipwdata[7]), .ip2(ic_sar[7]), .s(n588), .op(n1521) );
  mux2_1 U826 ( .ip1(ipwdata[0]), .ip2(ic_tar[0]), .s(n589), .op(n1520) );
  mux2_1 U827 ( .ip1(ipwdata[1]), .ip2(ic_tar[1]), .s(n589), .op(n1519) );
  mux2_1 U828 ( .ip1(ipwdata[2]), .ip2(ic_tar[2]), .s(n589), .op(n1518) );
  mux2_1 U829 ( .ip1(ipwdata[3]), .ip2(ic_tar[3]), .s(n589), .op(n1517) );
  mux2_1 U830 ( .ip1(ipwdata[4]), .ip2(ic_tar[4]), .s(n589), .op(n1516) );
  mux2_1 U831 ( .ip1(ipwdata[5]), .ip2(ic_tar[5]), .s(n589), .op(n1515) );
  mux2_1 U832 ( .ip1(ipwdata[6]), .ip2(ic_tar[6]), .s(n589), .op(n1514) );
  mux2_1 U833 ( .ip1(ipwdata[7]), .ip2(ic_tar[7]), .s(n589), .op(n1513) );
  nand2_1 U834 ( .ip1(ipwdata[0]), .ip2(n596), .op(n591) );
  nand2_1 U835 ( .ip1(hcr_ic_ss_hcnt[0]), .ip2(n597), .op(n590) );
  nand2_1 U836 ( .ip1(n591), .ip2(n590), .op(n1512) );
  inv_1 U837 ( .ip(ipwdata[1]), .op(n680) );
  nand2_1 U838 ( .ip1(n600), .ip2(n680), .op(n623) );
  mux2_1 U839 ( .ip1(n623), .ip2(hcr_ic_ss_hcnt[1]), .s(n597), .op(n1511) );
  nand2_1 U840 ( .ip1(n600), .ip2(n678), .op(n624) );
  mux2_1 U841 ( .ip1(n624), .ip2(hcr_ic_ss_hcnt[2]), .s(n597), .op(n1510) );
  nand2_1 U842 ( .ip1(ipwdata[3]), .ip2(n596), .op(n593) );
  nand2_1 U843 ( .ip1(hcr_ic_ss_hcnt[3]), .ip2(n597), .op(n592) );
  nand2_1 U844 ( .ip1(n593), .ip2(n592), .op(n1509) );
  nand2_1 U845 ( .ip1(ipwdata[4]), .ip2(n596), .op(n595) );
  nand2_1 U846 ( .ip1(hcr_ic_ss_hcnt[4]), .ip2(n597), .op(n594) );
  nand2_1 U847 ( .ip1(n595), .ip2(n594), .op(n1508) );
  mux2_1 U848 ( .ip1(ipwdata[5]), .ip2(hcr_ic_ss_hcnt[5]), .s(n597), .op(n1507) );
  mux2_1 U849 ( .ip1(ipwdata[6]), .ip2(hcr_ic_ss_hcnt[6]), .s(n597), .op(n1506) );
  nand2_1 U850 ( .ip1(ipwdata[7]), .ip2(n596), .op(n599) );
  nand2_1 U851 ( .ip1(hcr_ic_ss_hcnt[7]), .ip2(n597), .op(n598) );
  nand2_1 U852 ( .ip1(n599), .ip2(n598), .op(n1505) );
  inv_1 U853 ( .ip(n600), .op(n612) );
  nor2_1 U854 ( .ip1(n612), .ip2(n681), .op(n633) );
  mux2_1 U855 ( .ip1(n633), .ip2(hcr_ic_ss_lcnt[0]), .s(n601), .op(n1496) );
  nor2_1 U856 ( .ip1(n612), .ip2(n680), .op(n634) );
  mux2_1 U857 ( .ip1(n634), .ip2(hcr_ic_ss_lcnt[1]), .s(n601), .op(n1495) );
  nor2_1 U858 ( .ip1(n612), .ip2(n678), .op(n635) );
  mux2_1 U859 ( .ip1(n635), .ip2(hcr_ic_ss_lcnt[2]), .s(n601), .op(n1494) );
  or2_1 U860 ( .ip1(ipwdata[3]), .ip2(n612), .op(n636) );
  mux2_1 U861 ( .ip1(n636), .ip2(hcr_ic_ss_lcnt[3]), .s(n601), .op(n1493) );
  mux2_1 U862 ( .ip1(ipwdata[4]), .ip2(hcr_ic_ss_lcnt[4]), .s(n601), .op(n1492) );
  mux2_1 U863 ( .ip1(ipwdata[5]), .ip2(hcr_ic_ss_lcnt[5]), .s(n601), .op(n1491) );
  mux2_1 U864 ( .ip1(ipwdata[6]), .ip2(hcr_ic_ss_lcnt[6]), .s(n601), .op(n1490) );
  mux2_1 U865 ( .ip1(ipwdata[7]), .ip2(hcr_ic_ss_lcnt[7]), .s(n601), .op(n1489) );
  nand2_1 U866 ( .ip1(ipwdata[0]), .ip2(n608), .op(n603) );
  nand2_1 U867 ( .ip1(ic_fs_hcnt[0]), .ip2(n609), .op(n602) );
  nand2_1 U868 ( .ip1(n603), .ip2(n602), .op(n1480) );
  mux2_1 U869 ( .ip1(n623), .ip2(ic_fs_hcnt[1]), .s(n609), .op(n1479) );
  mux2_1 U870 ( .ip1(n624), .ip2(ic_fs_hcnt[2]), .s(n609), .op(n1478) );
  nand2_1 U871 ( .ip1(ipwdata[3]), .ip2(n608), .op(n605) );
  nand2_1 U872 ( .ip1(ic_fs_hcnt[3]), .ip2(n609), .op(n604) );
  nand2_1 U873 ( .ip1(n605), .ip2(n604), .op(n1477) );
  nand2_1 U874 ( .ip1(ipwdata[4]), .ip2(n608), .op(n607) );
  nand2_1 U875 ( .ip1(ic_fs_hcnt[4]), .ip2(n609), .op(n606) );
  nand2_1 U876 ( .ip1(n607), .ip2(n606), .op(n1476) );
  mux2_1 U877 ( .ip1(ipwdata[5]), .ip2(ic_fs_hcnt[5]), .s(n609), .op(n1475) );
  mux2_1 U878 ( .ip1(ipwdata[6]), .ip2(ic_fs_hcnt[6]), .s(n609), .op(n1474) );
  nand2_1 U879 ( .ip1(ipwdata[7]), .ip2(n608), .op(n611) );
  nand2_1 U880 ( .ip1(ic_fs_hcnt[7]), .ip2(n609), .op(n610) );
  nand2_1 U881 ( .ip1(n611), .ip2(n610), .op(n1473) );
  nor2_1 U882 ( .ip1(n612), .ip2(n620), .op(n617) );
  nand2_1 U883 ( .ip1(ipwdata[0]), .ip2(n617), .op(n614) );
  nand2_1 U884 ( .ip1(ic_fs_lcnt[0]), .ip2(n620), .op(n613) );
  nand2_1 U885 ( .ip1(n614), .ip2(n613), .op(n1464) );
  nand2_1 U886 ( .ip1(n617), .ip2(ipwdata[1]), .op(n616) );
  nand2_1 U887 ( .ip1(ic_fs_lcnt[1]), .ip2(n620), .op(n615) );
  nand2_1 U888 ( .ip1(n616), .ip2(n615), .op(n1463) );
  nand2_1 U889 ( .ip1(n617), .ip2(ipwdata[2]), .op(n619) );
  nand2_1 U890 ( .ip1(ic_fs_lcnt[2]), .ip2(n620), .op(n618) );
  nand2_1 U891 ( .ip1(n619), .ip2(n618), .op(n1462) );
  mux2_1 U892 ( .ip1(n636), .ip2(ic_fs_lcnt[3]), .s(n620), .op(n1461) );
  mux2_1 U893 ( .ip1(ipwdata[4]), .ip2(ic_fs_lcnt[4]), .s(n620), .op(n1460) );
  mux2_1 U894 ( .ip1(ipwdata[5]), .ip2(ic_fs_lcnt[5]), .s(n620), .op(n1459) );
  mux2_1 U895 ( .ip1(ipwdata[6]), .ip2(ic_fs_lcnt[6]), .s(n620), .op(n1458) );
  mux2_1 U896 ( .ip1(ipwdata[7]), .ip2(ic_fs_lcnt[7]), .s(n620), .op(n1457) );
  nand2_1 U897 ( .ip1(ipwdata[0]), .ip2(n629), .op(n622) );
  nand2_1 U898 ( .ip1(hcr_ic_hs_hcnt[0]), .ip2(n630), .op(n621) );
  nand2_1 U899 ( .ip1(n622), .ip2(n621), .op(n1448) );
  mux2_1 U900 ( .ip1(n623), .ip2(hcr_ic_hs_hcnt[1]), .s(n630), .op(n1447) );
  mux2_1 U901 ( .ip1(n624), .ip2(hcr_ic_hs_hcnt[2]), .s(n630), .op(n1446) );
  nand2_1 U902 ( .ip1(ipwdata[3]), .ip2(n629), .op(n626) );
  nand2_1 U903 ( .ip1(hcr_ic_hs_hcnt[3]), .ip2(n630), .op(n625) );
  nand2_1 U904 ( .ip1(n626), .ip2(n625), .op(n1445) );
  nand2_1 U905 ( .ip1(ipwdata[4]), .ip2(n629), .op(n628) );
  nand2_1 U906 ( .ip1(hcr_ic_hs_hcnt[4]), .ip2(n630), .op(n627) );
  nand2_1 U907 ( .ip1(n628), .ip2(n627), .op(n1444) );
  mux2_1 U908 ( .ip1(ipwdata[5]), .ip2(hcr_ic_hs_hcnt[5]), .s(n630), .op(n1443) );
  mux2_1 U909 ( .ip1(ipwdata[6]), .ip2(hcr_ic_hs_hcnt[6]), .s(n630), .op(n1442) );
  nand2_1 U910 ( .ip1(ipwdata[7]), .ip2(n629), .op(n632) );
  nand2_1 U911 ( .ip1(hcr_ic_hs_hcnt[7]), .ip2(n630), .op(n631) );
  nand2_1 U912 ( .ip1(n632), .ip2(n631), .op(n1441) );
  mux2_1 U913 ( .ip1(n633), .ip2(hcr_ic_hs_lcnt[0]), .s(n637), .op(n1432) );
  mux2_1 U914 ( .ip1(n634), .ip2(hcr_ic_hs_lcnt[1]), .s(n637), .op(n1431) );
  mux2_1 U915 ( .ip1(n635), .ip2(hcr_ic_hs_lcnt[2]), .s(n637), .op(n1430) );
  mux2_1 U916 ( .ip1(n636), .ip2(hcr_ic_hs_lcnt[3]), .s(n637), .op(n1429) );
  mux2_1 U917 ( .ip1(ipwdata[4]), .ip2(hcr_ic_hs_lcnt[4]), .s(n637), .op(n1428) );
  mux2_1 U918 ( .ip1(ipwdata[5]), .ip2(hcr_ic_hs_lcnt[5]), .s(n637), .op(n1427) );
  mux2_1 U919 ( .ip1(ipwdata[6]), .ip2(hcr_ic_hs_lcnt[6]), .s(n637), .op(n1426) );
  mux2_1 U920 ( .ip1(ipwdata[7]), .ip2(hcr_ic_hs_lcnt[7]), .s(n637), .op(n1425) );
  nand2_1 U921 ( .ip1(n638), .ip2(n689), .op(n640) );
  mux2_1 U922 ( .ip1(ipwdata[7]), .ip2(ic_fs_spklen[7]), .s(n640), .op(n1416)
         );
  mux2_1 U923 ( .ip1(ipwdata[6]), .ip2(ic_fs_spklen[6]), .s(n640), .op(n1415)
         );
  mux2_1 U924 ( .ip1(ipwdata[5]), .ip2(ic_fs_spklen[5]), .s(n640), .op(n1414)
         );
  mux2_1 U925 ( .ip1(ipwdata[4]), .ip2(ic_fs_spklen[4]), .s(n640), .op(n1413)
         );
  mux2_1 U926 ( .ip1(ipwdata[3]), .ip2(ic_fs_spklen[3]), .s(n640), .op(n1412)
         );
  mux2_1 U927 ( .ip1(ipwdata[2]), .ip2(ic_fs_spklen[2]), .s(n640), .op(n1411)
         );
  mux2_1 U928 ( .ip1(ipwdata[1]), .ip2(ic_fs_spklen[1]), .s(n640), .op(n1410)
         );
  nand3_1 U929 ( .ip1(n678), .ip2(n682), .ip3(n680), .op(n639) );
  inv_1 U930 ( .ip(ipwdata[0]), .op(n681) );
  nand2_1 U931 ( .ip1(n639), .ip2(n681), .op(n643) );
  mux2_1 U932 ( .ip1(n643), .ip2(ic_fs_spklen[0]), .s(n640), .op(n1409) );
  nand2_1 U933 ( .ip1(n641), .ip2(n689), .op(n642) );
  mux2_1 U934 ( .ip1(ipwdata[7]), .ip2(ic_hs_spklen[7]), .s(n642), .op(n1408)
         );
  mux2_1 U935 ( .ip1(ipwdata[6]), .ip2(ic_hs_spklen[6]), .s(n642), .op(n1407)
         );
  mux2_1 U936 ( .ip1(ipwdata[5]), .ip2(ic_hs_spklen[5]), .s(n642), .op(n1406)
         );
  mux2_1 U937 ( .ip1(ipwdata[4]), .ip2(ic_hs_spklen[4]), .s(n642), .op(n1405)
         );
  mux2_1 U938 ( .ip1(ipwdata[3]), .ip2(ic_hs_spklen[3]), .s(n642), .op(n1404)
         );
  mux2_1 U939 ( .ip1(ipwdata[2]), .ip2(ic_hs_spklen[2]), .s(n642), .op(n1403)
         );
  mux2_1 U940 ( .ip1(ipwdata[1]), .ip2(ic_hs_spklen[1]), .s(n642), .op(n1402)
         );
  mux2_1 U941 ( .ip1(n643), .ip2(ic_hs_spklen[0]), .s(n642), .op(n1401) );
  and2_1 U942 ( .ip1(n644), .ip2(wr_en), .op(n645) );
  mux2_1 U943 ( .ip1(ic_intr_mask[8]), .ip2(ipwdata[8]), .s(n645), .op(n1400)
         );
  mux2_1 U944 ( .ip1(ic_intr_mask[9]), .ip2(ipwdata[9]), .s(n645), .op(n1399)
         );
  mux2_1 U945 ( .ip1(ic_intr_mask[10]), .ip2(ipwdata[10]), .s(n645), .op(n1398) );
  mux2_1 U946 ( .ip1(ic_intr_mask[11]), .ip2(ipwdata[11]), .s(n645), .op(n1397) );
  mux2_1 U947 ( .ip1(ic_intr_mask[0]), .ip2(ipwdata[0]), .s(n645), .op(n1396)
         );
  mux2_1 U948 ( .ip1(ic_intr_mask[1]), .ip2(ipwdata[1]), .s(n645), .op(n1395)
         );
  mux2_1 U949 ( .ip1(ic_intr_mask[2]), .ip2(ipwdata[2]), .s(n645), .op(n1394)
         );
  mux2_1 U950 ( .ip1(ic_intr_mask[3]), .ip2(ipwdata[3]), .s(n645), .op(n1393)
         );
  mux2_1 U951 ( .ip1(ic_intr_mask[4]), .ip2(ipwdata[4]), .s(n645), .op(n1392)
         );
  mux2_1 U952 ( .ip1(ic_intr_mask[5]), .ip2(ipwdata[5]), .s(n645), .op(n1391)
         );
  mux2_1 U953 ( .ip1(ic_intr_mask[6]), .ip2(ipwdata[6]), .s(n645), .op(n1390)
         );
  mux2_1 U954 ( .ip1(ic_intr_mask[7]), .ip2(ipwdata[7]), .s(n645), .op(n1389)
         );
  nand2_1 U955 ( .ip1(n646), .ip2(n689), .op(n647) );
  mux2_1 U956 ( .ip1(ipwdata[23]), .ip2(ic_sda_hold[23]), .s(n647), .op(n1388)
         );
  mux2_1 U957 ( .ip1(ipwdata[22]), .ip2(ic_sda_hold[22]), .s(n648), .op(n1387)
         );
  mux2_1 U958 ( .ip1(ipwdata[21]), .ip2(ic_sda_hold[21]), .s(n648), .op(n1386)
         );
  mux2_1 U959 ( .ip1(ipwdata[20]), .ip2(ic_sda_hold[20]), .s(n647), .op(n1385)
         );
  mux2_1 U960 ( .ip1(ipwdata[19]), .ip2(ic_sda_hold[19]), .s(n648), .op(n1384)
         );
  mux2_1 U961 ( .ip1(ipwdata[18]), .ip2(ic_sda_hold[18]), .s(n648), .op(n1383)
         );
  mux2_1 U962 ( .ip1(ipwdata[17]), .ip2(ic_sda_hold[17]), .s(n647), .op(n1382)
         );
  mux2_1 U963 ( .ip1(ipwdata[16]), .ip2(ic_sda_hold[16]), .s(n648), .op(n1381)
         );
  mux2_1 U964 ( .ip1(ipwdata[15]), .ip2(ic_sda_hold[15]), .s(n648), .op(n1380)
         );
  mux2_1 U965 ( .ip1(ipwdata[14]), .ip2(ic_sda_hold[14]), .s(n648), .op(n1379)
         );
  mux2_1 U966 ( .ip1(ipwdata[13]), .ip2(ic_sda_hold[13]), .s(n648), .op(n1378)
         );
  mux2_1 U967 ( .ip1(ipwdata[12]), .ip2(ic_sda_hold[12]), .s(n647), .op(n1377)
         );
  mux2_1 U968 ( .ip1(ipwdata[11]), .ip2(ic_sda_hold[11]), .s(n647), .op(n1376)
         );
  mux2_1 U969 ( .ip1(ipwdata[10]), .ip2(ic_sda_hold[10]), .s(n648), .op(n1375)
         );
  mux2_1 U970 ( .ip1(ipwdata[9]), .ip2(ic_sda_hold[9]), .s(n648), .op(n1374)
         );
  mux2_1 U971 ( .ip1(ipwdata[8]), .ip2(ic_sda_hold[8]), .s(n648), .op(n1373)
         );
  mux2_1 U972 ( .ip1(ipwdata[7]), .ip2(ic_sda_hold[7]), .s(n648), .op(n1372)
         );
  mux2_1 U973 ( .ip1(ipwdata[6]), .ip2(ic_sda_hold[6]), .s(n648), .op(n1371)
         );
  mux2_1 U974 ( .ip1(ipwdata[5]), .ip2(ic_sda_hold[5]), .s(n648), .op(n1370)
         );
  mux2_1 U975 ( .ip1(ipwdata[4]), .ip2(ic_sda_hold[4]), .s(n648), .op(n1369)
         );
  mux2_1 U976 ( .ip1(ipwdata[3]), .ip2(ic_sda_hold[3]), .s(n648), .op(n1368)
         );
  mux2_1 U977 ( .ip1(ipwdata[2]), .ip2(ic_sda_hold[2]), .s(n648), .op(n1367)
         );
  mux2_1 U978 ( .ip1(ipwdata[1]), .ip2(ic_sda_hold[1]), .s(n648), .op(n1366)
         );
  mux2_1 U979 ( .ip1(ipwdata[0]), .ip2(ic_sda_hold[0]), .s(n648), .op(n1365)
         );
  nor3_1 U980 ( .ip1(slv_clr_leftover_flg_edg), .ip2(n703), .ip3(n649), .op(
        tx_fifo_rst_n) );
  inv_1 U981 ( .ip(tx_fifo_rst_n), .op(n652) );
  nor3_1 U982 ( .ip1(ic_txflr[0]), .ip2(ic_txflr[1]), .ip3(ic_txflr[2]), .op(
        n675) );
  inv_1 U983 ( .ip(ic_txflr[3]), .op(n698) );
  nand2_1 U984 ( .ip1(tx_fifo_rst_n), .ip2(tx_pop_sync), .op(n650) );
  not_ab_or_c_or_d U985 ( .ip1(n675), .ip2(n698), .ip3(tx_push), .ip4(n650), 
        .op(n676) );
  inv_1 U986 ( .ip(n676), .op(n653) );
  nor4_1 U987 ( .ip1(n652), .ip2(n651), .ip3(ic_txflr[3]), .ip4(tx_pop_sync), 
        .op(n663) );
  inv_1 U988 ( .ip(n663), .op(n672) );
  nand2_1 U989 ( .ip1(n653), .ip2(n672), .op(n659) );
  nor2_1 U990 ( .ip1(n652), .ip2(n659), .op(n660) );
  nor2_1 U991 ( .ip1(n653), .ip2(n675), .op(n654) );
  or2_1 U992 ( .ip1(n660), .ip2(n654), .op(n655) );
  nand2_1 U993 ( .ip1(ic_txflr[3]), .ip2(n655), .op(n658) );
  nand3_1 U994 ( .ip1(ic_txflr[0]), .ip2(ic_txflr[1]), .ip3(ic_txflr[2]), .op(
        n656) );
  mux2_1 U995 ( .ip1(ic_txflr[3]), .ip2(n698), .s(n656), .op(n697) );
  or2_1 U996 ( .ip1(n672), .ip2(n697), .op(n657) );
  nand2_1 U997 ( .ip1(n658), .ip2(n657), .op(n1364) );
  inv_1 U998 ( .ip(ic_txflr[0]), .op(n691) );
  mux2_1 U999 ( .ip1(n660), .ip2(n659), .s(n691), .op(n1363) );
  mux2_1 U1000 ( .ip1(n663), .ip2(n676), .s(n691), .op(n666) );
  or2_1 U1001 ( .ip1(n676), .ip2(n660), .op(n662) );
  or2_1 U1002 ( .ip1(ic_txflr[0]), .ip2(n660), .op(n661) );
  nand2_1 U1003 ( .ip1(n662), .ip2(n661), .op(n667) );
  nand2_1 U1004 ( .ip1(n663), .ip2(n691), .op(n664) );
  nand2_1 U1005 ( .ip1(n667), .ip2(n664), .op(n665) );
  mux2_1 U1006 ( .ip1(n666), .ip2(n665), .s(ic_txflr[1]), .op(n1362) );
  inv_1 U1007 ( .ip(ic_txflr[2]), .op(n702) );
  or2_1 U1008 ( .ip1(n667), .ip2(n702), .op(n670) );
  nand2_1 U1009 ( .ip1(ic_txflr[1]), .ip2(n676), .op(n668) );
  or2_1 U1010 ( .ip1(n668), .ip2(n702), .op(n669) );
  nand2_1 U1011 ( .ip1(n670), .ip2(n669), .op(n674) );
  nand2_1 U1012 ( .ip1(ic_txflr[0]), .ip2(ic_txflr[1]), .op(n671) );
  mux2_1 U1013 ( .ip1(ic_txflr[2]), .ip2(n702), .s(n671), .op(n701) );
  nor2_1 U1014 ( .ip1(n672), .ip2(n701), .op(n673) );
  ab_or_c_or_d U1015 ( .ip1(n676), .ip2(n675), .ip3(n674), .ip4(n673), .op(
        n1361) );
  nand2_1 U1016 ( .ip1(n677), .ip2(n689), .op(n706) );
  mux2_1 U1017 ( .ip1(ipwdata[2]), .ip2(ic_hs_maddr[2]), .s(n706), .op(n1167)
         );
  mux2_1 U1018 ( .ip1(ipwdata[1]), .ip2(ic_hs_maddr[1]), .s(n706), .op(n1165)
         );
  nand2_1 U1019 ( .ip1(n682), .ip2(n678), .op(n685) );
  nand2_1 U1020 ( .ip1(n679), .ip2(wr_en), .op(n683) );
  mux2_1 U1021 ( .ip1(n685), .ip2(ic_rx_tl_int[2]), .s(n683), .op(n1153) );
  nand2_1 U1022 ( .ip1(n682), .ip2(n680), .op(n686) );
  mux2_1 U1023 ( .ip1(n686), .ip2(ic_rx_tl_int[1]), .s(n683), .op(n1151) );
  nand2_1 U1024 ( .ip1(n682), .ip2(n681), .op(n688) );
  mux2_1 U1025 ( .ip1(n688), .ip2(ic_rx_tl_int[0]), .s(n683), .op(n1149) );
  and2_1 U1026 ( .ip1(n684), .ip2(wr_en), .op(n687) );
  mux2_1 U1027 ( .ip1(ic_tx_tl_2_), .ip2(n685), .s(n687), .op(n1137) );
  mux2_1 U1028 ( .ip1(ic_tx_tl_1_), .ip2(n686), .s(n687), .op(n1135) );
  mux2_1 U1029 ( .ip1(ic_tx_tl_0_), .ip2(n688), .s(n687), .op(n1133) );
  nand2_1 U1030 ( .ip1(n690), .ip2(n689), .op(n707) );
  mux2_1 U1031 ( .ip1(ipwdata[7]), .ip2(ic_sda_setup[7]), .s(n707), .op(n1131)
         );
  mux2_1 U1032 ( .ip1(ipwdata[4]), .ip2(ic_sda_setup[4]), .s(n707), .op(n1129)
         );
  mux2_1 U1033 ( .ip1(ipwdata[3]), .ip2(ic_sda_setup[3]), .s(n707), .op(n1127)
         );
  mux2_1 U1034 ( .ip1(ipwdata[1]), .ip2(ic_sda_setup[1]), .s(n707), .op(n1125)
         );
  mux2_1 U1035 ( .ip1(ipwdata[0]), .ip2(ic_sda_setup[0]), .s(n707), .op(n1123)
         );
  mux2_1 U1036 ( .ip1(n691), .ip2(ic_txflr[0]), .s(abrt_in_rcve_trns), .op(
        n693) );
  nor2_1 U1037 ( .ip1(ic_txflr_flushed[0]), .ip2(tx_abrt_flg_edg), .op(n692)
         );
  not_ab_or_c_or_d U1038 ( .ip1(tx_abrt_flg_edg), .ip2(n693), .ip3(n692), 
        .ip4(n703), .op(n1121) );
  nand2_1 U1039 ( .ip1(abrt_in_rcve_trns), .ip2(ic_txflr[0]), .op(n694) );
  xor2_1 U1040 ( .ip1(ic_txflr[1]), .ip2(n694), .op(n696) );
  nor2_1 U1041 ( .ip1(ic_txflr_flushed[1]), .ip2(tx_abrt_flg_edg), .op(n695)
         );
  not_ab_or_c_or_d U1042 ( .ip1(tx_abrt_flg_edg), .ip2(n696), .ip3(n695), 
        .ip4(n703), .op(n1119) );
  mux2_1 U1043 ( .ip1(n698), .ip2(n697), .s(abrt_in_rcve_trns), .op(n700) );
  nor2_1 U1044 ( .ip1(ic_txflr_flushed[3]), .ip2(tx_abrt_flg_edg), .op(n699)
         );
  not_ab_or_c_or_d U1045 ( .ip1(tx_abrt_flg_edg), .ip2(n700), .ip3(n699), 
        .ip4(n703), .op(n1117) );
  mux2_1 U1046 ( .ip1(n702), .ip2(n701), .s(abrt_in_rcve_trns), .op(n705) );
  nor2_1 U1047 ( .ip1(ic_txflr_flushed[2]), .ip2(tx_abrt_flg_edg), .op(n704)
         );
  not_ab_or_c_or_d U1048 ( .ip1(tx_abrt_flg_edg), .ip2(n705), .ip3(n704), 
        .ip4(n703), .op(n1115) );
  mux2_1 U1049 ( .ip1(ipwdata[0]), .ip2(ic_hs_maddr[0]), .s(n706), .op(n1113)
         );
  mux2_1 U1050 ( .ip1(ipwdata[6]), .ip2(ic_sda_setup[6]), .s(n707), .op(n1111)
         );
  mux2_1 U1051 ( .ip1(ipwdata[5]), .ip2(ic_sda_setup[5]), .s(n707), .op(n1109)
         );
  mux2_1 U1052 ( .ip1(ipwdata[2]), .ip2(ic_sda_setup[2]), .s(n707), .op(n1107)
         );
  nand2_1 U1053 ( .ip1(n708), .ip2(wr_en), .op(n709) );
  mux2_1 U1054 ( .ip1(ipwdata[0]), .ip2(ic_ack_general_call), .s(n709), .op(
        n1105) );
endmodule


module interconnect_ip ( HCLK_hclk, HRESETn_hresetn, PCLK_pclk, 
        PRESETn_presetn, ex_i_ahb_AHB_MASTER_CORTEXM0_haddr, 
        ex_i_ahb_AHB_MASTER_CORTEXM0_hburst, 
        ex_i_ahb_AHB_MASTER_CORTEXM0_hlock, ex_i_ahb_AHB_MASTER_CORTEXM0_hprot, 
        ex_i_ahb_AHB_MASTER_CORTEXM0_hsize, 
        ex_i_ahb_AHB_MASTER_CORTEXM0_htrans, 
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata, 
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite, 
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata, 
        ex_i_ahb_AHB_MASTER_CORTEXM0_hready, 
        ex_i_ahb_AHB_MASTER_CORTEXM0_hresp, ex_i_ahb_AHB_Slave_PID_hrdata, 
        ex_i_ahb_AHB_Slave_PID_hready_resp, ex_i_ahb_AHB_Slave_PID_hresp, 
        ex_i_ahb_AHB_Slave_PID_haddr, ex_i_ahb_AHB_Slave_PID_hburst, 
        ex_i_ahb_AHB_Slave_PID_hmastlock, ex_i_ahb_AHB_Slave_PID_hprot, 
        ex_i_ahb_AHB_Slave_PID_hready, ex_i_ahb_AHB_Slave_PID_hsel, 
        ex_i_ahb_AHB_Slave_PID_hsize, ex_i_ahb_AHB_Slave_PID_htrans, 
        ex_i_ahb_AHB_Slave_PID_hwdata, ex_i_ahb_AHB_Slave_PID_hwrite, 
        ex_i_ahb_AHB_Slave_PWM_hrdata, ex_i_ahb_AHB_Slave_PWM_hready_resp, 
        ex_i_ahb_AHB_Slave_PWM_hresp, ex_i_ahb_AHB_Slave_PWM_haddr, 
        ex_i_ahb_AHB_Slave_PWM_hburst, ex_i_ahb_AHB_Slave_PWM_hmastlock, 
        ex_i_ahb_AHB_Slave_PWM_hprot, ex_i_ahb_AHB_Slave_PWM_hready, 
        ex_i_ahb_AHB_Slave_PWM_hsel, ex_i_ahb_AHB_Slave_PWM_hsize, 
        ex_i_ahb_AHB_Slave_PWM_htrans, ex_i_ahb_AHB_Slave_PWM_hwdata, 
        ex_i_ahb_AHB_Slave_PWM_hwrite, ex_i_ahb_AHB_Slave_RAM_hrdata, 
        ex_i_ahb_AHB_Slave_RAM_hready_resp, ex_i_ahb_AHB_Slave_RAM_hresp, 
        ex_i_ahb_AHB_Slave_RAM_haddr, ex_i_ahb_AHB_Slave_RAM_hburst, 
        ex_i_ahb_AHB_Slave_RAM_hmastlock, ex_i_ahb_AHB_Slave_RAM_hprot, 
        ex_i_ahb_AHB_Slave_RAM_hready, ex_i_ahb_AHB_Slave_RAM_hsel, 
        ex_i_ahb_AHB_Slave_RAM_hsize, ex_i_ahb_AHB_Slave_RAM_htrans, 
        ex_i_ahb_AHB_Slave_RAM_hwdata, ex_i_ahb_AHB_Slave_RAM_hwrite, 
        i_apb_pclk_en, i_i2c_ic_clk, i_i2c_ic_clk_in_a, i_i2c_ic_data_in_a, 
        i_i2c_ic_rst_n, i_ssi_rxd, i_ssi_ss_in_n, i_ssi_ssi_clk, 
        i_ssi_ssi_rst_n, i_ahb_hmaster_data, i_i2c_debug_addr, 
        i_i2c_debug_addr_10bit, i_i2c_debug_data, i_i2c_debug_hs, 
        i_i2c_debug_master_act, i_i2c_debug_mst_cstate, i_i2c_debug_p_gen, 
        i_i2c_debug_rd, i_i2c_debug_s_gen, i_i2c_debug_slave_act, 
        i_i2c_debug_slv_cstate, i_i2c_debug_wr, i_i2c_ic_activity_intr, 
        i_i2c_ic_clk_oe, i_i2c_ic_current_src_en, i_i2c_ic_data_oe, 
        i_i2c_ic_en, i_i2c_ic_gen_call_intr, i_i2c_ic_rd_req_intr, 
        i_i2c_ic_rx_done_intr, i_i2c_ic_rx_full_intr, i_i2c_ic_rx_over_intr, 
        i_i2c_ic_rx_under_intr, i_i2c_ic_start_det_intr, 
        i_i2c_ic_stop_det_intr, i_i2c_ic_tx_abrt_intr, i_i2c_ic_tx_empty_intr, 
        i_i2c_ic_tx_over_intr, i_ssi_sclk_out, i_ssi_ss_0_n, 
        i_ssi_ssi_mst_intr_n, i_ssi_ssi_oe_n, i_ssi_ssi_rxf_intr_n, 
        i_ssi_ssi_rxo_intr_n, i_ssi_ssi_rxu_intr_n, i_ssi_ssi_sleep, 
        i_ssi_ssi_txe_intr_n, i_ssi_ssi_txo_intr_n, i_ssi_txd );
  input [31:0] ex_i_ahb_AHB_MASTER_CORTEXM0_haddr;
  input [2:0] ex_i_ahb_AHB_MASTER_CORTEXM0_hburst;
  input [3:0] ex_i_ahb_AHB_MASTER_CORTEXM0_hprot;
  input [2:0] ex_i_ahb_AHB_MASTER_CORTEXM0_hsize;
  input [1:0] ex_i_ahb_AHB_MASTER_CORTEXM0_htrans;
  input [31:0] ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata;
  output [31:0] ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata;
  output [1:0] ex_i_ahb_AHB_MASTER_CORTEXM0_hresp;
  input [31:0] ex_i_ahb_AHB_Slave_PID_hrdata;
  input [1:0] ex_i_ahb_AHB_Slave_PID_hresp;
  output [31:0] ex_i_ahb_AHB_Slave_PID_haddr;
  output [2:0] ex_i_ahb_AHB_Slave_PID_hburst;
  output [3:0] ex_i_ahb_AHB_Slave_PID_hprot;
  output [2:0] ex_i_ahb_AHB_Slave_PID_hsize;
  output [1:0] ex_i_ahb_AHB_Slave_PID_htrans;
  output [31:0] ex_i_ahb_AHB_Slave_PID_hwdata;
  input [31:0] ex_i_ahb_AHB_Slave_PWM_hrdata;
  input [1:0] ex_i_ahb_AHB_Slave_PWM_hresp;
  output [31:0] ex_i_ahb_AHB_Slave_PWM_haddr;
  output [2:0] ex_i_ahb_AHB_Slave_PWM_hburst;
  output [3:0] ex_i_ahb_AHB_Slave_PWM_hprot;
  output [2:0] ex_i_ahb_AHB_Slave_PWM_hsize;
  output [1:0] ex_i_ahb_AHB_Slave_PWM_htrans;
  output [31:0] ex_i_ahb_AHB_Slave_PWM_hwdata;
  input [31:0] ex_i_ahb_AHB_Slave_RAM_hrdata;
  input [1:0] ex_i_ahb_AHB_Slave_RAM_hresp;
  output [31:0] ex_i_ahb_AHB_Slave_RAM_haddr;
  output [2:0] ex_i_ahb_AHB_Slave_RAM_hburst;
  output [3:0] ex_i_ahb_AHB_Slave_RAM_hprot;
  output [2:0] ex_i_ahb_AHB_Slave_RAM_hsize;
  output [1:0] ex_i_ahb_AHB_Slave_RAM_htrans;
  output [31:0] ex_i_ahb_AHB_Slave_RAM_hwdata;
  output [3:0] i_ahb_hmaster_data;
  output [4:0] i_i2c_debug_mst_cstate;
  output [3:0] i_i2c_debug_slv_cstate;
  input HCLK_hclk, HRESETn_hresetn, PCLK_pclk, PRESETn_presetn,
         ex_i_ahb_AHB_MASTER_CORTEXM0_hlock,
         ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite,
         ex_i_ahb_AHB_Slave_PID_hready_resp,
         ex_i_ahb_AHB_Slave_PWM_hready_resp,
         ex_i_ahb_AHB_Slave_RAM_hready_resp, i_apb_pclk_en, i_i2c_ic_clk,
         i_i2c_ic_clk_in_a, i_i2c_ic_data_in_a, i_i2c_ic_rst_n, i_ssi_rxd,
         i_ssi_ss_in_n, i_ssi_ssi_clk, i_ssi_ssi_rst_n;
  output ex_i_ahb_AHB_MASTER_CORTEXM0_hready, ex_i_ahb_AHB_Slave_PID_hmastlock,
         ex_i_ahb_AHB_Slave_PID_hready, ex_i_ahb_AHB_Slave_PID_hsel,
         ex_i_ahb_AHB_Slave_PID_hwrite, ex_i_ahb_AHB_Slave_PWM_hmastlock,
         ex_i_ahb_AHB_Slave_PWM_hready, ex_i_ahb_AHB_Slave_PWM_hsel,
         ex_i_ahb_AHB_Slave_PWM_hwrite, ex_i_ahb_AHB_Slave_RAM_hmastlock,
         ex_i_ahb_AHB_Slave_RAM_hready, ex_i_ahb_AHB_Slave_RAM_hsel,
         ex_i_ahb_AHB_Slave_RAM_hwrite, i_i2c_debug_addr,
         i_i2c_debug_addr_10bit, i_i2c_debug_data, i_i2c_debug_hs,
         i_i2c_debug_master_act, i_i2c_debug_p_gen, i_i2c_debug_rd,
         i_i2c_debug_s_gen, i_i2c_debug_slave_act, i_i2c_debug_wr,
         i_i2c_ic_activity_intr, i_i2c_ic_clk_oe, i_i2c_ic_current_src_en,
         i_i2c_ic_data_oe, i_i2c_ic_en, i_i2c_ic_gen_call_intr,
         i_i2c_ic_rd_req_intr, i_i2c_ic_rx_done_intr, i_i2c_ic_rx_full_intr,
         i_i2c_ic_rx_over_intr, i_i2c_ic_rx_under_intr,
         i_i2c_ic_start_det_intr, i_i2c_ic_stop_det_intr,
         i_i2c_ic_tx_abrt_intr, i_i2c_ic_tx_empty_intr, i_i2c_ic_tx_over_intr,
         i_ssi_sclk_out, i_ssi_ss_0_n, i_ssi_ssi_mst_intr_n, i_ssi_ssi_oe_n,
         i_ssi_ssi_rxf_intr_n, i_ssi_ssi_rxo_intr_n, i_ssi_ssi_rxu_intr_n,
         i_ssi_ssi_sleep, i_ssi_ssi_txe_intr_n, i_ssi_ssi_txo_intr_n,
         i_ssi_txd;
  wire   ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite, ex_i_ahb_AHB_Slave_PID_hmastlock,
         i_apb_hready_resp, i_apb_penable, i_apb_pwrite, i_ahb_hresp_none_0_,
         i_apb_psel_en, i_i2c_tx_full, i_i2c_rx_full, i_i2c_tx_push,
         i_i2c_rx_pop, i_i2c_rx_push_sync, i_i2c_tx_pop_sync,
         i_i2c_tx_fifo_rst_n, i_i2c_fifo_rst_n, i_i2c_abrt_in_rcve_trns,
         i_i2c_split_start_en, i_i2c_ack_det, i_i2c_ic_bus_idle,
         i_i2c_slv_addressed, i_i2c_slv_ack_det, i_i2c_p_det, i_i2c_wr_en,
         i_i2c_sda_vld, i_i2c_slv_rx_2addr, i_i2c_rx_hs_mcode,
         i_i2c_rx_addr_match, i_i2c_slv_rxbyte_rdy, i_i2c_rx_slv_read,
         i_i2c_mst_rxbyte_rdy, i_i2c_slv_rx_ack_vld, i_i2c_mst_rx_bwen,
         i_i2c_rx_scl_hcnt_en, i_i2c_rx_scl_lcnt_en, i_i2c_mst_rx_data_scl,
         i_i2c_mst_rx_ack_vld, i_i2c_slv_tx_ack_vld, i_i2c_mst_tx_ack_vld,
         i_i2c_scl_p_setup_cmplt, i_i2c_scl_s_setup_cmplt,
         i_i2c_scl_s_hld_cmplt, i_i2c_scl_lcnt_cmplt, i_i2c_scl_p_setup_en,
         i_i2c_scl_s_setup_en, i_i2c_scl_hcnt_en, i_i2c_slv_tx_cmplt,
         i_i2c_slv_tx_ready_unconn, i_i2c_scl_hld_low_en, i_i2c_byte_wait_scl,
         i_i2c_slv_fifo_filled_and_flushed_sync, i_i2c_slv_rx_aborted_sync,
         i_i2c_activity, i_i2c_slv_activity_sync, i_i2c_mst_activity_sync,
         i_i2c_tx_abrt_flg_edg, i_i2c_ic_clr_gen_call_en,
         i_i2c_ic_clr_start_det_en, i_i2c_ic_clr_stop_det_en,
         i_i2c_ic_clr_activity_en, i_i2c_ic_clr_rx_done_en,
         i_i2c_ic_clr_tx_abrt_en, i_i2c_ic_clr_rd_req_en,
         i_i2c_ic_clr_tx_over_en, i_i2c_ic_clr_rx_over_en,
         i_i2c_ic_clr_rx_under_en, i_i2c_ic_clr_intr_en, i_i2c_tx_empty_ctrl,
         i_i2c_slv_fifo_filled_and_flushed, i_i2c_slv_rx_aborted,
         i_i2c_ic_ack_general_call_sync, i_i2c_ic_slave_en_sync,
         i_i2c_p_det_ifaddr_sync, i_i2c_ic_ss_sync, i_i2c_ic_fs_sync,
         i_i2c_ic_abort_sync, i_i2c_ic_ack_general_call, i_i2c_p_det_ifaddr,
         i_i2c_ic_slave_en, i_i2c_ic_rstrt_en, i_i2c_ic_10bit_slv, i_i2c_ic_ss,
         i_i2c_ic_fs, i_i2c_ic_hs, i_i2c_ic_10bit_mst, i_i2c_ic_master,
         i_i2c_set_tx_empty_en_flg, i_i2c_slv_clr_leftover_flg,
         i_i2c_rx_push_flg, i_i2c_tx_pop_flg, i_i2c_rx_gen_call_flg,
         i_i2c_s_det_flg, i_i2c_p_det_flg, i_i2c_ic_rd_req_flg,
         i_i2c_rx_done_flg, i_i2c_tx_abrt_flg, i_i2c_rx_addr_10bit,
         i_i2c_hs_mcode_en, i_i2c_ic_enable_sync, i_i2c_re_start_en,
         i_i2c_start_en, i_i2c_rx_current_src_en, i_i2c_tx_current_src_en,
         i_i2c_set_tx_empty_en, i_i2c_rx_push, i_i2c_tx_pop, i_i2c_rx_gen_call,
         i_i2c_s_det, i_i2c_p_det_intr, i_i2c_slv_activity, i_i2c_mst_activity,
         i_ssi_mst_contention, i_ssi_load_start_bit, i_ssi_rx_push,
         i_ssi_tx_pop, i_ssi_sclk_fe, i_ssi_sclk_re, i_ssi_start_xfer,
         i_ssi_baud2, i_ssi_ser_0_, i_ssi_sclk_active, i_ssi_fsm_multi_mst,
         i_ssi_ssi_en_int, i_ssi_rx_full, i_ssi_tx_full, i_ssi_tx_pop_sync,
         i_ssi_fsm_busy, i_ssi_fsm_sleep, i_ahb_U_dfltslv_N4,
         i_ahb_U_dfltslv_next_state, i_ahb_U_dfltslv_current_state,
         i_apb_U_DW_apb_ahbsif_N727, i_apb_U_DW_apb_ahbsif_use_saved_c,
         i_apb_U_DW_apb_ahbsif_piped_hwrite_c,
         i_apb_U_DW_apb_ahbsif_pipeline_c,
         i_apb_U_DW_apb_ahbsif_use_saved_data, i_i2c_U_DW_apb_i2c_toggle_N33,
         i_i2c_U_DW_apb_i2c_toggle_N32, i_i2c_U_DW_apb_i2c_toggle_N31,
         i_i2c_U_DW_apb_i2c_toggle_N30, i_i2c_U_DW_apb_i2c_toggle_N29,
         i_i2c_U_DW_apb_i2c_toggle_rx_gen_call_r,
         i_i2c_U_DW_apb_i2c_toggle_tx_abrt_r,
         i_i2c_U_DW_apb_i2c_toggle_tx_abrt,
         i_i2c_U_DW_apb_i2c_sync_tx_empty_sync_r,
         i_i2c_U_DW_apb_i2c_sync_ic_rstrt_en_sync_inv,
         i_i2c_U_DW_apb_i2c_sync_ic_10bit_slv_sync_inv,
         i_i2c_U_DW_apb_i2c_sync_tx_empty_int_inv,
         i_i2c_U_DW_apb_i2c_sync_ic_10bit_mst_sync_inv,
         i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv,
         i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv,
         i_i2c_U_DW_apb_i2c_intctl_N4,
         i_i2c_U_DW_apb_i2c_intctl_set_tx_empty_en_flg_sync_q,
         i_i2c_U_DW_apb_i2c_intctl_slv_clr_leftover_flg_sync_q,
         i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync_q,
         i_i2c_U_DW_apb_i2c_intctl_s_det_flg_sync_q,
         i_i2c_U_DW_apb_i2c_intctl_p_det_flg_sync_q,
         i_i2c_U_DW_apb_i2c_intctl_ic_rd_req_flg_sync_q,
         i_i2c_U_DW_apb_i2c_intctl_rx_done_flg_sync_q,
         i_i2c_U_DW_apb_i2c_intctl_tx_abrt_flg_sync_q,
         i_i2c_U_DW_apb_i2c_intctl_set_tx_empty_en_flg_sync,
         i_i2c_U_DW_apb_i2c_intctl_slv_clr_leftover_flg_sync,
         i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync,
         i_i2c_U_DW_apb_i2c_intctl_s_det_flg_sync,
         i_i2c_U_DW_apb_i2c_intctl_p_det_flg_sync,
         i_i2c_U_DW_apb_i2c_intctl_ic_rd_req_flg_sync,
         i_i2c_U_DW_apb_i2c_intctl_rx_done_flg_sync,
         i_i2c_U_DW_apb_i2c_intctl_tx_abrt_flg_sync,
         i_i2c_U_DW_apb_i2c_tx_shift_N402,
         i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly2,
         i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly1,
         i_i2c_U_DW_apb_i2c_tx_shift_N281,
         i_i2c_U_DW_apb_i2c_tx_shift_stop_sda_gate_r,
         i_i2c_U_DW_apb_i2c_tx_shift_N272,
         i_i2c_U_DW_apb_i2c_tx_shift_start_sda_gate_r,
         i_i2c_U_DW_apb_i2c_tx_shift_slv_data_sda,
         i_i2c_U_DW_apb_i2c_tx_shift_data_sda,
         i_i2c_U_DW_apb_i2c_tx_shift_data_sda_prev_r,
         i_i2c_U_DW_apb_i2c_tx_shift_stop_sda,
         i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda,
         i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda_r,
         i_i2c_U_DW_apb_i2c_tx_shift_start_sda,
         i_i2c_U_DW_apb_i2c_tx_shift_byte_wait_en,
         i_i2c_U_DW_apb_i2c_tx_shift_mst_tx_bwen,
         i_i2c_U_DW_apb_i2c_tx_shift_N90,
         i_i2c_U_DW_apb_i2c_tx_shift_data_scl_lcnt_en,
         i_i2c_U_DW_apb_i2c_tx_shift_re_scl_s_hld_en,
         i_i2c_U_DW_apb_i2c_tx_shift_st_scl_s_hld_en,
         i_i2c_U_DW_apb_i2c_tx_shift_N85,
         i_i2c_U_DW_apb_i2c_tx_shift_mst_slv_ack_ext_r,
         i_i2c_U_DW_apb_i2c_tx_shift_mst_slv_ack_ext,
         i_i2c_U_DW_apb_i2c_tx_shift_N74,
         i_i2c_U_DW_apb_i2c_tx_shift_ic_data_oe_early,
         i_i2c_U_DW_apb_i2c_tx_shift_scl_hld_low_en_r,
         i_i2c_U_DW_apb_i2c_tx_shift_stop_scl_lcnt_en,
         i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl_lcnt_en,
         i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl,
         i_i2c_U_DW_apb_i2c_tx_shift_stop_scl,
         i_i2c_U_DW_apb_i2c_tx_shift_data_scl,
         i_i2c_U_DW_apb_i2c_rx_shift_rx_slv_read_s,
         i_i2c_U_DW_apb_i2c_rx_shift_N30,
         i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_3_,
         i_i2c_U_DW_apb_i2c_slvfsm_N284,
         i_i2c_U_DW_apb_i2c_slvfsm_ic_enable_sync_vld,
         i_i2c_U_DW_apb_i2c_slvfsm_slv_tx_flush, i_i2c_U_DW_apb_i2c_slvfsm_N39,
         i_i2c_U_DW_apb_i2c_slvfsm_N38, i_i2c_U_DW_apb_i2c_slvfsm_N37,
         i_i2c_U_DW_apb_i2c_mstfsm_N487,
         i_i2c_U_DW_apb_i2c_mstfsm_mst_gen_ack_en_r,
         i_i2c_U_DW_apb_i2c_mstfsm_N421, i_i2c_U_DW_apb_i2c_mstfsm_N382,
         i_i2c_U_DW_apb_i2c_mstfsm_N252,
         i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_sync_d,
         i_i2c_U_DW_apb_i2c_mstfsm_delay_stop_en,
         i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_chk_win,
         i_i2c_U_DW_apb_i2c_mstfsm_tx_empty_hld,
         i_i2c_U_DW_apb_i2c_mstfsm_abrt_in_idle,
         i_i2c_U_DW_apb_i2c_mstfsm_mst_tx_flush,
         i_i2c_U_DW_apb_i2c_mstfsm_byte_waiting_q,
         i_i2c_U_DW_apb_i2c_mstfsm_old_is_read, i_i2c_U_DW_apb_i2c_mstfsm_N76,
         i_i2c_U_DW_apb_i2c_mstfsm_N75, i_i2c_U_DW_apb_i2c_mstfsm_N74,
         i_i2c_U_DW_apb_i2c_mstfsm_N73, i_i2c_U_DW_apb_i2c_mstfsm_N72,
         i_i2c_U_DW_apb_i2c_mstfsm_addr_1byte_sent,
         i_i2c_U_DW_apb_i2c_mstfsm_addr_2byte_sent,
         i_i2c_U_DW_apb_i2c_rx_filter_N241,
         i_i2c_U_DW_apb_i2c_rx_filter_slv_arb_lost,
         i_i2c_U_DW_apb_i2c_rx_filter_mst_arb_lost,
         i_i2c_U_DW_apb_i2c_rx_filter_N207,
         i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_q,
         i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_qq,
         i_i2c_U_DW_apb_i2c_rx_filter_sda_post_hold_done,
         i_i2c_U_DW_apb_i2c_rx_filter_N130, i_i2c_U_DW_apb_i2c_rx_filter_N129,
         i_i2c_U_DW_apb_i2c_rx_filter_N128, i_i2c_U_DW_apb_i2c_rx_filter_N127,
         i_i2c_U_DW_apb_i2c_rx_filter_N126, i_i2c_U_DW_apb_i2c_rx_filter_N125,
         i_i2c_U_DW_apb_i2c_rx_filter_N124, i_i2c_U_DW_apb_i2c_rx_filter_N123,
         i_i2c_U_DW_apb_i2c_rx_filter_sda_data_int,
         i_i2c_U_DW_apb_i2c_rx_filter_N89, i_i2c_U_DW_apb_i2c_rx_filter_N88,
         i_i2c_U_DW_apb_i2c_rx_filter_N87, i_i2c_U_DW_apb_i2c_rx_filter_N86,
         i_i2c_U_DW_apb_i2c_rx_filter_N85, i_i2c_U_DW_apb_i2c_rx_filter_N84,
         i_i2c_U_DW_apb_i2c_rx_filter_N83,
         i_i2c_U_DW_apb_i2c_rx_filter_scl_clk_int,
         i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r,
         i_i2c_U_DW_apb_i2c_rx_filter_ic_hs, i_i2c_U_DW_apb_i2c_rx_filter_N50,
         i_i2c_U_DW_apb_i2c_rx_filter_hs_mcode_fed_dtctd_r,
         i_i2c_U_DW_apb_i2c_rx_filter_hs_mcode_en_r,
         i_i2c_U_DW_apb_i2c_rx_filter_rx_hs_mcode_r,
         i_i2c_U_DW_apb_i2c_rx_filter_scl_edg_hl_q,
         i_i2c_U_DW_apb_i2c_rx_filter_s_det_int,
         i_i2c_U_DW_apb_i2c_rx_filter_sda_int_q,
         i_i2c_U_DW_apb_i2c_rx_filter_scl_int_q,
         i_i2c_U_DW_apb_i2c_clk_gen_scl_int_d,
         i_i2c_U_DW_apb_i2c_clk_gen_scl_hcnt_cmplt_int,
         i_i2c_U_DW_apb_i2c_clk_gen_N77, i_i2c_U_DW_apb_i2c_clk_gen_N76,
         i_i2c_U_DW_apb_i2c_clk_gen_N75, i_i2c_U_DW_apb_i2c_clk_gen_N74,
         i_i2c_U_DW_apb_i2c_clk_gen_N73, i_i2c_U_DW_apb_i2c_clk_gen_N72,
         i_i2c_U_DW_apb_i2c_clk_gen_N71, i_i2c_U_DW_apb_i2c_clk_gen_N70,
         i_i2c_U_DW_apb_i2c_clk_gen_N69, i_i2c_U_DW_apb_i2c_clk_gen_N68,
         i_i2c_U_DW_apb_i2c_clk_gen_N67, i_i2c_U_DW_apb_i2c_clk_gen_N66,
         i_i2c_U_DW_apb_i2c_clk_gen_N65, i_i2c_U_DW_apb_i2c_clk_gen_N64,
         i_i2c_U_DW_apb_i2c_clk_gen_N63, i_i2c_U_DW_apb_i2c_clk_gen_N62,
         i_i2c_U_DW_apb_i2c_clk_gen_N51, i_i2c_U_DW_apb_i2c_clk_gen_count_en,
         i_i2c_U_DW_apb_i2c_fifo_i_rx_almost_full,
         i_i2c_U_DW_apb_i2c_fifo_rx_error_ir,
         i_i2c_U_DW_apb_i2c_fifo_tx_error_ir,
         i_i2c_U_DW_apb_i2c_fifo_rx_push_sync_dly,
         i_i2c_U_DW_apb_i2c_fifo_rx_pop_dly,
         i_i2c_U_DW_apb_i2c_fifo_tx_pop_sync_dly,
         i_i2c_U_DW_apb_i2c_fifo_tx_push_dly,
         i_i2c_U_DW_apb_i2c_fifo_rx_push_flg_sync_q,
         i_i2c_U_DW_apb_i2c_fifo_tx_pop_flg_sync_q,
         i_i2c_U_DW_apb_i2c_fifo_rx_push_flg_sync,
         i_i2c_U_DW_apb_i2c_fifo_tx_pop_flg_sync, i_ssi_U_regfile_N452,
         i_ssi_U_regfile_N451, i_ssi_U_regfile_multi_mst_edge,
         i_ssi_U_regfile_sr_6_, i_ssi_U_regfile_ctrlr0_ir_int_7,
         i_ssi_U_sclkgen_N75, i_ssi_U_sclkgen_N74, i_ssi_U_sclkgen_N55,
         i_ssi_U_sclkgen_N54, i_ssi_U_sclkgen_N53, i_ssi_U_sclkgen_N52,
         i_ssi_U_sclkgen_N51, i_ssi_U_sclkgen_N50, i_ssi_U_sclkgen_N49,
         i_ssi_U_sclkgen_N48, i_ssi_U_sclkgen_N47, i_ssi_U_sclkgen_N46,
         i_ssi_U_sclkgen_N45, i_ssi_U_sclkgen_N44, i_ssi_U_sclkgen_N43,
         i_ssi_U_sclkgen_N42, i_ssi_U_sclkgen_N41,
         i_ssi_U_fifo_switch_almost_full, i_ssi_U_fifo_rx_push_edge,
         i_ssi_U_fifo_tx_pop_edge, i_ssi_U_fifo_rx_error_ir,
         i_ssi_U_fifo_tx_error_ir, i_ssi_U_fifo_rx_push_sync_dly,
         i_ssi_U_fifo_rx_pop_dly, i_ssi_U_fifo_tx_pop_sync_dly,
         i_ssi_U_fifo_tx_push_dly, i_ssi_U_mstfsm_abort_ir,
         i_ssi_U_mstfsm_N222, i_ssi_U_mstfsm_N221, i_ssi_U_mstfsm_N220,
         i_ssi_U_mstfsm_N219, i_ssi_U_mstfsm_last_frame,
         i_ssi_U_mstfsm_spi1_control, i_ssi_U_mstfsm_spi0_control,
         i_ssi_U_mstfsm_c_done_ir, i_ssi_U_mstfsm_ss_in_n_sync,
         i_ssi_U_mstfsm_tx_load_en_int, i_ssi_U_intctl_N33,
         i_i2c_U_DW_apb_i2c_sync_U_ic_enable_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_abort_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_gen_call_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_master_1_sync_N2,
         i_i2c_U_DW_apb_i2c_sync_U_ic_master_1_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_hs_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_fs_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_ss_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_mst_1_sync_N2,
         i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_mst_1_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_tx_empty_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_slv_1_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_rstrt_en_1_sync_N2,
         i_i2c_U_DW_apb_i2c_sync_U_ic_rstrt_en_1_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_ic_slave_en_1_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_sync_U_p_det_ifaddr_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_rx_done_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_ic_rd_req_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_p_det_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_s_det_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_rx_gen_call_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_slv_clr_leftover_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_set_tx_empty_en_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_mst_activity_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_slv_activity_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_slv_rx_aborted_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_intctl_U_slv_fifo_filled_and_flushed_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_data_d_int_0_,
         i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_data_d_int_0_,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_pop_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_push_flg_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N48,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N46,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N45,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N44,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N43,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N42,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N41,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N40,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N39,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N38,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N37,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N34,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N33,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_almost_empty_n,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_rd_addr_at_max,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_wr_addr_at_max,
         i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_empty_n,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N49,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N48,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N47,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N46,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N45,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N44,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N43,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N42,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N41,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N40,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N39,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N38,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N37,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N36,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N33,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_rd_addr_at_max,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_wr_addr_at_max,
         i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_empty_n, i_ssi_U_fifo_U_tx_fifo_N46,
         i_ssi_U_fifo_U_tx_fifo_N45, i_ssi_U_fifo_U_tx_fifo_N43,
         i_ssi_U_fifo_U_tx_fifo_N42, i_ssi_U_fifo_U_tx_fifo_N40,
         i_ssi_U_fifo_U_tx_fifo_N39, i_ssi_U_fifo_U_tx_fifo_N38,
         i_ssi_U_fifo_U_tx_fifo_N34, i_ssi_U_fifo_U_tx_fifo_N33,
         i_ssi_U_fifo_U_tx_fifo_almost_empty_n,
         i_ssi_U_fifo_U_tx_fifo_rd_addr_at_max,
         i_ssi_U_fifo_U_tx_fifo_wr_addr_at_max, i_ssi_U_fifo_U_tx_fifo_empty_n,
         i_ssi_U_fifo_U_rx_fifo_N46, i_ssi_U_fifo_U_rx_fifo_N45,
         i_ssi_U_fifo_U_rx_fifo_N43, i_ssi_U_fifo_U_rx_fifo_N42,
         i_ssi_U_fifo_U_rx_fifo_N40, i_ssi_U_fifo_U_rx_fifo_N39,
         i_ssi_U_fifo_U_rx_fifo_N38, i_ssi_U_fifo_U_rx_fifo_N33,
         i_ssi_U_fifo_U_rx_fifo_rd_addr_at_max,
         i_ssi_U_fifo_U_rx_fifo_wr_addr_at_max, i_ssi_U_fifo_U_rx_fifo_empty_n,
         i_ssi_U_shift_U_tx_shifter_load_start_bit_ir,
         i_ssi_U_mstfsm_U_ss_in_n_sync_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_U_SYNC_N2,
         i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_U_SYNC_next_sample_syncm1_0_,
         i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_U_SYNC_N2,
         i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_U_SYNC_next_sample_syncm1_0_,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4187,
         n4189, n4190, n4191, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4817,
         n4818, n4819, n4835, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5103, n5104, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5234, n5235, n5240, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11794, n11795, n11816, n11829, n11830,
         n11831, ex_i_ahb_AHB_Slave_PID_hready, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         ex_i_ahb_AHB_MASTER_CORTEXM0_hready, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14;
  wire   [31:12] i_apb_paddr;
  wire   [31:0] i_ssi_prdata;
  wire   [30:0] i_i2c_prdata;
  wire   [23:0] i_apb_pwdata_int;
  wire   [2:0] i_i2c_rx_rd_addr;
  wire   [2:0] i_i2c_rx_wr_addr;
  wire   [2:0] i_i2c_tx_rd_addr;
  wire   [2:0] i_i2c_tx_wr_addr;
  wire   [7:0] i_i2c_rx_pop_data;
  wire   [2:0] i_i2c_ic_tx_tl;
  wire   [2:0] i_i2c_ic_rx_tl;
  wire   [15:0] i_i2c_ic_fs_hcnt;
  wire   [15:0] i_i2c_ic_fs_lcnt;
  wire   [15:0] i_i2c_ic_lcnt;
  wire   [15:0] i_i2c_ic_hcnt;
  wire   [7:0] i_i2c_ic_fs_spklen;
  wire   [7:0] i_i2c_ic_hs_spklen;
  wire   [10:0] i_i2c_ic_tar;
  wire   [2:0] i_i2c_ic_hs_maddr;
  wire   [7:0] i_i2c_ic_sda_setup;
  wire   [30:0] i_i2c_iprdata;
  wire   [7:0] i_i2c_rx_push_data;
  wire   [9:0] i_i2c_ic_sar;
  wire   [3:0] i_i2c_mst_rx_bit_count;
  wire   [8:0] i_i2c_tx_fifo_data_buf;
  wire   [16:0] i_i2c_ic_tx_abrt_source;
  wire   [11:0] i_i2c_ic_raw_intr_stat;
  wire   [11:0] i_i2c_ic_intr_stat;
  wire   [11:0] i_i2c_ic_intr_mask;
  wire   [7:0] i_i2c_ic_sda_rx_hold_sync;
  wire   [15:0] i_i2c_ic_sda_tx_hold_sync;
  wire   [23:0] i_i2c_ic_sda_hold;
  wire   [1:0] i_i2c_ic_enable;
  wire   [16:0] i_i2c_tx_abrt_source;
  wire   [3:0] i_i2c_slv_debug_cstate;
  wire   [4:0] i_i2c_mst_debug_cstate;
  wire   [15:0] i_ssi_rx_push_data;
  wire   [2:0] i_ssi_rx_rd_addr;
  wire   [2:0] i_ssi_rx_wr_addr;
  wire   [2:0] i_ssi_tx_rd_addr;
  wire   [2:0] i_ssi_tx_wr_addr;
  wire   [2:0] i_ssi_rxftlr;
  wire   [2:0] i_ssi_txftlr;
  wire   [15:1] i_ssi_baudr;
  wire   [2:0] i_ssi_mwcr;
  wire   [5:0] i_ssi_imr;
  wire   [5:0] i_ssi_risr;
  wire   [5:0] i_ssi_reg_addr;
  wire   [3:0] i_ssi_cfs;
  wire   [1:0] i_ssi_tmod;
  wire   [11:10] i_ssi_ctrlr0;
  wire   [3:0] i_ssi_dfs;
  wire   [4:1] i_ahb_U_mux_hsel_prev;
  wire   [23:0] i_apb_U_DW_apb_ahbsif_saved_hwdata32_c;
  wire   [31:2] i_apb_U_DW_apb_ahbsif_saved_haddr_c;
  wire   [16:2] i_apb_U_DW_apb_ahbsif_piped_haddr_c;
  wire   [2:0] i_apb_U_DW_apb_ahbsif_nextstate;
  wire   [2:0] i_apb_U_DW_apb_ahbsif_state;
  wire   [16:0] i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q;
  wire   [16:0] i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync;
  wire   [15:0] i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r;
  wire   [7:0] i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf;
  wire   [3:0] i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count;
  wire   [3:0] i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count;
  wire   [3:0] i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr;
  wire   [7:0] i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg;
  wire   [7:0] i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg;
  wire   [2:0] i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0;
  wire   [7:0] i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count;
  wire  
         [3:0] i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en
;
  wire   [1:0] i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt;
  wire   [7:0] i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt;
  wire   [7:0] i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt;
  wire   [7:0] i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt;
  wire   [15:0] i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr;
  wire   [15:0] i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr;
  wire   [15:0] i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr;
  wire   [15:0] i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr;
  wire   [15:0] i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr;
  wire   [15:0] i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr;
  wire   [15:0] i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr;
  wire   [2:0] i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn;
  wire   [2:0] i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn;
  wire   [7:0] i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr;
  wire   [63:0] i_i2c_U_dff_rx_mem;
  wire   [71:0] i_i2c_U_dff_tx_mem;
  wire   [3:0] i_ssi_U_regfile_rxflr;
  wire   [3:0] i_ssi_U_regfile_txflr;
  wire   [15:0] i_ssi_U_regfile_ctrlr1_int;
  wire   [5:4] i_ssi_U_regfile_ctrlr0_ir_int;
  wire   [15:0] i_ssi_U_sclkgen_ssi_cnt;
  wire   [2:0] i_ssi_U_fifo_unconnected_rx_wrd_count;
  wire   [2:0] i_ssi_U_fifo_unconnected_tx_wrd_count;
  wire   [16:0] i_ssi_U_mstfsm_frame_cnt;
  wire   [3:0] i_ssi_U_mstfsm_c_state;
  wire   [3:0] i_ssi_U_mstfsm_ctrl_cnt;
  wire   [4:0] i_ssi_U_mstfsm_bit_cnt;
  wire   [127:0] i_ssi_U_dff_rx_mem;
  wire   [127:0] i_ssi_U_dff_tx_mem;
  wire   [23:0] i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1;
  wire  
         [16:0] i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1
;
  wire   [15:0] i_ssi_U_shift_U_tx_shifter_tx_buffer;
  wire   [15:0] i_ssi_U_shift_U_tx_shifter_tx_shift_reg;
  wire   [15:0] i_ssi_U_shift_U_rx_shifter_rx_shift_reg;
  assign ex_i_ahb_AHB_Slave_RAM_haddr[31] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[31];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[31] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[31];
  assign ex_i_ahb_AHB_Slave_PID_haddr[31] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[31];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[30] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[30];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[30] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[30];
  assign ex_i_ahb_AHB_Slave_PID_haddr[30] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[30];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[29] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[29];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[29] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[29];
  assign ex_i_ahb_AHB_Slave_PID_haddr[29] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[29];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[28] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[28];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[28] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[28];
  assign ex_i_ahb_AHB_Slave_PID_haddr[28] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[28];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[27] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[27];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[27] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[27];
  assign ex_i_ahb_AHB_Slave_PID_haddr[27] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[27];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[26] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[26];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[26] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[26];
  assign ex_i_ahb_AHB_Slave_PID_haddr[26] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[26];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[25] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[25];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[25] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[25];
  assign ex_i_ahb_AHB_Slave_PID_haddr[25] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[25];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[24] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[24];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[24] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[24];
  assign ex_i_ahb_AHB_Slave_PID_haddr[24] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[24];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[23] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[23];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[23] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[23];
  assign ex_i_ahb_AHB_Slave_PID_haddr[23] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[23];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[22] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[22];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[22] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[22];
  assign ex_i_ahb_AHB_Slave_PID_haddr[22] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[22];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[21] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[21];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[21] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[21];
  assign ex_i_ahb_AHB_Slave_PID_haddr[21] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[21];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[20] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[20];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[20] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[20];
  assign ex_i_ahb_AHB_Slave_PID_haddr[20] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[20];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[19] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[19];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[19] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[19];
  assign ex_i_ahb_AHB_Slave_PID_haddr[19] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[19];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[18] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[18];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[18] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[18];
  assign ex_i_ahb_AHB_Slave_PID_haddr[18] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[18];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[17] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[17];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[17] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[17];
  assign ex_i_ahb_AHB_Slave_PID_haddr[17] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[17];
  assign ex_i_ahb_AHB_Slave_PID_haddr[16] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[16];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[16] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[16];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[16] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[16];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[15] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[15];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[15] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[15];
  assign ex_i_ahb_AHB_Slave_PID_haddr[15] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[15];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[14] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[14];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[14] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[14];
  assign ex_i_ahb_AHB_Slave_PID_haddr[14] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[14];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[13] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[13];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[13] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[13];
  assign ex_i_ahb_AHB_Slave_PID_haddr[13] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[13];
  assign ex_i_ahb_AHB_Slave_PID_haddr[12] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[12];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[12] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[12];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[12] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[12];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[11] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[11];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[11] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[11];
  assign ex_i_ahb_AHB_Slave_PID_haddr[11] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[11];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[10] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[10];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[10] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[10];
  assign ex_i_ahb_AHB_Slave_PID_haddr[10] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[10];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[9] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[9];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[9] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[9];
  assign ex_i_ahb_AHB_Slave_PID_haddr[9] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[9];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[8] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[8];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[8] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[8];
  assign ex_i_ahb_AHB_Slave_PID_haddr[8] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[8];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[7] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[7];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[7] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[7];
  assign ex_i_ahb_AHB_Slave_PID_haddr[7] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[7];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[6] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[6];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[6] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[6];
  assign ex_i_ahb_AHB_Slave_PID_haddr[6] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[6];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[5] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[5];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[5] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[5];
  assign ex_i_ahb_AHB_Slave_PID_haddr[5] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[5];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[4] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[4];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[4] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[4];
  assign ex_i_ahb_AHB_Slave_PID_haddr[4] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[4];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[3] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[3];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[3] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[3];
  assign ex_i_ahb_AHB_Slave_PID_haddr[3] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[3];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[2];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[2];
  assign ex_i_ahb_AHB_Slave_PID_haddr[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[2];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[1];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[1];
  assign ex_i_ahb_AHB_Slave_PID_haddr[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[1];
  assign ex_i_ahb_AHB_Slave_RAM_haddr[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[0];
  assign ex_i_ahb_AHB_Slave_PWM_haddr[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[0];
  assign ex_i_ahb_AHB_Slave_PID_haddr[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[0];
  assign ex_i_ahb_AHB_Slave_RAM_hburst[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hburst[2];
  assign ex_i_ahb_AHB_Slave_PWM_hburst[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hburst[2];
  assign ex_i_ahb_AHB_Slave_PID_hburst[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hburst[2];
  assign ex_i_ahb_AHB_Slave_RAM_hburst[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hburst[1];
  assign ex_i_ahb_AHB_Slave_PWM_hburst[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hburst[1];
  assign ex_i_ahb_AHB_Slave_PID_hburst[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hburst[1];
  assign ex_i_ahb_AHB_Slave_RAM_hburst[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hburst[0];
  assign ex_i_ahb_AHB_Slave_PWM_hburst[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hburst[0];
  assign ex_i_ahb_AHB_Slave_PID_hburst[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hburst[0];
  assign ex_i_ahb_AHB_Slave_RAM_hprot[3] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[3];
  assign ex_i_ahb_AHB_Slave_PWM_hprot[3] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[3];
  assign ex_i_ahb_AHB_Slave_PID_hprot[3] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[3];
  assign ex_i_ahb_AHB_Slave_RAM_hprot[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[2];
  assign ex_i_ahb_AHB_Slave_PWM_hprot[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[2];
  assign ex_i_ahb_AHB_Slave_PID_hprot[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[2];
  assign ex_i_ahb_AHB_Slave_RAM_hprot[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[1];
  assign ex_i_ahb_AHB_Slave_PWM_hprot[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[1];
  assign ex_i_ahb_AHB_Slave_PID_hprot[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[1];
  assign ex_i_ahb_AHB_Slave_RAM_hprot[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[0];
  assign ex_i_ahb_AHB_Slave_PWM_hprot[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[0];
  assign ex_i_ahb_AHB_Slave_PID_hprot[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hprot[0];
  assign ex_i_ahb_AHB_Slave_RAM_hsize[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hsize[2];
  assign ex_i_ahb_AHB_Slave_PWM_hsize[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hsize[2];
  assign ex_i_ahb_AHB_Slave_PID_hsize[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hsize[2];
  assign ex_i_ahb_AHB_Slave_RAM_hsize[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hsize[1];
  assign ex_i_ahb_AHB_Slave_PWM_hsize[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hsize[1];
  assign ex_i_ahb_AHB_Slave_PID_hsize[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hsize[1];
  assign ex_i_ahb_AHB_Slave_RAM_hsize[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hsize[0];
  assign ex_i_ahb_AHB_Slave_PWM_hsize[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hsize[0];
  assign ex_i_ahb_AHB_Slave_PID_hsize[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hsize[0];
  assign ex_i_ahb_AHB_Slave_RAM_htrans[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_htrans[1];
  assign ex_i_ahb_AHB_Slave_PWM_htrans[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_htrans[1];
  assign ex_i_ahb_AHB_Slave_PID_htrans[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_htrans[1];
  assign ex_i_ahb_AHB_Slave_RAM_htrans[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_htrans[0];
  assign ex_i_ahb_AHB_Slave_PWM_htrans[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_htrans[0];
  assign ex_i_ahb_AHB_Slave_PID_htrans[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_htrans[0];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[31] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[31];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[31] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[31];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[31] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[31];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[30] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[30];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[30] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[30];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[30] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[30];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[29] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[29];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[29] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[29];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[29] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[29];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[28] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[28];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[28] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[28];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[28] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[28];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[27] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[27];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[27] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[27];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[27] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[27];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[26] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[26];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[26] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[26];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[26] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[26];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[25] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[25];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[25] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[25];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[25] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[25];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[24] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[24];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[24] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[24];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[24] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[24];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[23] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[23];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[23] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[23];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[23] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[23];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[22] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[22];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[22] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[22];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[22] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[22];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[21] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[21];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[21] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[21];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[21] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[21];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[20] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[20];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[20] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[20];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[20] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[20];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[19] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[19];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[19] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[19];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[19] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[19];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[18] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[18];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[18] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[18];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[18] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[18];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[17] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[17];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[17] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[17];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[17] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[17];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[16] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[16];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[16] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[16];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[16] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[16];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[15] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[15];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[15] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[15];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[15] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[15];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[14] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[14];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[14] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[14];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[14] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[14];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[13] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[13];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[13] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[13];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[13] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[13];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[12] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[12];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[12] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[12];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[12] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[12];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[11] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[11];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[11] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[11];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[11] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[11];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[10] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[10];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[10] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[10];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[10] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[10];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[9] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[9];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[9] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[9];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[9] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[9];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[8] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[8];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[8] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[8];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[8] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[8];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[7] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[7];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[7] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[7];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[7] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[7];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[6] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[6];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[6] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[6];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[6] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[6];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[5] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[5];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[5] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[5];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[5] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[5];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[4] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[4];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[4] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[4];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[4] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[4];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[3] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[3];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[3] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[3];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[3] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[3];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[2];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[2];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[2] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[2];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[1];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[1];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[1] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[1];
  assign ex_i_ahb_AHB_Slave_RAM_hwdata[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[0];
  assign ex_i_ahb_AHB_Slave_PWM_hwdata[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[0];
  assign ex_i_ahb_AHB_Slave_PID_hwdata[0] = ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[0];
  assign ex_i_ahb_AHB_Slave_RAM_hwrite = ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite;
  assign ex_i_ahb_AHB_Slave_PWM_hwrite = ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite;
  assign ex_i_ahb_AHB_Slave_PID_hwrite = ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite;
  assign ex_i_ahb_AHB_Slave_RAM_hmastlock = ex_i_ahb_AHB_Slave_PID_hmastlock;
  assign ex_i_ahb_AHB_Slave_PWM_hmastlock = ex_i_ahb_AHB_Slave_PID_hmastlock;
  assign i_ahb_hmaster_data[0] = 1'b1;
  assign i_ahb_hmaster_data[3] = 1'b0;
  assign i_ahb_hmaster_data[2] = 1'b0;
  assign i_ahb_hmaster_data[1] = 1'b0;
  assign ex_i_ahb_AHB_Slave_PWM_hready = ex_i_ahb_AHB_Slave_PID_hready;
  assign ex_i_ahb_AHB_Slave_RAM_hready = ex_i_ahb_AHB_MASTER_CORTEXM0_hready;

  i_i2c_DW_apb_i2c_regfile i_i2c_U_DW_apb_i2c_regfile ( .pclk(PCLK_pclk), 
        .presetn(PRESETn_presetn), .wr_en(i_i2c_wr_en), .rd_en(n11839), 
        .byte_en({1'b1, 1'b1, 1'b1, 1'b1}), .reg_addr(i_ssi_reg_addr), 
        .ipwdata({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        i_apb_pwdata_int}), .iprdata({SYNOPSYS_UNCONNECTED_1, 
        i_i2c_iprdata[30:29], SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        i_i2c_iprdata[26:0]}), .ic_clr_intr_en(i_i2c_ic_clr_intr_en), 
        .ic_clr_rx_under_en(i_i2c_ic_clr_rx_under_en), .ic_clr_rx_over_en(
        i_i2c_ic_clr_rx_over_en), .ic_clr_tx_over_en(i_i2c_ic_clr_tx_over_en), 
        .ic_clr_rd_req_en(i_i2c_ic_clr_rd_req_en), .ic_clr_tx_abrt_en(
        i_i2c_ic_clr_tx_abrt_en), .ic_clr_rx_done_en(i_i2c_ic_clr_rx_done_en), 
        .ic_clr_activity_en(i_i2c_ic_clr_activity_en), .ic_clr_stop_det_en(
        i_i2c_ic_clr_stop_det_en), .ic_clr_start_det_en(
        i_i2c_ic_clr_start_det_en), .ic_clr_gen_call_en(
        i_i2c_ic_clr_gen_call_en), .mst_activity(i_i2c_mst_activity_sync), 
        .slv_activity(i_i2c_slv_activity_sync), .activity(i_i2c_activity), 
        .ic_tx_abrt_source(i_i2c_ic_tx_abrt_source), .ic_en(i_i2c_ic_en), 
        .slv_rx_aborted_sync(i_i2c_slv_rx_aborted_sync), 
        .slv_fifo_filled_and_flushed_sync(
        i_i2c_slv_fifo_filled_and_flushed_sync), .ic_tar({
        i_i2c_U_DW_apb_i2c_mstfsm_N252, i_i2c_ic_tar}), .ic_sar(i_i2c_ic_sar), 
        .ic_hs_maddr(i_i2c_ic_hs_maddr), .ic_fs_hcnt(i_i2c_ic_fs_hcnt), 
        .ic_fs_lcnt(i_i2c_ic_fs_lcnt), .ic_intr_mask({SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, i_i2c_ic_intr_mask}), .ic_rx_tl_int(
        i_i2c_ic_rx_tl), .ic_enable(i_i2c_ic_enable), .ic_hcnt(i_i2c_ic_hcnt), 
        .ic_lcnt(i_i2c_ic_lcnt), .ic_fs_spklen(i_i2c_ic_fs_spklen), 
        .ic_hs_spklen(i_i2c_ic_hs_spklen), .ic_intr_stat({1'b0, 1'b0, 
        i_i2c_ic_intr_stat}), .ic_raw_intr_stat({1'b0, 1'b0, 
        i_i2c_ic_raw_intr_stat}), .ic_hs(i_i2c_ic_hs), .ic_fs(i_i2c_ic_fs), 
        .ic_ss(i_i2c_ic_ss), .ic_master(i_i2c_ic_master), .ic_10bit_mst(
        i_i2c_ic_10bit_mst), .ic_10bit_slv(i_i2c_ic_10bit_slv), .ic_slave_en(
        i_i2c_ic_slave_en), .p_det_ifaddr(i_i2c_p_det_ifaddr), .tx_empty_ctrl(
        i_i2c_tx_empty_ctrl), .rx_pop_data(i_i2c_rx_pop_data), .tx_push_data({
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14}), .fifo_rst_n(
        i_i2c_fifo_rst_n), .tx_fifo_rst_n(i_i2c_tx_fifo_rst_n), .tx_pop_sync(
        i_i2c_tx_pop_sync), .rx_push_sync(i_i2c_rx_push_sync), .rx_pop(
        i_i2c_rx_pop), .tx_push(i_i2c_tx_push), .tx_empty(n11862), .rx_full(
        i_i2c_rx_full), .tx_full(i_i2c_tx_full), .rx_empty(n5240), 
        .tx_abrt_flg_edg(i_i2c_tx_abrt_flg_edg), .abrt_in_rcve_trns(
        i_i2c_abrt_in_rcve_trns), .slv_clr_leftover_flg_edg(n7398), 
        .ic_rstrt_en(i_i2c_ic_rstrt_en), .ic_sda_setup(i_i2c_ic_sda_setup), 
        .ic_sda_hold(i_i2c_ic_sda_hold), .ic_ack_general_call(
        i_i2c_ic_ack_general_call), .ic_tx_tl_2_(i_i2c_ic_tx_tl[2]), 
        .ic_tx_tl_1_(i_i2c_ic_tx_tl[1]), .ic_tx_tl_0_(i_i2c_ic_tx_tl[0]) );
  drsp_1 i_ssi_U_mstfsm_tx_load_en_reg ( .ip(n4579), .ck(i_ssi_ssi_clk), .rb(
        1'b1), .s(n11841), .q(i_ssi_U_mstfsm_tx_load_en_int) );
  drsp_1 i_i2c_U_DW_apb_i2c_rx_filter_scl_clk_int_reg ( .ip(n5130), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11842), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_scl_clk_int) );
  drp_1 i_ahb_U_dfltslv_current_state_reg ( .ip(i_ahb_U_dfltslv_next_state), 
        .ck(HCLK_hclk), .rb(HRESETn_hresetn), .q(i_ahb_U_dfltslv_current_state) );
  drp_1 i_ahb_U_dfltslv_hresp_none_reg_0_ ( .ip(i_ahb_U_dfltslv_N4), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(i_ahb_hresp_none_0_) );
  drp_1 i_ahb_U_mux_hsel_prev_reg_3_ ( .ip(n4851), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ahb_U_mux_hsel_prev[3]) );
  drp_1 i_ahb_U_mux_hsel_prev_reg_2_ ( .ip(n4850), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ahb_U_mux_hsel_prev[2]) );
  drp_1 i_ahb_U_mux_hsel_prev_reg_1_ ( .ip(n4849), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ahb_U_mux_hsel_prev[1]) );
  drp_1 i_ahb_U_arblite_hmastlock_reg ( .ip(n4848), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(ex_i_ahb_AHB_Slave_PID_hmastlock) );
  drp_1 i_apb_U_DW_apb_ahbsif_state_reg_0_ ( .ip(
        i_apb_U_DW_apb_ahbsif_nextstate[0]), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_state[0]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pipeline_reg ( .ip(n4847), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_pipeline_c) );
  drp_1 i_apb_U_DW_apb_ahbsif_state_reg_1_ ( .ip(
        i_apb_U_DW_apb_ahbsif_nextstate[1]), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_state[1]) );
  drp_1 i_apb_U_DW_apb_ahbsif_state_reg_2_ ( .ip(
        i_apb_U_DW_apb_ahbsif_nextstate[2]), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_state[2]) );
  drp_1 i_apb_U_DW_apb_ahbsif_piped_hwrite_reg ( .ip(n4846), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_piped_hwrite_c) );
  drp_1 i_apb_U_DW_apb_ahbsif_piped_haddr_reg_2_ ( .ip(n4845), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_piped_haddr_c[2]) );
  drp_1 i_apb_U_DW_apb_ahbsif_piped_haddr_reg_3_ ( .ip(n4844), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_piped_haddr_c[3]) );
  drp_1 i_apb_U_DW_apb_ahbsif_piped_haddr_reg_4_ ( .ip(n4843), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_piped_haddr_c[4]) );
  drp_1 i_apb_U_DW_apb_ahbsif_piped_haddr_reg_5_ ( .ip(n4842), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_piped_haddr_c[5]) );
  drp_1 i_apb_U_DW_apb_ahbsif_piped_haddr_reg_6_ ( .ip(n4841), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_piped_haddr_c[6]) );
  drp_1 i_apb_U_DW_apb_ahbsif_piped_haddr_reg_7_ ( .ip(n4840), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_piped_haddr_c[7]) );
  drp_1 i_apb_U_DW_apb_ahbsif_piped_haddr_reg_12_ ( .ip(n4839), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_piped_haddr_c[12]) );
  drp_1 i_apb_U_DW_apb_ahbsif_piped_haddr_reg_16_ ( .ip(n4835), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_piped_haddr_c[16]) );
  drp_1 i_apb_U_DW_apb_ahbsif_use_saved_reg ( .ip(n4819), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_use_saved_c) );
  drp_1 i_apb_U_DW_apb_ahbsif_use_saved_data_reg ( .ip(
        i_apb_U_DW_apb_ahbsif_N727), .ck(HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_use_saved_data) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_0_ ( .ip(n4815), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[0]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_1_ ( .ip(n4814), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[1]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_2_ ( .ip(n4813), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[2]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_3_ ( .ip(n4812), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[3]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_4_ ( .ip(n4811), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[4]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_5_ ( .ip(n4810), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[5]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_6_ ( .ip(n4809), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[6]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_7_ ( .ip(n4808), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[7]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_8_ ( .ip(n4807), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[8]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_9_ ( .ip(n4806), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[9]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_10_ ( .ip(n4805), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[10]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_11_ ( .ip(n4804), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[11]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_12_ ( .ip(n4803), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[12]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_13_ ( .ip(n4802), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[13]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_14_ ( .ip(n4801), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[14]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_15_ ( .ip(n4800), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[15]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_16_ ( .ip(n4799), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[16]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_17_ ( .ip(n4798), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[17]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_18_ ( .ip(n4797), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[18]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_19_ ( .ip(n4796), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[19]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_20_ ( .ip(n4795), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[20]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_21_ ( .ip(n4794), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[21]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_22_ ( .ip(n4793), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[22]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_hwdata32_reg_23_ ( .ip(n4792), .ck(
        HCLK_hclk), .rb(HRESETn_hresetn), .q(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[23]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_2_ ( .ip(n4752), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[2]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_3_ ( .ip(n4751), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[3]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_4_ ( .ip(n4750), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[4]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_5_ ( .ip(n4749), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[5]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_6_ ( .ip(n4748), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[6]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_7_ ( .ip(n4747), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[7]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_12_ ( .ip(n4746), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[12]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_13_ ( .ip(n4745), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[13]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_14_ ( .ip(n4744), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[14]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_15_ ( .ip(n4743), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[15]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_16_ ( .ip(n4742), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[16]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_17_ ( .ip(n4741), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[17]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_18_ ( .ip(n4740), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[18]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_19_ ( .ip(n4739), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[19]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_20_ ( .ip(n4738), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[20]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_21_ ( .ip(n4737), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[21]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_22_ ( .ip(n4736), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[22]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_23_ ( .ip(n4735), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[23]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_24_ ( .ip(n4734), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[24]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_25_ ( .ip(n4733), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[25]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_26_ ( .ip(n4732), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[26]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_27_ ( .ip(n4731), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[27]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_28_ ( .ip(n4730), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[28]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_29_ ( .ip(n4729), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[29]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_30_ ( .ip(n4728), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[30]) );
  drp_1 i_apb_U_DW_apb_ahbsif_saved_haddr_reg_31_ ( .ip(n4727), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_U_DW_apb_ahbsif_saved_haddr_c[31]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_0_ ( .ip(n4784), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[0]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_1_ ( .ip(n4783), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[1]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_2_ ( .ip(n4782), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[2]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_3_ ( .ip(n4781), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[3]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_4_ ( .ip(n4780), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[4]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_5_ ( .ip(n4779), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[5]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_6_ ( .ip(n4778), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[6]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_7_ ( .ip(n4777), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[7]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_8_ ( .ip(n4776), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[8]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_9_ ( .ip(n4775), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[9]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_10_ ( .ip(n4774), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[10]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_11_ ( .ip(n4773), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[11]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_12_ ( .ip(n4772), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[12]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_13_ ( .ip(n4771), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[13]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_14_ ( .ip(n4770), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[14]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_15_ ( .ip(n4769), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[15]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_16_ ( .ip(n4768), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[16]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_17_ ( .ip(n4767), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[17]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_18_ ( .ip(n4766), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[18]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_19_ ( .ip(n4765), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[19]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_20_ ( .ip(n4764), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[20]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_21_ ( .ip(n4763), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[21]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_22_ ( .ip(n4762), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[22]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwdata_int_reg_23_ ( .ip(n4761), .ck(HCLK_hclk), 
        .rb(HRESETn_hresetn), .q(i_apb_pwdata_int[23]) );
  drp_1 i_apb_U_DW_apb_ahbsif_pwrite_reg ( .ip(n4818), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_pwrite) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_2_ ( .ip(n4726), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ssi_reg_addr[0]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_3_ ( .ip(n4725), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ssi_reg_addr[1]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_4_ ( .ip(n4724), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ssi_reg_addr[2]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_5_ ( .ip(n4723), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ssi_reg_addr[3]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_6_ ( .ip(n4722), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ssi_reg_addr[4]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_7_ ( .ip(n4721), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ssi_reg_addr[5]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_12_ ( .ip(n4720), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[12]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_13_ ( .ip(n4719), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[13]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_14_ ( .ip(n4718), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[14]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_15_ ( .ip(n4717), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[15]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_16_ ( .ip(n4716), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[16]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_17_ ( .ip(n4715), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[17]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_18_ ( .ip(n4714), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[18]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_19_ ( .ip(n4713), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[19]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_20_ ( .ip(n4712), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[20]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_21_ ( .ip(n4711), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[21]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_22_ ( .ip(n4710), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[22]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_23_ ( .ip(n4709), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[23]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_24_ ( .ip(n4708), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[24]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_25_ ( .ip(n4707), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[25]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_26_ ( .ip(n4706), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[26]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_27_ ( .ip(n4705), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[27]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_28_ ( .ip(n4704), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[28]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_29_ ( .ip(n4703), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[29]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_30_ ( .ip(n4702), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[30]) );
  drp_1 i_apb_U_DW_apb_ahbsif_paddr_reg_31_ ( .ip(n4701), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_paddr[31]) );
  drp_1 i_ssi_U_biu_prdata_reg_16_ ( .ip(n4221), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[16]) );
  drp_1 i_ssi_U_biu_prdata_reg_17_ ( .ip(n4220), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[17]) );
  drp_1 i_ssi_U_biu_prdata_reg_18_ ( .ip(n4219), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[18]) );
  drp_1 i_ssi_U_biu_prdata_reg_19_ ( .ip(n4218), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[19]) );
  drp_1 i_ssi_U_biu_prdata_reg_20_ ( .ip(n4217), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[20]) );
  drp_1 i_ssi_U_biu_prdata_reg_21_ ( .ip(n4216), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[21]) );
  drp_1 i_ssi_U_biu_prdata_reg_22_ ( .ip(n4215), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[22]) );
  drp_1 i_ssi_U_biu_prdata_reg_23_ ( .ip(n4214), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[23]) );
  drp_1 i_ssi_U_biu_prdata_reg_24_ ( .ip(n4213), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[24]) );
  drp_1 i_ssi_U_biu_prdata_reg_25_ ( .ip(n4212), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[25]) );
  drp_1 i_ssi_U_biu_prdata_reg_26_ ( .ip(n4211), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[26]) );
  drp_1 i_ssi_U_biu_prdata_reg_27_ ( .ip(n4210), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[27]) );
  drp_1 i_ssi_U_biu_prdata_reg_28_ ( .ip(n4209), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[28]) );
  drp_1 i_ssi_U_biu_prdata_reg_29_ ( .ip(n4208), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[29]) );
  drp_1 i_ssi_U_biu_prdata_reg_30_ ( .ip(n4207), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[30]) );
  drp_1 i_ssi_U_biu_prdata_reg_31_ ( .ip(n4206), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[31]) );
  drp_1 i_ssi_U_regfile_ser_reg_0_ ( .ip(n4627), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_ser_0_) );
  drp_1 i_ssi_U_regfile_rxftlr_reg_0_ ( .ip(n4637), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_rxftlr[0]) );
  drp_1 i_ssi_U_regfile_rxftlr_reg_1_ ( .ip(n4636), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_rxftlr[1]) );
  drp_1 i_ssi_U_regfile_rxftlr_reg_2_ ( .ip(n4635), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_rxftlr[2]) );
  drp_1 i_ssi_U_regfile_txftlr_reg_0_ ( .ip(n4634), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_txftlr[0]) );
  drp_1 i_ssi_U_regfile_txftlr_reg_1_ ( .ip(n4633), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_txftlr[1]) );
  drp_1 i_ssi_U_regfile_txftlr_reg_2_ ( .ip(n4632), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_txftlr[2]) );
  drp_1 i_ssi_U_regfile_ssienr_reg ( .ip(n4631), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_ssi_en_int) );
  drp_1 i_ssi_U_regfile_mwcr_ir_reg_0_ ( .ip(n4630), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_mwcr[0]) );
  drp_1 i_ssi_U_regfile_mwcr_ir_reg_1_ ( .ip(n4629), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_mwcr[1]) );
  drp_1 i_ssi_U_regfile_mwcr_ir_reg_2_ ( .ip(n4628), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_mwcr[2]) );
  drp_1 i_ssi_U_regfile_baudr_reg_4_ ( .ip(n4623), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[4]) );
  drp_1 i_ssi_U_regfile_baudr_reg_8_ ( .ip(n4619), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[8]) );
  drp_1 i_ssi_U_regfile_baudr_reg_9_ ( .ip(n4618), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[9]) );
  drp_1 i_ssi_U_regfile_baudr_reg_10_ ( .ip(n4617), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[10]) );
  drp_1 i_ssi_U_regfile_baudr_reg_11_ ( .ip(n4616), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[11]) );
  drp_1 i_ssi_U_regfile_baudr_reg_12_ ( .ip(n4615), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[12]) );
  drp_1 i_ssi_U_regfile_baudr_reg_13_ ( .ip(n4614), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[13]) );
  drp_1 i_ssi_U_regfile_baudr_reg_14_ ( .ip(n4613), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[14]) );
  drp_1 i_ssi_U_regfile_baudr_reg_15_ ( .ip(n4612), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[15]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_0_ ( .ip(n4603), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[0]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_1_ ( .ip(n4602), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[1]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_2_ ( .ip(n4601), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[2]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_4_ ( .ip(n4599), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[4]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_5_ ( .ip(n4598), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[5]) );
  drp_1 i_ssi_U_biu_prdata_reg_7_ ( .ip(n4230), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[7]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_12_ ( .ip(n4607), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[12]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_13_ ( .ip(n4606), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[13]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_14_ ( .ip(n4605), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[14]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_4_ ( .ip(n4585), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr0_ir_int[4]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_5_ ( .ip(n4586), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr0_ir_int[5]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_7_ ( .ip(n4587), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr0_ir_int_7) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_8_ ( .ip(n4588), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_tmod[0]) );
  drp_1 i_ssi_U_biu_prdata_reg_8_ ( .ip(n4229), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[8]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_9_ ( .ip(n4589), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_tmod[1]) );
  drp_1 i_ssi_U_biu_prdata_reg_9_ ( .ip(n4228), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[9]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_10_ ( .ip(n4590), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_ctrlr0[10]) );
  drp_1 i_ssi_U_biu_prdata_reg_10_ ( .ip(n4227), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[10]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_11_ ( .ip(n4591), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_ctrlr0[11]) );
  drp_1 i_ssi_U_biu_prdata_reg_11_ ( .ip(n4226), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[11]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_12_ ( .ip(n4592), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_cfs[0]) );
  drp_1 i_ssi_U_biu_prdata_reg_12_ ( .ip(n4225), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[12]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_13_ ( .ip(n4593), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_cfs[1]) );
  drp_1 i_ssi_U_biu_prdata_reg_13_ ( .ip(n4224), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[13]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_14_ ( .ip(n4594), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_cfs[2]) );
  drp_1 i_ssi_U_biu_prdata_reg_14_ ( .ip(n4223), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[14]) );
  drp_1 i_ssi_U_regfile_ctrlr0_ir_reg_15_ ( .ip(n4595), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_cfs[3]) );
  drp_1 i_ssi_U_biu_prdata_reg_15_ ( .ip(n4222), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[15]) );
  drp_1 i_ssi_U_sclkgen_sclk_fe_ir_reg ( .ip(i_ssi_U_sclkgen_N75), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_sclk_fe) );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_5_ ( .ip(i_ssi_U_sclkgen_N45), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[5])
         );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_6_ ( .ip(i_ssi_U_sclkgen_N46), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[6])
         );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_7_ ( .ip(i_ssi_U_sclkgen_N47), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[7])
         );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_8_ ( .ip(i_ssi_U_sclkgen_N48), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[8])
         );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_10_ ( .ip(i_ssi_U_sclkgen_N50), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[10])
         );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_11_ ( .ip(i_ssi_U_sclkgen_N51), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[11])
         );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_12_ ( .ip(i_ssi_U_sclkgen_N52), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[12])
         );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_13_ ( .ip(i_ssi_U_sclkgen_N53), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[13])
         );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_14_ ( .ip(i_ssi_U_sclkgen_N54), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[14])
         );
  drp_1 i_ssi_U_sclkgen_ssi_cnt_reg_15_ ( .ip(i_ssi_U_sclkgen_N55), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[15])
         );
  drp_1 i_ssi_U_fifo_tx_push_dly_reg ( .ip(n11854), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_fifo_tx_push_dly) );
  drp_1 i_ssi_U_fifo_rx_pop_dly_reg ( .ip(n6937), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_fifo_rx_pop_dly) );
  drp_1 i_ssi_U_mstfsm_U_ss_in_n_sync_sample_meta_reg_0_ ( .ip(i_ssi_ss_in_n), 
        .ck(i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_mstfsm_U_ss_in_n_sync_next_sample_syncm1_0_) );
  drp_1 i_ssi_U_mstfsm_U_ss_in_n_sync_sample_syncl_reg_0_ ( .ip(
        i_ssi_U_mstfsm_U_ss_in_n_sync_next_sample_syncm1_0_), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_ss_in_n_sync)
         );
  drp_1 i_ssi_U_mstfsm_c_state_reg_0_ ( .ip(i_ssi_U_mstfsm_N219), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_c_state[0]) );
  drp_1 i_ssi_U_mstfsm_c_state_reg_1_ ( .ip(i_ssi_U_mstfsm_N220), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_c_state[1]) );
  drp_1 i_ssi_U_mstfsm_c_state_reg_2_ ( .ip(i_ssi_U_mstfsm_N221), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_c_state[2]) );
  drp_1 i_ssi_U_mstfsm_c_state_reg_3_ ( .ip(i_ssi_U_mstfsm_N222), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_c_state[3]) );
  drp_1 i_ssi_U_mstfsm_c_done_ir_reg ( .ip(n11831), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_c_done_ir) );
  drp_1 i_ssi_U_shift_tx_pop_tgl_reg ( .ip(n4578), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_tx_pop) );
  drp_1 i_ssi_U_fifo_tx_pop_edge_reg ( .ip(i_ssi_tx_pop), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_fifo_tx_pop_edge) );
  drp_1 i_ssi_U_fifo_tx_pop_sync_dly_reg ( .ip(i_ssi_tx_pop_sync), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_ssi_U_fifo_tx_pop_sync_dly) );
  drp_1 i_ssi_U_intctl_irisr_tx_empty_reg ( .ip(n10803), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_risr[0]) );
  drp_1 i_ssi_U_intctl_irisr_tx_fifo_overflow_reg ( .ip(n4577), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_ssi_risr[1]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__0_ ( .ip(n4576), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[0]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__1_ ( .ip(n4575), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[1]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__2_ ( .ip(n4574), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[2]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__3_ ( .ip(n4573), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[3]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__4_ ( .ip(n4572), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[4]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__5_ ( .ip(n4571), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[5]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__6_ ( .ip(n4570), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[6]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__7_ ( .ip(n4569), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[7]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__8_ ( .ip(n4568), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[8]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__9_ ( .ip(n4567), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[9]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__10_ ( .ip(n4566), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[10]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__11_ ( .ip(n4565), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[11]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__12_ ( .ip(n4564), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[12]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__13_ ( .ip(n4563), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[13]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__14_ ( .ip(n4562), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[14]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_7__15_ ( .ip(n4561), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[15]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__0_ ( .ip(n4544), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[32]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__1_ ( .ip(n4543), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[33]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__2_ ( .ip(n4542), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[34]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__3_ ( .ip(n4541), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[35]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__4_ ( .ip(n4540), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[36]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__5_ ( .ip(n4539), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[37]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__6_ ( .ip(n4538), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[38]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__7_ ( .ip(n4537), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[39]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__8_ ( .ip(n4536), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[40]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__9_ ( .ip(n4535), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[41]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__10_ ( .ip(n4534), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[42]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__11_ ( .ip(n4533), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[43]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__12_ ( .ip(n4532), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[44]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__13_ ( .ip(n4531), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[45]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__14_ ( .ip(n4530), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[46]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_5__15_ ( .ip(n4529), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[47]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__0_ ( .ip(n4512), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[64]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__1_ ( .ip(n4511), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[65]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__2_ ( .ip(n4510), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[66]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__3_ ( .ip(n4509), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[67]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__4_ ( .ip(n4508), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[68]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__5_ ( .ip(n4507), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[69]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__6_ ( .ip(n4506), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[70]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__7_ ( .ip(n4505), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[71]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__8_ ( .ip(n4504), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[72]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__9_ ( .ip(n4503), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[73]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__10_ ( .ip(n4502), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[74]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__11_ ( .ip(n4501), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[75]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__12_ ( .ip(n4500), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[76]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__13_ ( .ip(n4499), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[77]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__14_ ( .ip(n4498), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[78]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_3__15_ ( .ip(n4497), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[79]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__0_ ( .ip(n4480), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[96]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__1_ ( .ip(n4479), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[97]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__2_ ( .ip(n4478), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[98]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__3_ ( .ip(n4477), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[99]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__4_ ( .ip(n4476), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[100]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__5_ ( .ip(n4475), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[101]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__6_ ( .ip(n4474), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[102]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__7_ ( .ip(n4473), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[103]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__8_ ( .ip(n4472), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[104]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__9_ ( .ip(n4471), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[105]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__10_ ( .ip(n4470), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[106]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__11_ ( .ip(n4469), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[107]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__12_ ( .ip(n4468), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[108]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__13_ ( .ip(n4467), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[109]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__14_ ( .ip(n4466), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[110]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_1__15_ ( .ip(n4465), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[111]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__0_ ( .ip(n4560), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[16]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__1_ ( .ip(n4559), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[17]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__2_ ( .ip(n4558), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[18]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__3_ ( .ip(n4557), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[19]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__4_ ( .ip(n4556), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[20]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__5_ ( .ip(n4555), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[21]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__6_ ( .ip(n4554), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[22]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__7_ ( .ip(n4553), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[23]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__8_ ( .ip(n4552), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[24]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__9_ ( .ip(n4551), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[25]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__10_ ( .ip(n4550), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[26]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__11_ ( .ip(n4549), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[27]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__12_ ( .ip(n4548), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[28]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__13_ ( .ip(n4547), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[29]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__14_ ( .ip(n4546), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[30]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_6__15_ ( .ip(n4545), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[31]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__0_ ( .ip(n4528), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[48]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__1_ ( .ip(n4527), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[49]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__2_ ( .ip(n4526), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[50]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__3_ ( .ip(n4525), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[51]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__4_ ( .ip(n4524), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[52]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__5_ ( .ip(n4523), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[53]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__6_ ( .ip(n4522), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[54]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__7_ ( .ip(n4521), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[55]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__8_ ( .ip(n4520), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[56]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__9_ ( .ip(n4519), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[57]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__10_ ( .ip(n4518), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[58]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__11_ ( .ip(n4517), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[59]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__12_ ( .ip(n4516), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[60]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__13_ ( .ip(n4515), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[61]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__14_ ( .ip(n4514), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[62]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_4__15_ ( .ip(n4513), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[63]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__0_ ( .ip(n4496), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[80]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__1_ ( .ip(n4495), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[81]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__2_ ( .ip(n4494), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[82]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__3_ ( .ip(n4493), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[83]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__4_ ( .ip(n4492), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[84]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__5_ ( .ip(n4491), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[85]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__6_ ( .ip(n4490), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[86]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__7_ ( .ip(n4489), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[87]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__8_ ( .ip(n4488), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[88]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__9_ ( .ip(n4487), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[89]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__10_ ( .ip(n4486), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[90]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__11_ ( .ip(n4485), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[91]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__12_ ( .ip(n4484), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[92]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__13_ ( .ip(n4483), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[93]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__14_ ( .ip(n4482), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[94]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_2__15_ ( .ip(n4481), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[95]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__0_ ( .ip(n4464), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[112]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__1_ ( .ip(n4463), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[113]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__2_ ( .ip(n4462), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[114]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__3_ ( .ip(n4461), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[115]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__4_ ( .ip(n4460), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[116]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__5_ ( .ip(n4459), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[117]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__6_ ( .ip(n4458), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[118]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__7_ ( .ip(n4457), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[119]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__8_ ( .ip(n4456), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[120]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__9_ ( .ip(n4455), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[121]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__10_ ( .ip(n4454), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[122]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__11_ ( .ip(n4453), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[123]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__12_ ( .ip(n4452), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[124]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__13_ ( .ip(n4451), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[125]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__14_ ( .ip(n4450), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[126]) );
  drp_1 i_ssi_U_dff_tx_mem_reg_0__15_ ( .ip(n4449), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_tx_mem[127]) );
  drp_1 i_ssi_U_regfile_txflr_reg_0_ ( .ip(n4447), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_txflr[0]) );
  drp_1 i_ssi_U_regfile_txflr_reg_1_ ( .ip(n4446), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_txflr[1]) );
  drp_1 i_ssi_U_regfile_txflr_reg_2_ ( .ip(n4445), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_txflr[2]) );
  drp_1 i_ssi_U_regfile_txflr_reg_3_ ( .ip(n4448), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_txflr[3]) );
  drp_1 i_ssi_U_mstfsm_last_frame_reg ( .ip(n4422), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_last_frame) );
  drp_1 i_ssi_U_mstfsm_abort_ir_reg ( .ip(n4421), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_abort_ir) );
  drp_1 i_ssi_U_shift_U_tx_shifter_load_start_bit_ir_reg ( .ip(
        i_ssi_load_start_bit), .ck(i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_load_start_bit_ir) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_0_ ( .ip(n4420), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[0]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_1_ ( .ip(n4419), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[1]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_2_ ( .ip(n4418), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[2]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_3_ ( .ip(n4417), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[3]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_4_ ( .ip(n4416), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[4]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_5_ ( .ip(n4415), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[5]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_6_ ( .ip(n4414), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[6]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_7_ ( .ip(n4413), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[7]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_8_ ( .ip(n4412), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[8]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_9_ ( .ip(n4411), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[9]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_10_ ( .ip(n4410), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[10]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_11_ ( .ip(n4409), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[11]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_12_ ( .ip(n4408), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[12]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_13_ ( .ip(n4407), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[13]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_14_ ( .ip(n4406), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[14]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_buffer_reg_15_ ( .ip(n4405), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_buffer[15]) );
  drp_1 i_ssi_U_shift_rx_push_tgl_reg ( .ip(n4444), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_rx_push) );
  drp_1 i_ssi_U_fifo_rx_push_edge_reg ( .ip(i_ssi_rx_push), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_ssi_U_fifo_rx_push_edge) );
  drp_1 i_ssi_U_fifo_rx_push_sync_dly_reg ( .ip(n11837), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_fifo_rx_push_sync_dly) );
  drp_1 i_ssi_U_intctl_irisr_rx_full_reg ( .ip(i_ssi_U_intctl_N33), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_ssi_risr[4]) );
  drp_1 i_ssi_U_biu_prdata_reg_4_ ( .ip(n4233), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[4]) );
  drp_1 i_ssi_U_intctl_irisr_rx_fifo_overflow_reg ( .ip(n4443), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_ssi_risr[3]) );
  drp_1 i_ssi_U_intctl_irisr_rx_fifo_underflow_reg ( .ip(n4442), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(i_ssi_risr[2]) );
  drp_1 i_ssi_U_regfile_rxflr_reg_0_ ( .ip(n4440), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_rxflr[0]) );
  drp_1 i_ssi_U_regfile_rxflr_reg_1_ ( .ip(n4439), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_rxflr[1]) );
  drp_1 i_ssi_U_biu_prdata_reg_1_ ( .ip(n4236), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[1]) );
  drp_1 i_ssi_U_regfile_rxflr_reg_2_ ( .ip(n4438), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_rxflr[2]) );
  drp_1 i_ssi_U_regfile_rxflr_reg_3_ ( .ip(n4441), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_rxflr[3]) );
  drp_1 i_ssi_U_biu_prdata_reg_3_ ( .ip(n4234), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[3]) );
  drp_1 i_ssi_U_biu_prdata_reg_2_ ( .ip(n4235), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[2]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_1_ ( .ip(n4437), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[1]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__1_ ( .ip(n4362), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[1]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__1_ ( .ip(n4361), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[17]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__1_ ( .ip(n4360), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[33]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__1_ ( .ip(n4359), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[49]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__1_ ( .ip(n4358), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[65]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__1_ ( .ip(n4357), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[81]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__1_ ( .ip(n4356), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[97]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__1_ ( .ip(n4355), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[113]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_2_ ( .ip(n4436), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[2]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__2_ ( .ip(n4354), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[2]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__2_ ( .ip(n4353), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[18]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__2_ ( .ip(n4352), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[34]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__2_ ( .ip(n4351), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[50]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__2_ ( .ip(n4350), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[66]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__2_ ( .ip(n4349), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[82]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__2_ ( .ip(n4348), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[98]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__2_ ( .ip(n4347), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[114]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_3_ ( .ip(n4435), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[3]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__3_ ( .ip(n4346), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[3]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__3_ ( .ip(n4345), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[19]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__3_ ( .ip(n4344), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[35]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__3_ ( .ip(n4343), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[51]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__3_ ( .ip(n4342), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[67]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__3_ ( .ip(n4341), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[83]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__3_ ( .ip(n4340), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[99]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__3_ ( .ip(n4339), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[115]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_4_ ( .ip(n4434), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[4]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__4_ ( .ip(n4338), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[4]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__4_ ( .ip(n4337), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[20]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__4_ ( .ip(n4336), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[36]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__4_ ( .ip(n4335), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[52]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__4_ ( .ip(n4334), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[68]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__4_ ( .ip(n4333), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[84]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__4_ ( .ip(n4332), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[100]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__4_ ( .ip(n4331), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[116]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_5_ ( .ip(n4433), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[5]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__5_ ( .ip(n4330), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[5]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__5_ ( .ip(n4329), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[21]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__5_ ( .ip(n4328), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[37]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__5_ ( .ip(n4327), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[53]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__5_ ( .ip(n4326), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[69]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__5_ ( .ip(n4325), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[85]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__5_ ( .ip(n4324), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[101]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__5_ ( .ip(n4323), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[117]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_6_ ( .ip(n4432), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[6]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__6_ ( .ip(n4322), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[6]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__6_ ( .ip(n4321), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[22]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__6_ ( .ip(n4320), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[38]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__6_ ( .ip(n4319), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[54]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__6_ ( .ip(n4318), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[70]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__6_ ( .ip(n4317), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[86]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__6_ ( .ip(n4316), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[102]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__6_ ( .ip(n4315), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[118]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_7_ ( .ip(n4431), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[7]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__7_ ( .ip(n4314), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[7]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__7_ ( .ip(n4313), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[23]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__7_ ( .ip(n4312), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[39]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__7_ ( .ip(n4311), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[55]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__7_ ( .ip(n4310), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[71]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__7_ ( .ip(n4309), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[87]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__7_ ( .ip(n4308), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[103]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__7_ ( .ip(n4307), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[119]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_8_ ( .ip(n4430), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[8]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__8_ ( .ip(n4306), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[8]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__8_ ( .ip(n4305), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[24]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__8_ ( .ip(n4304), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[40]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__8_ ( .ip(n4303), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[56]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__8_ ( .ip(n4302), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[72]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__8_ ( .ip(n4301), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[88]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__8_ ( .ip(n4300), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[104]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__8_ ( .ip(n4299), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[120]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_9_ ( .ip(n4429), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[9]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__9_ ( .ip(n4298), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[9]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__9_ ( .ip(n4297), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[25]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__9_ ( .ip(n4296), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[41]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__9_ ( .ip(n4295), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[57]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__9_ ( .ip(n4294), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[73]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__9_ ( .ip(n4293), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[89]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__9_ ( .ip(n4292), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[105]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__9_ ( .ip(n4291), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[121]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_10_ ( .ip(n4428), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[10]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__10_ ( .ip(n4290), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[10]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__10_ ( .ip(n4289), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[26]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__10_ ( .ip(n4288), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[42]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__10_ ( .ip(n4287), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[58]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__10_ ( .ip(n4286), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[74]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__10_ ( .ip(n4285), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[90]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__10_ ( .ip(n4284), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[106]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__10_ ( .ip(n4283), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[122]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_11_ ( .ip(n4427), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[11]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__11_ ( .ip(n4282), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[11]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__11_ ( .ip(n4281), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[27]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__11_ ( .ip(n4280), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[43]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__11_ ( .ip(n4279), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[59]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__11_ ( .ip(n4278), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[75]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__11_ ( .ip(n4277), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[91]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__11_ ( .ip(n4276), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[107]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__11_ ( .ip(n4275), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[123]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_12_ ( .ip(n4426), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[12]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__12_ ( .ip(n4274), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[12]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__12_ ( .ip(n4273), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[28]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__12_ ( .ip(n4272), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[44]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__12_ ( .ip(n4271), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[60]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__12_ ( .ip(n4270), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[76]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__12_ ( .ip(n4269), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[92]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__12_ ( .ip(n4268), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[108]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__12_ ( .ip(n4267), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[124]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_13_ ( .ip(n4425), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[13]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__13_ ( .ip(n4266), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[13]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__13_ ( .ip(n4265), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[29]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__13_ ( .ip(n4264), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[45]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__13_ ( .ip(n4263), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[61]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__13_ ( .ip(n4262), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[77]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__13_ ( .ip(n4261), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[93]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__13_ ( .ip(n4260), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[109]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__13_ ( .ip(n4259), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[125]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_14_ ( .ip(n4424), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[14]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__14_ ( .ip(n4258), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[14]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__14_ ( .ip(n4257), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[30]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__14_ ( .ip(n4256), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[46]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__14_ ( .ip(n4255), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[62]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__14_ ( .ip(n4254), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[78]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__14_ ( .ip(n4253), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[94]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__14_ ( .ip(n4252), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[110]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__14_ ( .ip(n4251), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[126]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__15_ ( .ip(n4250), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[15]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__15_ ( .ip(n4249), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[31]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__15_ ( .ip(n4248), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[47]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__15_ ( .ip(n4247), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[63]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__15_ ( .ip(n4246), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[79]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__15_ ( .ip(n4245), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[95]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__15_ ( .ip(n4244), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[111]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__15_ ( .ip(n4243), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[127]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_1_ ( .ip(n4402), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[1]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_2_ ( .ip(n4401), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[2]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_3_ ( .ip(n4400), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[3]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_4_ ( .ip(n4399), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[4]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_6_ ( .ip(n4397), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[6]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_7_ ( .ip(n4396), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[7]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_8_ ( .ip(n4395), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[8]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_10_ ( .ip(n4393), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[10]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_12_ ( .ip(n4391), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[12]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_13_ ( .ip(n4390), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[13]) );
  drp_1 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_14_ ( .ip(n4404), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[14]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_0_ ( .ip(n4387), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[0]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_1_ ( .ip(n4386), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[1]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_2_ ( .ip(n4385), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[2]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_3_ ( .ip(n4384), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[3]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_4_ ( .ip(n4383), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[4]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_5_ ( .ip(n4382), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[5]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_6_ ( .ip(n4381), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[6]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_7_ ( .ip(n4380), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[7]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_8_ ( .ip(n4379), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[8]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_9_ ( .ip(n4378), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[9]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_10_ ( .ip(n4377), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[10]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_11_ ( .ip(n4376), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[11]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_12_ ( .ip(n4375), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[12]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_13_ ( .ip(n4374), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[13]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_14_ ( .ip(n4373), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[14]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_shift_reg_reg_15_ ( .ip(n4372), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[15]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_0_ ( .ip(n4371), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[0]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_7__0_ ( .ip(n4370), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[0]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_6__0_ ( .ip(n4369), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[16]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_5__0_ ( .ip(n4368), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[32]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_4__0_ ( .ip(n4367), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[48]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_3__0_ ( .ip(n4366), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[64]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_2__0_ ( .ip(n4365), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[80]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_1__0_ ( .ip(n4364), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[96]) );
  drp_1 i_ssi_U_dff_rx_mem_reg_0__0_ ( .ip(n4363), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_dff_rx_mem[112]) );
  drp_1 i_ssi_U_mstfsm_fsm_sleep_reg ( .ip(n5226), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_fsm_sleep) );
  drp_1 i_ssi_U_regfile_ssi_sleep_ir_reg ( .ip(i_ssi_U_regfile_N451), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_ssi_ssi_sleep) );
  drp_1 i_ssi_U_mstfsm_fsm_busy_reg ( .ip(n11851), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_fsm_busy) );
  drp_1 i_ssi_U_regfile_multi_mst_edge_reg ( .ip(i_ssi_fsm_multi_mst), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_ssi_U_regfile_multi_mst_edge)
         );
  drp_1 i_ssi_U_intctl_irisr_mst_collision_reg ( .ip(n4240), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_ssi_risr[5]) );
  drp_1 i_ssi_U_biu_prdata_reg_0_ ( .ip(n4237), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[0]) );
  drp_1 i_ssi_U_biu_prdata_reg_5_ ( .ip(n4232), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[5]) );
  drp_1 i_ssi_U_intctl_mst_contention_reg ( .ip(n4239), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_mst_contention) );
  drp_1 i_ssi_U_regfile_i_sr_reg ( .ip(n4238), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_sr_6_) );
  drp_1 i_ssi_U_biu_prdata_reg_6_ ( .ip(n4231), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_prdata[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_U_SYNC_sample_meta_reg_0_ ( 
        .ip(i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_U_SYNC_N2), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_U_SYNC_next_sample_syncm1_0_)
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_U_SYNC_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_U_SYNC_next_sample_syncm1_0_), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_data_d_int_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_U_SYNC_sample_meta_reg_0_ ( 
        .ip(i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_U_SYNC_N2), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_U_SYNC_next_sample_syncm1_0_)
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_U_SYNC_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_U_SYNC_next_sample_syncm1_0_), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_data_d_int_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_mst_arb_lost_reg ( .ip(n4932), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_mst_arb_lost) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_12_ ( 
        .ip(i_i2c_tx_abrt_source[12]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_12_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[12]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_12_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[12]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_mst_gen_ack_en_r_reg ( .ip(n11858), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_mst_gen_ack_en_r) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_ic_data_oe_early_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_N85), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_tx_shift_ic_data_oe_early) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_ic_data_oe_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_ic_data_oe_early), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_ic_data_oe) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_ic_rd_req_tog_reg ( .ip(n5030), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ic_rd_req_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_ic_rd_req_flg_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_ic_rd_req_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_ic_rd_req_flg_sync_next_sample_syncm1_0_)
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_ic_rd_req_flg_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_ic_rd_req_flg_sync_next_sample_syncm1_0_), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_ic_rd_req_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_rd_req_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_ic_rd_req_flg_sync), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_DW_apb_i2c_intctl_ic_rd_req_flg_sync_q)
         );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_mst_tx_flush_reg ( .ip(n4857), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_mst_tx_flush) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_sbyte_norstrt_tog_reg ( .ip(n4854), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_9_ ( 
        .ip(i_i2c_tx_abrt_source[9]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[9])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_9_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[9]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_9_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[9]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_9_ ( .ip(n4691), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_gen_call_sample_meta_reg_0_ ( .ip(
        i_i2c_ic_ack_general_call), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_U_DW_apb_i2c_sync_U_ic_gen_call_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_gen_call_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_gen_call_next_sample_syncm1_0_), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ic_ack_general_call_sync)
         );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_ic_sda_hold[0]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[0]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_1_ ( .ip(
        i_i2c_ic_sda_hold[1]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[1]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_2_ ( .ip(
        i_i2c_ic_sda_hold[2]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[2]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_3_ ( .ip(
        i_i2c_ic_sda_hold[3]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_3_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[3]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_4_ ( .ip(
        i_i2c_ic_sda_hold[4]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_4_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[4]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_5_ ( .ip(
        i_i2c_ic_sda_hold[5]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_5_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[5]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_6_ ( .ip(
        i_i2c_ic_sda_hold[6]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_6_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[6]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_7_ ( .ip(
        i_i2c_ic_sda_hold[7]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_7_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[7]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_8_ ( .ip(
        i_i2c_ic_sda_hold[8]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_8_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[8]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_9_ ( .ip(
        i_i2c_ic_sda_hold[9]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_9_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[9]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_10_ ( .ip(
        i_i2c_ic_sda_hold[10]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_10_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[10]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_11_ ( .ip(
        i_i2c_ic_sda_hold[11]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_11_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[11]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_12_ ( .ip(
        i_i2c_ic_sda_hold[12]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_12_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[12]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_13_ ( .ip(
        i_i2c_ic_sda_hold[13]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_13_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[13]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_14_ ( .ip(
        i_i2c_ic_sda_hold[14]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_14_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[14]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_15_ ( .ip(
        i_i2c_ic_sda_hold[15]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_15_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[15]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_tx_hold_sync[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_16_ ( .ip(
        i_i2c_ic_sda_hold[16]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[16]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_16_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[16]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_rx_hold_sync[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_17_ ( .ip(
        i_i2c_ic_sda_hold[17]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[17]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_17_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[17]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_rx_hold_sync[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_18_ ( .ip(
        i_i2c_ic_sda_hold[18]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[18]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_18_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[18]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_rx_hold_sync[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_19_ ( .ip(
        i_i2c_ic_sda_hold[19]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[19]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_19_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[19]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_rx_hold_sync[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_20_ ( .ip(
        i_i2c_ic_sda_hold[20]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[20]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_20_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[20]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_rx_hold_sync[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_21_ ( .ip(
        i_i2c_ic_sda_hold[21]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[21]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_21_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[21]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_rx_hold_sync[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_22_ ( .ip(
        i_i2c_ic_sda_hold[22]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[22]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_22_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[22]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_rx_hold_sync[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_meta_reg_23_ ( .ip(
        i_i2c_ic_sda_hold[23]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[23]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_sample_syncl_reg_23_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_sda_hold_sync_next_sample_syncm1[23]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_ic_sda_rx_hold_sync[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_rstrt_en_1_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_rstrt_en_1_sync_N2), .ck(i_i2c_ic_clk), 
        .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_rstrt_en_1_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_rstrt_en_1_sync_sample_syncl_reg_0_ ( 
        .ip(i_i2c_U_DW_apb_i2c_sync_U_ic_rstrt_en_1_sync_next_sample_syncm1_0_), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_ic_rstrt_en_sync_inv) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_push_dly_reg ( .ip(i_i2c_tx_push), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_push_dly) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_rx_pop_dly_reg ( .ip(i_i2c_rx_pop), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_rx_pop_dly) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_p_det_ifaddr_sample_meta_reg_0_ ( .ip(
        i_i2c_p_det_ifaddr), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_p_det_ifaddr_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_p_det_ifaddr_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_p_det_ifaddr_next_sample_syncm1_0_), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_p_det_ifaddr_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_slave_en_1_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_ic_slave_en), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_slave_en_1_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_slave_en_1_sync_sample_syncl_reg_0_ ( 
        .ip(i_i2c_U_DW_apb_i2c_sync_U_ic_slave_en_1_sync_next_sample_syncm1_0_), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ic_slave_en_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_slv_1_sync_sample_meta_reg_0_ ( 
        .ip(n11868), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_slv_1_sync_next_sample_syncm1_0_)
         );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_slv_1_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_slv_1_sync_next_sample_syncm1_0_), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_ic_10bit_slv_sync_inv) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_mst_1_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_mst_1_sync_N2), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_mst_1_sync_next_sample_syncm1_0_)
         );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_mst_1_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_mst_1_sync_next_sample_syncm1_0_), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_ic_10bit_mst_sync_inv) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_master_1_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_master_1_sync_N2), .ck(i_i2c_ic_clk), 
        .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_master_1_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_master_1_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_master_1_sync_next_sample_syncm1_0_), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_master_dis_tog_reg ( .ip(n4855), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_11_ ( 
        .ip(i_i2c_tx_abrt_source[11]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_11_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[11]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_11_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[11]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_ss_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_ic_ss), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_ss_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_fs_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_ic_fs), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_fs_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_fs_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_fs_sync_next_sample_syncm1_0_), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ic_fs_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_hs_sync_sample_meta_reg_0_ ( .ip(n11840), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_hs_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_hs_norstrt_tog_reg ( .ip(n4856), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_8_ ( 
        .ip(i_i2c_tx_abrt_source[8]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[8])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_8_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[8]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_8_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[8]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_enable_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_ic_enable[0]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_enable_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_enable_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_enable_sync_next_sample_syncm1_0_), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ic_enable_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_ic_bus_idle_reg ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N51), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ic_bus_idle) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_abort_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_ic_enable[1]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_ic_abort_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_abort_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_abort_sync_next_sample_syncm1_0_), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ic_abort_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_sync_d_reg ( .ip(
        i_i2c_ic_abort_sync), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_sync_d) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_split_start_en_int_reg ( .ip(n5225), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_split_start_en) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_start_en_int_reg ( .ip(n5110), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_start_en) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_st_scl_s_hld_en_reg ( .ip(i_i2c_start_en), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_st_scl_s_hld_en) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cmplt_reg ( .ip(n5188), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_scl_s_hld_cmplt) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl_lcnt_en_reg ( .ip(n4955), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl_lcnt_en) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_lcnt_cmplt_reg ( .ip(n8523), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_scl_lcnt_cmplt) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_re_start_en_int_reg ( .ip(n5192), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_re_start_en) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_s_gen_reg ( .ip(
        i_i2c_U_DW_apb_i2c_toggle_N30), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_s_gen) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_byte_wait_scl_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_byte_wait_en), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_byte_wait_scl) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_rd_reg ( .ip(n11863), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_debug_rd) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_bit_count_reg_1_ ( .ip(n5108), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_mst_rx_bit_count[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_ack_int_reg ( .ip(n4952), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_mst_rx_ack_vld) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rxbyte_rdy_reg ( .ip(n4931), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_mst_rxbyte_rdy) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_byte_waiting_q_reg ( .ip(n5184), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_byte_waiting_q) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_mst_current_state_reg_3_ ( .ip(
        i_i2c_U_DW_apb_i2c_mstfsm_N75), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_mst_debug_cstate[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_mst_cstate_reg_3_ ( .ip(
        i_i2c_mst_debug_cstate[3]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_mst_cstate[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_mst_activity_reg ( .ip(
        i_i2c_U_DW_apb_i2c_mstfsm_N487), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_mst_activity) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_master_act_reg ( .ip(
        i_i2c_mst_activity), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_debug_master_act) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_mst_activity_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_mst_activity), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_mst_activity_sync_next_sample_syncm1_0_)
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_mst_activity_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_mst_activity_sync_next_sample_syncm1_0_), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_mst_activity_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_mst_current_state_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_mstfsm_N72), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_mst_debug_cstate[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_mst_cstate_reg_0_ ( .ip(
        i_i2c_mst_debug_cstate[0]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_mst_cstate[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_mst_cstate_reg_1_ ( .ip(
        i_i2c_mst_debug_cstate[1]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_mst_cstate[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_mst_cstate_reg_2_ ( .ip(
        i_i2c_mst_debug_cstate[2]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_mst_cstate[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_addr_2byte_sent_reg ( .ip(n5199), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_addr_2byte_sent) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_pop_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_tx_pop) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_pop_flg_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_tx_pop_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_pop_flg_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_pop_flg_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_pop_flg_sync_next_sample_syncm1_0_), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_pop_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_pop_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_tx_pop_flg_sync), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_DW_apb_i2c_fifo_tx_pop_flg_sync_q) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_pop_sync_dly_reg ( .ip(i_i2c_tx_pop_sync), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_pop_sync_dly) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_tx_empty_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_empty_n), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_U_tx_empty_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_tx_empty_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_tx_empty_sync_next_sample_syncm1_0_), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_tx_empty_int_inv) );
  drp_1 i_i2c_U_dff_tx_mem_reg_7__0_ ( .ip(n5028), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[0]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_7__1_ ( .ip(n5020), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[1]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_7__2_ ( .ip(n5012), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[2]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_7__3_ ( .ip(n5004), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[3]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_7__4_ ( .ip(n4996), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[4]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_7__5_ ( .ip(n4988), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[5]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_7__6_ ( .ip(n4980), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[6]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_7__7_ ( .ip(n4972), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[7]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_7__8_ ( .ip(n4964), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[8]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_5__0_ ( .ip(n5026), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[18]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_5__1_ ( .ip(n5018), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[19]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_5__2_ ( .ip(n5010), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[20]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_5__3_ ( .ip(n5002), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[21]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_5__4_ ( .ip(n4994), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[22]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_5__5_ ( .ip(n4986), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[23]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_5__6_ ( .ip(n4978), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[24]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_5__7_ ( .ip(n4970), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[25]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_5__8_ ( .ip(n4962), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[26]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_3__0_ ( .ip(n5024), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[36]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_3__1_ ( .ip(n5016), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[37]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_3__2_ ( .ip(n5008), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[38]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_3__3_ ( .ip(n5000), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[39]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_3__4_ ( .ip(n4992), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[40]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_3__5_ ( .ip(n4984), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[41]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_3__6_ ( .ip(n4976), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[42]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_3__7_ ( .ip(n4968), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[43]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_3__8_ ( .ip(n4960), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[44]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_1__0_ ( .ip(n5022), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[54]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_1__1_ ( .ip(n5014), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[55]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_1__2_ ( .ip(n5006), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[56]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_1__3_ ( .ip(n4998), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[57]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_1__4_ ( .ip(n4990), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[58]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_1__5_ ( .ip(n4982), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[59]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_1__6_ ( .ip(n4974), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[60]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_1__7_ ( .ip(n4966), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[61]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_1__8_ ( .ip(n4958), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[62]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_6__0_ ( .ip(n5027), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[9]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_6__1_ ( .ip(n5019), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[10]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_6__2_ ( .ip(n5011), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[11]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_6__3_ ( .ip(n5003), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[12]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_6__4_ ( .ip(n4995), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[13]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_6__5_ ( .ip(n4987), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[14]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_6__6_ ( .ip(n4979), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[15]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_6__7_ ( .ip(n4971), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[16]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_6__8_ ( .ip(n4963), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[17]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_4__0_ ( .ip(n5025), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[27]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_4__1_ ( .ip(n5017), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[28]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_4__2_ ( .ip(n5009), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[29]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_4__3_ ( .ip(n5001), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[30]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_4__4_ ( .ip(n4993), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[31]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_4__5_ ( .ip(n4985), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[32]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_4__6_ ( .ip(n4977), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[33]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_4__7_ ( .ip(n4969), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[34]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_4__8_ ( .ip(n4961), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[35]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_2__0_ ( .ip(n5023), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[45]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_2__1_ ( .ip(n5015), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[46]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_2__2_ ( .ip(n5007), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[47]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_2__3_ ( .ip(n4999), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[48]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_2__4_ ( .ip(n4991), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[49]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_2__5_ ( .ip(n4983), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[50]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_2__6_ ( .ip(n4975), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[51]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_2__7_ ( .ip(n4967), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[52]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_2__8_ ( .ip(n4959), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[53]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_0__0_ ( .ip(n5021), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[63]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_0__1_ ( .ip(n5013), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[64]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_0__2_ ( .ip(n5005), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[65]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_0__3_ ( .ip(n4997), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[66]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_0__4_ ( .ip(n4989), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[67]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_0__5_ ( .ip(n4981), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[68]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_0__6_ ( .ip(n4973), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[69]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_0__7_ ( .ip(n4965), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[70]) );
  drp_1 i_i2c_U_dff_tx_mem_reg_0__8_ ( .ip(n4957), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_tx_mem[71]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_fifo_data_buf_reg_0_ ( .ip(n5222), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_fifo_data_buf[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_fifo_data_buf_reg_1_ ( .ip(n5221), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_fifo_data_buf[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_fifo_data_buf_reg_2_ ( .ip(n5220), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_fifo_data_buf[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_fifo_data_buf_reg_3_ ( .ip(n5219), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_fifo_data_buf[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_fifo_data_buf_reg_4_ ( .ip(n5218), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_fifo_data_buf[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_fifo_data_buf_reg_5_ ( .ip(n5217), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_fifo_data_buf[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_fifo_data_buf_reg_6_ ( .ip(n5216), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_fifo_data_buf[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_fifo_data_buf_reg_7_ ( .ip(n5215), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_fifo_data_buf[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_fifo_data_buf_reg_8_ ( .ip(n5214), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_fifo_data_buf[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_data_capture_reg ( .ip(n11834), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_debug_wr) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_scl_p_stp_int_reg ( .ip(n5061), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_scl_p_setup_en) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cmplt_reg ( .ip(n5044), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_scl_p_setup_cmplt) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_mst_current_state_reg_4_ ( .ip(
        i_i2c_U_DW_apb_i2c_mstfsm_N76), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_mst_debug_cstate[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_mst_cstate_reg_4_ ( .ip(
        i_i2c_mst_debug_cstate[4]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_mst_cstate[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_abrt_in_rcve_trns_reg ( .ip(n5183), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_abrt_in_rcve_trns) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_addr_1byte_sent_reg ( .ip(n5200), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_addr_1byte_sent) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_delay_stop_en_reg ( .ip(
        i_i2c_U_DW_apb_i2c_mstfsm_N421), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_mstfsm_delay_stop_en) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_p_gen_reg ( .ip(n11857), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_debug_p_gen) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_old_is_read_reg ( .ip(n5201), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_old_is_read) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_hs_mcode_en_r_reg ( .ip(n5562), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_hs_mcode_en_r) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_hs_mcode_fed_dtctd_r_reg ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N50), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_hs_mcode_fed_dtctd_r)
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt_reg_0_ ( .ip(n11865), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N83), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[1])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt_reg_3_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N85), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[3])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt_reg_7_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N89), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[7])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N123), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[0])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N124), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[1])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N125), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[2])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt_reg_3_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N126), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[3])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt_reg_4_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N127), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[4])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt_reg_5_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N128), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[5])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt_reg_6_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N129), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[6])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt_reg_7_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N130), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[7])
         );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_int_d_reg ( .ip(n6352), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_int_d) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_p_det_reg ( .ip(n11864), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_p_det) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_sda_vld_int_reg ( .ip(n5227), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_sda_vld) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_s_det_reg ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_s_det_int), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_s_det) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_s_det_flg_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_s_det_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_s_det_flg_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_s_det_flg_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_s_det_flg_sync_next_sample_syncm1_0_), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_s_det_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_s_det_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_s_det_flg_sync), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_DW_apb_i2c_intctl_s_det_flg_sync_q) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N62), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N63), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N64), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_3_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N65), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_4_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N66), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_5_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N67), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_6_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N68), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_7_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N69), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_8_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N70), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_9_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N71), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_10_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N72), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_11_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N73), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_13_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N75), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_15_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N77), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt_reg_0_ ( .ip(n5096), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt_reg_1_ ( .ip(n5095), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt_reg_2_ ( .ip(n5094), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt_reg_3_ ( .ip(n5093), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt_reg_4_ ( .ip(n5092), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt_reg_5_ ( .ip(n5091), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt_reg_6_ ( .ip(n5090), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt_reg_7_ ( .ip(n5089), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_scl_edg_hl_q_reg ( .ip(n11835), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_scl_edg_hl_q) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_qq_reg ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_q), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_qq) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count_reg_3_ ( .ip(n5098), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_cmplt_reg ( .ip(n8091), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_tx_cmplt) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_current_state_reg_0_ ( .ip(n9603), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_debug_cstate[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_slv_cstate_reg_0_ ( .ip(
        i_i2c_slv_debug_cstate[0]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_slv_cstate[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly1_reg ( .ip(n11859), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly1) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ack_vld_reg ( .ip(n5104), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_tx_ack_vld) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_slv_ack_det_reg ( .ip(n5065), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_ack_det) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_rx_done_tog_reg ( .ip(n5064), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_done_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_rx_done_flg_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_rx_done_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_rx_done_flg_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_rx_done_flg_sync_sample_syncl_reg_0_ ( 
        .ip(i_i2c_U_DW_apb_i2c_intctl_U_rx_done_flg_sync_next_sample_syncm1_0_), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_rx_done_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_rx_done_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_rx_done_flg_sync), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_DW_apb_i2c_intctl_rx_done_flg_sync_q) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_tx_flush_reg ( .ip(n5223), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_slv_tx_flush) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_current_state_reg_3_ ( .ip(
        i_i2c_U_DW_apb_i2c_slvfsm_N39), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_slv_debug_cstate[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_slv_cstate_reg_3_ ( .ip(
        i_i2c_slv_debug_cstate[3]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_slv_cstate[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_current_state_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_slvfsm_N38), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_slv_debug_cstate[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_slv_cstate_reg_2_ ( .ip(
        i_i2c_slv_debug_cstate[2]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_slv_cstate[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_data_reg ( .ip(
        i_i2c_U_DW_apb_i2c_toggle_N31), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_data) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_reg_0_ ( .ip(n5077), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_reg_1_ ( .ip(n5076), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_reg_2_ ( .ip(n5075), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_reg_3_ ( .ip(n5074), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_3_) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg_reg_0_ ( .ip(n5073), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg_reg_2_ ( .ip(n5071), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg_reg_4_ ( .ip(n5069), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg_reg_6_ ( .ip(n5067), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg_reg_1_ ( .ip(n5072), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg_reg_3_ ( .ip(n5070), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg_reg_5_ ( .ip(n5068), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg_reg_7_ ( .ip(n5066), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_gen_call_reg ( .ip(n5084), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_gen_call) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_rx_gen_call_r_reg ( .ip(i_i2c_rx_gen_call), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_toggle_rx_gen_call_r) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_rx_gen_call_flg_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_rx_gen_call_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_rx_gen_call_flg_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_rx_gen_call_flg_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_rx_gen_call_flg_sync_next_sample_syncm1_0_), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync_q)
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_hs_mcode_reg ( .ip(n5083), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_hs_mcode) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_rx_hs_mcode_r_reg ( .ip(i_i2c_rx_hs_mcode), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_rx_hs_mcode_r) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_addr_10bit_reg ( .ip(n5086), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_addr_10bit) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_addr_10bit_reg ( .ip(
        i_i2c_rx_addr_10bit), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_debug_addr_10bit) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_slv_read_reg ( .ip(
        i_i2c_U_DW_apb_i2c_rx_shift_rx_slv_read_s), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_rx_slv_read) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_addr_match_reg ( .ip(n5085), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_addr_match) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_current_state_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_slvfsm_N37), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_slv_debug_cstate[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_slv_cstate_reg_1_ ( .ip(
        i_i2c_slv_debug_cstate[1]), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_slv_cstate[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_rx_2addr_reg ( .ip(n5224), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_rx_2addr) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rxbyte_rdy_reg ( .ip(n9563), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_rxbyte_rdy) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_addr_reg ( .ip(
        i_i2c_U_DW_apb_i2c_toggle_N32), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_addr) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_activity_reg ( .ip(
        i_i2c_U_DW_apb_i2c_slvfsm_N284), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_activity) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_slave_act_reg ( .ip(i_i2c_slv_activity), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_debug_slave_act) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_slv_activity_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_slv_activity), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_slv_activity_sync_next_sample_syncm1_0_)
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_slv_activity_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_slv_activity_sync_next_sample_syncm1_0_), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_slv_activity_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_en_reg ( .ip(i_i2c_U_DW_apb_i2c_intctl_N4), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_en) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_empty_intr_reg ( .ip(
        i_i2c_ic_intr_stat[4]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_tx_empty_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_slvrd_intx_tog_reg ( .ip(n5111), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_15_ ( 
        .ip(i_i2c_tx_abrt_source[15]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_15_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[15]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_15_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[15]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_rx_aborted_reg ( .ip(n5203), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_rx_aborted) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_slv_rx_aborted_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_slv_rx_aborted), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_slv_rx_aborted_sync_next_sample_syncm1_0_)
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_slv_rx_aborted_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_slv_rx_aborted_sync_next_sample_syncm1_0_), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_slv_rx_aborted_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_push_reg ( .ip(
        i_i2c_U_DW_apb_i2c_rx_shift_N30), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_rx_push) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_push_flg_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_rx_push_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_push_flg_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_push_flg_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_push_flg_sync_next_sample_syncm1_0_), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_rx_push_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_rx_push_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_rx_push_flg_sync), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_DW_apb_i2c_fifo_rx_push_flg_sync_q) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_rx_push_sync_dly_reg ( .ip(i_i2c_rx_push_sync), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_rx_push_sync_dly) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_rx_full_intr_reg ( .ip(
        i_i2c_ic_intr_stat[2]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_rx_full_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_fifo_filled_and_flushed_reg ( .ip(n5079), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_slv_fifo_filled_and_flushed) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_slv_fifo_filled_and_flushed_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_slv_fifo_filled_and_flushed), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_slv_fifo_filled_and_flushed_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_slv_fifo_filled_and_flushed_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_slv_fifo_filled_and_flushed_sync_next_sample_syncm1_0_), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_slv_fifo_filled_and_flushed_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_slv_addressed_reg ( .ip(n5078), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_addressed) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_p_det_intr_reg ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N241), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_p_det_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_p_det_flg_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_p_det_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_p_det_flg_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_p_det_flg_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_p_det_flg_sync_next_sample_syncm1_0_), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_p_det_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_p_det_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_p_det_flg_sync), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_DW_apb_i2c_intctl_p_det_flg_sync_q) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_ack_vld_reg ( .ip(n5082), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_rx_ack_vld) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_ic_enable_sync_vld_reg ( .ip(n5081), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_ic_enable_sync_vld) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count_reg_0_ ( .ip(n5211), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count_reg_1_ ( .ip(n5210), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count_reg_2_ ( .ip(n5209), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count_reg_3_ ( .ip(n5208), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count_reg_4_ ( .ip(n5207), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count_reg_5_ ( .ip(n5206), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count_reg_6_ ( .ip(n5205), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count_reg_7_ ( .ip(n5204), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_scl_hld_low_en_r_reg ( .ip(
        i_i2c_scl_hld_low_en), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_scl_hld_low_en_r) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_tx_abrt_r_reg ( .ip(
        i_i2c_U_DW_apb_i2c_toggle_tx_abrt), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_toggle_tx_abrt_r) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_tx_abrt_tog_reg ( .ip(n5196), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_flg_sync_sample_meta_reg_0_ ( .ip(
        i_i2c_tx_abrt_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_flg_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_flg_sync_sample_syncl_reg_0_ ( 
        .ip(i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_flg_sync_next_sample_syncm1_0_), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_flg_sync), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_flg_sync_q) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_slvflush_txfifo_tog_reg ( .ip(n5032), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[13])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_13_ ( 
        .ip(i_i2c_tx_abrt_source[13]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_13_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[13]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_13_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[13]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_slv_clr_leftover_tog_reg ( .ip(n5031), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_slv_clr_leftover_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_slv_clr_leftover_flg_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_slv_clr_leftover_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_slv_clr_leftover_flg_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_slv_clr_leftover_flg_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_slv_clr_leftover_flg_sync_next_sample_syncm1_0_), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_slv_clr_leftover_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_slv_clr_leftover_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_slv_clr_leftover_flg_sync), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_slv_clr_leftover_flg_sync_q) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly2_reg ( .ip(n11860), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly2) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_N402), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_slv_tx_ready_unconn) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count_reg_0_ ( .ip(n5101), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count_reg_1_ ( .ip(n5100), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count_reg_2_ ( .ip(n5099), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_debug_hs_reg ( .ip(
        i_i2c_U_DW_apb_i2c_toggle_N33), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_debug_hs) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_15_ ( .ip(n5128), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_1_ ( .ip(n5126), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_2_ ( .ip(n5125), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_3_ ( .ip(n5124), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_4_ ( .ip(n5123), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_5_ ( .ip(n5122), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_7_ ( .ip(n5120), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_8_ ( .ip(n5119), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_9_ ( .ip(n5118), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_10_ ( .ip(n5117), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_11_ ( .ip(n5116), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_12_ ( .ip(n5115), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_13_ ( .ip(n5114), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_14_ ( .ip(n5113), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cmplt_reg ( .ip(n5112), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_mstfsm_N382)
         );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_15_ ( .ip(n5060), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_0_ ( .ip(n5059), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_1_ ( .ip(n5058), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_2_ ( .ip(n5057), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_3_ ( .ip(n5056), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_4_ ( .ip(n5055), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_5_ ( .ip(n5054), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_6_ ( .ip(n5053), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_7_ ( .ip(n5052), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_8_ ( .ip(n5051), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_9_ ( .ip(n5050), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_10_ ( .ip(n5049), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_11_ ( .ip(n5048), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_12_ ( .ip(n5047), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_13_ ( .ip(n5046), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr_reg_14_ ( .ip(n5045), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_stop_scl_lcnt_en_reg ( .ip(n5041), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_stop_scl_lcnt_en) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_hs_ackdet_tog_reg ( .ip(n5182), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_6_ ( 
        .ip(i_i2c_tx_abrt_source[6]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[6])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_6_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[6]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_6_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[6]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_sbyte_ackdet_tog_reg ( .ip(n5180), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_7_ ( 
        .ip(i_i2c_tx_abrt_source[7]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[7])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_7_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[7]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_7_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[7]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_7b_addr_noack_tog_reg ( .ip(n5187), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_tx_abrt_source[0]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[0])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[0]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[0]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_txdata_noack_tog_reg ( .ip(n5186), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_3_ ( 
        .ip(i_i2c_tx_abrt_source[3]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[3])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_3_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[3]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_3_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[3]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_10addr1_noack_tog_reg ( .ip(n5185), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_1_ ( 
        .ip(i_i2c_tx_abrt_source[1]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[1])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_1_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[1]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[1]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_10addr2_noack_tog_reg ( .ip(n5181), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_2_ ( 
        .ip(i_i2c_tx_abrt_source[2]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[2])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_2_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[2]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[2]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_gcall_noack_tog_reg ( .ip(n5179), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_4_ ( 
        .ip(i_i2c_tx_abrt_source[4]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[4])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_4_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[4]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_4_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[4]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_10b_rd_norstrt_tog_reg ( .ip(n5202), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[10])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_10_ ( 
        .ip(i_i2c_tx_abrt_source[10]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_10_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[10]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_10_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[10]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_slv_arblost_tog_reg ( .ip(n5213), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_14_ ( 
        .ip(i_i2c_tx_abrt_source[14]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_14_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[14]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_14_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[14]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf_reg_0_ ( .ip(n5040), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf_reg_1_ ( .ip(n5039), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf_reg_2_ ( .ip(n5038), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf_reg_3_ ( .ip(n5037), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf_reg_4_ ( .ip(n5036), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf_reg_5_ ( .ip(n5035), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf_reg_6_ ( .ip(n5034), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf_reg_7_ ( .ip(n5033), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_tx_empty_hld_reg ( .ip(n5029), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_tx_empty_hld) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_user_abrt_tog_reg ( .ip(n5198), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[16]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_16_ ( 
        .ip(i_i2c_tx_abrt_source[16]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[16]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_16_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[16]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[16]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_16_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[16]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[16]) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_abrt_in_idle_reg ( .ip(n5197), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_abrt_in_idle) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_scl_lcnt_en_reg ( .ip(n5194), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_scl_lcnt_en) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_bit_count_reg_0_ ( .ip(n5109), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_mst_rx_bit_count[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_bit_count_reg_2_ ( .ip(n5107), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_mst_rx_bit_count[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_bit_count_reg_3_ ( .ip(n5106), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_mst_rx_bit_count[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_current_src_en_reg ( .ip(n5063), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_current_src_en) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_scl_hcnt_en_reg ( .ip(n5195), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_scl_hcnt_en) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_set_tx_empty_en_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_N74), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_set_tx_empty_en) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_set_tx_empty_en_flg_sync_sample_meta_reg_0_ ( 
        .ip(i_i2c_set_tx_empty_en_flg), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_set_tx_empty_en_flg_sync_next_sample_syncm1_0_) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_set_tx_empty_en_flg_sync_sample_syncl_reg_0_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_set_tx_empty_en_flg_sync_next_sample_syncm1_0_), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_set_tx_empty_en_flg_sync) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_set_tx_empty_en_flg_sync_q_reg ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_set_tx_empty_en_flg_sync), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_set_tx_empty_en_flg_sync_q) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_current_src_en_reg ( .ip(n5062), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_current_src_en) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_ic_current_src_en_reg ( .ip(
        i_i2c_U_DW_apb_i2c_toggle_N29), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_ic_current_src_en) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en_reg_0_ ( 
        .ip(i_i2c_U_DW_apb_i2c_rx_filter_N207), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[0])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en_reg_1_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[0]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[1])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en_reg_2_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[1]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[2])
         );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en_reg_3_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[2]), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[3])
         );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_scl_s_stp_int_reg ( .ip(n5191), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_scl_s_setup_en) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cmplt_reg ( .ip(n5190), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_scl_s_setup_cmplt) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_0_ ( .ip(n5146), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_1_ ( .ip(n5145), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_2_ ( .ip(n5144), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_3_ ( .ip(n5143), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_4_ ( .ip(n5142), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_5_ ( .ip(n5141), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_6_ ( .ip(n5140), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_7_ ( .ip(n5139), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_8_ ( .ip(n5138), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_10_ ( .ip(n5136), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_11_ ( .ip(n5135), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_12_ ( .ip(n5134), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_13_ ( .ip(n5133), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_14_ ( .ip(n5132), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_15_ ( .ip(n7160), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_re_scl_s_hld_en_reg ( .ip(n5189), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_re_scl_s_hld_en) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_abrt_gcall_read_tog_reg ( .ip(n4933), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_meta_reg_5_ ( 
        .ip(i_i2c_tx_abrt_source[5]), .ck(PCLK_pclk), .rb(PRESETn_presetn), 
        .q(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[5])
         );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_sample_syncl_reg_5_ ( 
        .ip(
        i_i2c_U_DW_apb_i2c_intctl_U_tx_abrt_source_sync_next_sample_syncm1[5]), 
        .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q_reg_5_ ( .ip(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[5]), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_0_ ( .ip(n5178), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_1_ ( .ip(n5177), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_2_ ( .ip(n5176), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_3_ ( .ip(n5175), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_4_ ( .ip(n5174), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_5_ ( .ip(n5173), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_6_ ( .ip(n5172), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_7_ ( .ip(n5171), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_8_ ( .ip(n5170), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_9_ ( .ip(n5169), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_10_ ( .ip(n5168), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_11_ ( .ip(n5167), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_12_ ( .ip(n5166), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_13_ ( .ip(n5165), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_14_ ( .ip(n5164), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr_reg_15_ ( .ip(n5163), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_0_ ( .ip(n5162), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_1_ ( .ip(n5161), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_2_ ( .ip(n5160), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_3_ ( .ip(n5159), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_4_ ( .ip(n5158), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_5_ ( .ip(n5157), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_6_ ( .ip(n5156), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_7_ ( .ip(n5155), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_8_ ( .ip(n5154), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_9_ ( .ip(n5153), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_11_ ( .ip(n5151), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_12_ ( .ip(n5150), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_13_ ( .ip(n5149), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_14_ ( .ip(n5148), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_15_ ( .ip(n5147), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_ic_clk_oe_reg ( .ip(n4951), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ic_clk_oe) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_0_ ( .ip(n4950), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_1_ ( .ip(n4949), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_2_ ( .ip(n4948), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_3_ ( .ip(n4947), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_4_ ( .ip(n4946), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_6_ ( .ip(n4944), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_7_ ( .ip(n4943), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_8_ ( .ip(n4942), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_14_ ( .ip(n4936), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_start_sda_gate_r_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_N272), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_tx_shift_start_sda_gate_r) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_mst_slv_ack_ext_r_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_mst_slv_ack_ext), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_tx_shift_mst_slv_ack_ext_r) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_gen_call_reg ( .ip(n4653), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_gen_call_intr_reg ( .ip(
        i_i2c_ic_intr_stat[11]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_gen_call_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_activity_reg ( .ip(n4650), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_activity_intr_reg ( .ip(
        i_i2c_ic_intr_stat[8]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_activity_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_stop_det_reg ( .ip(n4652), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_stop_det_intr_reg ( .ip(
        i_i2c_ic_intr_stat[9]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_stop_det_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_start_det_reg ( .ip(n4651), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_start_det_intr_reg ( .ip(
        i_i2c_ic_intr_stat[10]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_start_det_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_rx_done_reg ( .ip(n4649), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_rx_done_intr_reg ( .ip(
        i_i2c_ic_intr_stat[7]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_rx_done_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_16_ ( .ip(n5212), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[16]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_0_ ( .ip(n4700), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_1_ ( .ip(n4699), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_2_ ( .ip(n4698), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_3_ ( .ip(n4697), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_4_ ( .ip(n4696), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_5_ ( .ip(n4695), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_6_ ( .ip(n4694), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_7_ ( .ip(n4693), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_8_ ( .ip(n4692), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_10_ ( .ip(n4690), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_11_ ( .ip(n4689), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_12_ ( .ip(n4688), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_13_ ( .ip(n4687), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_14_ ( .ip(n4686), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_source_reg_15_ ( .ip(n4685), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_tx_abrt_source[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_tx_abrt_reg ( .ip(n4648), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_abrt_intr_reg ( .ip(
        i_i2c_ic_intr_stat[6]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_tx_abrt_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_rd_req_reg ( .ip(n4647), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_rd_req_intr_reg ( .ip(
        i_i2c_ic_intr_stat[5]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_rd_req_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_rx_under_reg ( .ip(n4646), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_rx_under_intr_reg ( .ip(
        i_i2c_ic_intr_stat[0]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_rx_under_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_rx_over_reg ( .ip(n4645), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_rx_over_intr_reg ( .ip(
        i_i2c_ic_intr_stat[1]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_rx_over_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_raw_tx_over_reg ( .ip(n4644), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_ic_raw_intr_stat[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_intctl_ic_tx_over_intr_reg ( .ip(
        i_i2c_ic_intr_stat[3]), .ck(PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_ic_tx_over_intr) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_0_ ( .ip(n4654), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_1_ ( .ip(n4655), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_2_ ( .ip(n4656), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_3_ ( .ip(n4657), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_4_ ( .ip(n4658), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_5_ ( .ip(n4659), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_6_ ( .ip(n4660), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_7_ ( .ip(n4661), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_8_ ( .ip(n4662), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_9_ ( .ip(n4663), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_10_ ( .ip(n4664), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_11_ ( .ip(n4665), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_12_ ( .ip(n4666), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_13_ ( .ip(n4667), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_14_ ( .ip(n4668), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_15_ ( .ip(n4669), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_16_ ( .ip(n4670), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[16]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_17_ ( .ip(n4671), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[17]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_18_ ( .ip(n4672), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[18]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_19_ ( .ip(n4673), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[19]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_20_ ( .ip(n4674), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[20]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_21_ ( .ip(n4675), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[21]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_22_ ( .ip(n4676), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[22]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_23_ ( .ip(n4677), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[23]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_24_ ( .ip(n4678), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[24]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_25_ ( .ip(n4679), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[25]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_26_ ( .ip(n4680), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[26]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_28_ ( .ip(n4682), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[28]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_29_ ( .ip(n4683), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[29]) );
  drp_1 i_i2c_U_DW_apb_i2c_biu_prdata_reg_30_ ( .ip(n4684), .ck(PCLK_pclk), 
        .rb(PRESETn_presetn), .q(i_i2c_prdata[30]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg_reg_0_ ( .ip(n4929), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[0]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_7__0_ ( .ip(n4921), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[0]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_6__0_ ( .ip(n4920), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[8]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_5__0_ ( .ip(n4919), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[16]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_4__0_ ( .ip(n4918), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[24]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_3__0_ ( .ip(n4917), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[32]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_2__0_ ( .ip(n4916), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[40]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_1__0_ ( .ip(n4915), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[48]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_0__0_ ( .ip(n4914), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[56]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg_reg_1_ ( .ip(n4928), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[1]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_7__1_ ( .ip(n4913), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[1]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_6__1_ ( .ip(n4912), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[9]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_5__1_ ( .ip(n4911), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[17]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_4__1_ ( .ip(n4910), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[25]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_3__1_ ( .ip(n4909), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[33]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_2__1_ ( .ip(n4908), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[41]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_1__1_ ( .ip(n4907), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[49]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_0__1_ ( .ip(n4906), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[57]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg_reg_2_ ( .ip(n4927), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[2]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_7__2_ ( .ip(n4905), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[2]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_6__2_ ( .ip(n4904), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[10]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_5__2_ ( .ip(n4903), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[18]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_4__2_ ( .ip(n4902), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[26]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_3__2_ ( .ip(n4901), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[34]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_2__2_ ( .ip(n4900), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[42]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_1__2_ ( .ip(n4899), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[50]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_0__2_ ( .ip(n4898), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[58]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg_reg_3_ ( .ip(n4926), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[3]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_7__3_ ( .ip(n4897), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[3]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_6__3_ ( .ip(n4896), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[11]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_5__3_ ( .ip(n4895), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[19]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_4__3_ ( .ip(n4894), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[27]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_3__3_ ( .ip(n4893), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[35]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_2__3_ ( .ip(n4892), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[43]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_1__3_ ( .ip(n4891), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[51]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_0__3_ ( .ip(n4890), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[59]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg_reg_4_ ( .ip(n4925), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[4]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_7__4_ ( .ip(n4889), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[4]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_6__4_ ( .ip(n4888), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[12]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_5__4_ ( .ip(n4887), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[20]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_4__4_ ( .ip(n4886), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[28]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_3__4_ ( .ip(n4885), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[36]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_2__4_ ( .ip(n4884), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[44]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_1__4_ ( .ip(n4883), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[52]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_0__4_ ( .ip(n4882), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[60]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg_reg_5_ ( .ip(n4924), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[5]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_7__5_ ( .ip(n4881), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[5]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_6__5_ ( .ip(n4880), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[13]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_5__5_ ( .ip(n4879), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[21]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_4__5_ ( .ip(n4878), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[29]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_3__5_ ( .ip(n4877), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[37]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_2__5_ ( .ip(n4876), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[45]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_1__5_ ( .ip(n4875), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[53]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_0__5_ ( .ip(n4874), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[61]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg_reg_6_ ( .ip(n4923), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[6]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_7__6_ ( .ip(n4873), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[6]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_6__6_ ( .ip(n4872), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[14]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_5__6_ ( .ip(n4871), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[22]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_4__6_ ( .ip(n4870), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[30]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_3__6_ ( .ip(n4869), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[38]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_2__6_ ( .ip(n4868), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[46]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_1__6_ ( .ip(n4867), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[54]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_0__6_ ( .ip(n4866), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[62]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg_reg_7_ ( .ip(n4922), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[7]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_7__7_ ( .ip(n4865), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[7]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_6__7_ ( .ip(n4864), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[15]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_5__7_ ( .ip(n4863), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[23]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_4__7_ ( .ip(n4862), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[31]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_3__7_ ( .ip(n4861), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[39]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_2__7_ ( .ip(n4860), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[47]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_1__7_ ( .ip(n4859), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[55]) );
  drp_1 i_i2c_U_dff_rx_mem_reg_0__7_ ( .ip(n4858), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_i2c_U_dff_rx_mem[63]) );
  drp_1 i_apb_U_DW_apb_ahbsif_psel_en_reg ( .ip(n4205), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_psel_en) );
  drp_1 i_apb_U_DW_apb_ahbsif_penable_reg ( .ip(n4204), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_apb_penable) );
  drp_1 i_ssi_U_mstfsm_ctrl_cnt_reg_0_ ( .ip(n4203), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_ctrl_cnt[0]) );
  drp_1 i_ssi_U_mstfsm_ctrl_cnt_reg_1_ ( .ip(n4202), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_ctrl_cnt[1]) );
  drp_1 i_ssi_U_mstfsm_ctrl_cnt_reg_2_ ( .ip(n4201), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_ctrl_cnt[2]) );
  drp_1 i_ssi_U_mstfsm_ctrl_cnt_reg_3_ ( .ip(n4200), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_ctrl_cnt[3]) );
  drp_1 i_ssi_U_mstfsm_bit_cnt_reg_0_ ( .ip(n4199), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_bit_cnt[0]) );
  drp_1 i_ssi_U_mstfsm_bit_cnt_reg_1_ ( .ip(n4198), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_bit_cnt[1]) );
  drp_1 i_ssi_U_mstfsm_bit_cnt_reg_2_ ( .ip(n4197), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_bit_cnt[2]) );
  drp_1 i_ssi_U_mstfsm_bit_cnt_reg_3_ ( .ip(n4196), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_bit_cnt[3]) );
  drp_1 i_ssi_U_mstfsm_bit_cnt_reg_4_ ( .ip(n4195), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_bit_cnt[4]) );
  drp_1 i_ssi_U_mstfsm_spi1_control_reg ( .ip(n4194), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_spi1_control) );
  drp_1 i_ssi_U_mstfsm_spi0_control_reg ( .ip(n4193), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_spi0_control) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_15_ ( .ip(n4191), .ck(i_ssi_ssi_clk), 
        .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[15]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_14_ ( .ip(n4190), .ck(i_ssi_ssi_clk), 
        .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[14]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_13_ ( .ip(n4189), .ck(i_ssi_ssi_clk), 
        .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[13]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_12_ ( .ip(n6036), .ck(i_ssi_ssi_clk), 
        .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[12]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_11_ ( .ip(n4187), .ck(i_ssi_ssi_clk), 
        .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[11]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_9_ ( .ip(n4185), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[9]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_8_ ( .ip(n4184), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[8]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_7_ ( .ip(n4183), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[7]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_6_ ( .ip(n4182), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[6]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_5_ ( .ip(n4181), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[5]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_4_ ( .ip(n4180), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[4]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_3_ ( .ip(n4179), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[3]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_2_ ( .ip(n4178), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[2]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_1_ ( .ip(n4177), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[1]) );
  drp_1 i_ssi_U_mstfsm_frame_cnt_reg_0_ ( .ip(n4176), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_mstfsm_frame_cnt[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_arb_lost_tog_reg ( .ip(n4175), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_abrt_source[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_chk_win_reg ( .ip(n4174), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_chk_win) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_tx_pop_tog_reg ( .ip(n4173), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_tx_pop_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_mst_tx_ack_int_reg ( .ip(n4172), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_mst_tx_ack_vld) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_s_det_tog_reg ( .ip(n4171), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_s_det_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_q_reg ( .ip(n4170), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_q) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr_reg_0_ ( .ip(n4169), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr_reg_1_ ( .ip(n4168), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr_reg_2_ ( .ip(n4167), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr_reg_3_ ( .ip(n4166), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_rx_gen_call_tog_reg ( .ip(n4165), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_gen_call_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_slv_arb_lost_reg ( .ip(n4164), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_slv_arb_lost) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_rx_push_tog_reg ( .ip(n4163), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_push_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_p_det_tog_reg ( .ip(n4162), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_p_det_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ack_det_reg ( .ip(n4161), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ack_det) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_bwen_reg ( .ip(n4160), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_mst_rx_bwen) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_hcnt_cmplt_int_reg ( .ip(n8331), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_hcnt_cmplt_int) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_0_ ( .ip(n4158), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_1_ ( .ip(n4157), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_2_ ( .ip(n4156), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_4_ ( .ip(n4154), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_5_ ( .ip(n4153), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_7_ ( .ip(n4151), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_8_ ( .ip(n4150), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[8]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_9_ ( .ip(n4149), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_10_ ( .ip(n4148), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_11_ ( .ip(n4147), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_12_ ( .ip(n4146), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_13_ ( .ip(n4145), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_scl_hcnt_en_int_reg ( .ip(n4142), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_scl_hcnt_en) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_data_scl_lcnt_en_reg ( .ip(n4141), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_data_scl_lcnt_en) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count_reg_0_ ( .ip(n4140), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count_reg_1_ ( .ip(n4139), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count_reg_2_ ( .ip(n4138), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count_reg_3_ ( .ip(n4137), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_toggle_set_tx_empty_en_tog_reg ( .ip(n4136), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_set_tx_empty_en_flg) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr_reg_0_ ( .ip(n4135), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr_reg_1_ ( .ip(n4134), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr_reg_2_ ( .ip(n4133), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr_reg_3_ ( .ip(n4132), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr_reg_4_ ( .ip(n4131), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr_reg_5_ ( .ip(n4130), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr_reg_6_ ( .ip(n4129), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr_reg_7_ ( .ip(n4128), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[7]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_mst_tx_bwen_reg ( .ip(n4127), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_mst_tx_bwen) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_push_data_reg_0_ ( .ip(n4126), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_push_data[0]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_push_data_reg_1_ ( .ip(n4125), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_push_data[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_push_data_reg_2_ ( .ip(n4124), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_push_data[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_push_data_reg_3_ ( .ip(n4123), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_push_data[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_push_data_reg_4_ ( .ip(n4122), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_push_data[4]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_push_data_reg_5_ ( .ip(n4121), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_push_data[5]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_push_data_reg_6_ ( .ip(n4120), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_push_data[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_shift_rx_push_data_reg_7_ ( .ip(n4119), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_rx_push_data[7]) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_empty_n_reg ( .ip(i_ssi_U_fifo_U_tx_fifo_N33), 
        .ck(PCLK_pclk), .q(i_ssi_U_fifo_U_tx_fifo_empty_n) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_rd_addr_int_reg_2_ ( .ip(
        i_ssi_U_fifo_U_tx_fifo_N46), .ck(PCLK_pclk), .q(i_ssi_tx_rd_addr[2])
         );
  dp_1 i_ssi_U_fifo_U_tx_fifo_word_count_reg_2_ ( .ip(n11852), .ck(PCLK_pclk), 
        .q(i_ssi_U_fifo_unconnected_tx_wrd_count[2]) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_almost_empty_n_reg ( .ip(
        i_ssi_U_fifo_U_tx_fifo_N34), .ck(PCLK_pclk), .q(
        i_ssi_U_fifo_U_tx_fifo_almost_empty_n) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_wr_addr_at_max_reg ( .ip(
        i_ssi_U_fifo_U_tx_fifo_N40), .ck(PCLK_pclk), .q(
        i_ssi_U_fifo_U_tx_fifo_wr_addr_at_max) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_wr_addr_int_reg_2_ ( .ip(
        i_ssi_U_fifo_U_tx_fifo_N43), .ck(PCLK_pclk), .q(i_ssi_tx_wr_addr[2])
         );
  dp_1 i_ssi_U_fifo_U_rx_fifo_almost_full_int_reg ( .ip(n11830), .ck(PCLK_pclk), .q(i_ssi_U_fifo_switch_almost_full) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_empty_n_reg ( .ip(i_ssi_U_fifo_U_rx_fifo_N33), 
        .ck(PCLK_pclk), .q(i_ssi_U_fifo_U_rx_fifo_empty_n) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_wr_addr_int_reg_2_ ( .ip(
        i_ssi_U_fifo_U_rx_fifo_N43), .ck(PCLK_pclk), .q(i_ssi_rx_wr_addr[2])
         );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_wr_addr_int_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N43), .ck(PCLK_pclk), .q(
        i_i2c_rx_wr_addr[2]) );
  drp_2 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_0_ ( .ip(n4403), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[0]) );
  drp_2 i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt_reg_5_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N87), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[5])
         );
  drsp_1 i_apb_U_DW_apb_ahbsif_hready_resp_reg ( .ip(n4817), .ck(HCLK_hclk), 
        .rb(1'b1), .s(n11829), .q(i_apb_hready_resp) );
  drsp_1 i_ssi_U_regfile_sclk_active_reg ( .ip(n5235), .ck(PCLK_pclk), .rb(
        1'b1), .s(n11845), .q(i_ssi_sclk_active) );
  drsp_1 i_ssi_U_regfile_imr_ir_reg_3_ ( .ip(n4640), .ck(PCLK_pclk), .rb(1'b1), 
        .s(n11845), .q(i_ssi_imr[3]) );
  drsp_1 i_ssi_U_regfile_imr_ir_reg_1_ ( .ip(n4642), .ck(PCLK_pclk), .rb(1'b1), 
        .s(n11845), .q(i_ssi_imr[1]) );
  drsp_1 i_ssi_U_regfile_imr_ir_reg_4_ ( .ip(n4639), .ck(PCLK_pclk), .rb(1'b1), 
        .s(n11845), .q(i_ssi_imr[4]) );
  drsp_1 i_ssi_U_regfile_imr_ir_reg_0_ ( .ip(n4643), .ck(PCLK_pclk), .rb(1'b1), 
        .s(n11845), .q(i_ssi_imr[0]) );
  drsp_1 i_ssi_U_regfile_imr_ir_reg_2_ ( .ip(n4641), .ck(PCLK_pclk), .rb(1'b1), 
        .s(n11845), .q(i_ssi_imr[2]) );
  drsp_1 i_ssi_U_regfile_imr_ir_reg_5_ ( .ip(n4638), .ck(PCLK_pclk), .rb(1'b1), 
        .s(n11845), .q(i_ssi_imr[5]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_rd_addr_int_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N44), .ck(PCLK_pclk), .q(
        i_i2c_tx_rd_addr[0]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_rd_addr_int_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N46), .ck(PCLK_pclk), .q(
        i_i2c_tx_rd_addr[2]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_rd_addr_int_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N45), .ck(PCLK_pclk), .q(
        i_i2c_tx_rd_addr[1]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_rd_addr_at_max_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N39), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_rd_addr_at_max) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_error_int_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N38), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_tx_error_ir) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_full_int_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N37), .ck(PCLK_pclk), .q(
        i_i2c_tx_full) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_wr_addr_int_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N41), .ck(PCLK_pclk), .q(
        i_i2c_tx_wr_addr[0]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_wr_addr_at_max_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N40), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_wr_addr_at_max) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_wr_addr_int_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N42), .ck(PCLK_pclk), .q(
        i_i2c_tx_wr_addr[1]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_word_count_reg_2_ ( .ip(n11866), .ck(
        PCLK_pclk), .q(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[2]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_word_count_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N48), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[1]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_wr_addr_int_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N43), .ck(PCLK_pclk), .q(
        i_i2c_tx_wr_addr[2]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_word_count_reg_0_ ( .ip(n11867), .ck(
        PCLK_pclk), .q(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[0]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_empty_n_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N33), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_empty_n) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_almost_empty_n_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N34), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_almost_empty_n) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_full_int_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N37), .ck(PCLK_pclk), .q(
        i_i2c_rx_full) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_error_int_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N38), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_rx_error_ir) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_rd_addr_int_reg_2_ ( .ip(
        i_ssi_U_fifo_U_rx_fifo_N46), .ck(PCLK_pclk), .q(i_ssi_rx_rd_addr[2])
         );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_rd_addr_int_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N44), .ck(PCLK_pclk), .q(
        i_i2c_rx_rd_addr[0]) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_rd_addr_int_reg_1_ ( .ip(
        i_ssi_U_fifo_U_rx_fifo_N45), .ck(PCLK_pclk), .q(i_ssi_rx_rd_addr[1])
         );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_wr_addr_int_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N41), .ck(PCLK_pclk), .q(
        i_i2c_rx_wr_addr[0]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_rd_addr_int_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N45), .ck(PCLK_pclk), .q(
        i_i2c_rx_rd_addr[1]) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_rd_addr_int_reg_0_ ( .ip(n11849), .ck(PCLK_pclk), 
        .q(i_ssi_rx_rd_addr[0]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_wr_addr_int_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N42), .ck(PCLK_pclk), .q(
        i_i2c_rx_wr_addr[1]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_rd_addr_int_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N46), .ck(PCLK_pclk), .q(
        i_i2c_rx_rd_addr[2]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_wr_addr_at_max_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N40), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_wr_addr_at_max) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_rd_addr_at_max_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N39), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_rd_addr_at_max) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_rd_addr_at_max_reg ( .ip(
        i_ssi_U_fifo_U_rx_fifo_N39), .ck(PCLK_pclk), .q(
        i_ssi_U_fifo_U_rx_fifo_rd_addr_at_max) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_word_count_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N47), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[0]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_word_count_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N48), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[1]) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_error_int_reg ( .ip(i_ssi_U_fifo_U_rx_fifo_N38), 
        .ck(PCLK_pclk), .q(i_ssi_U_fifo_rx_error_ir) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_word_count_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N49), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[2]) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_error_int_reg ( .ip(i_ssi_U_fifo_U_tx_fifo_N38), 
        .ck(PCLK_pclk), .q(i_ssi_U_fifo_tx_error_ir) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_full_int_reg ( .ip(n11871), .ck(PCLK_pclk), .q(
        i_ssi_rx_full) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_almost_full_int_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N36), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_i_rx_almost_full) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_rd_addr_int_reg_0_ ( .ip(n11847), .ck(PCLK_pclk), 
        .q(i_ssi_tx_rd_addr[0]) );
  dp_1 i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_empty_n_reg ( .ip(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N33), .ck(PCLK_pclk), .q(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_empty_n) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_word_count_reg_0_ ( .ip(n11869), .ck(PCLK_pclk), 
        .q(i_ssi_U_fifo_unconnected_rx_wrd_count[0]) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_rd_addr_at_max_reg ( .ip(
        i_ssi_U_fifo_U_tx_fifo_N39), .ck(PCLK_pclk), .q(
        i_ssi_U_fifo_U_tx_fifo_rd_addr_at_max) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_wr_addr_int_reg_0_ ( .ip(n11846), .ck(PCLK_pclk), 
        .q(i_ssi_rx_wr_addr[0]) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_word_count_reg_1_ ( .ip(n11870), .ck(PCLK_pclk), 
        .q(i_ssi_U_fifo_unconnected_rx_wrd_count[1]) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_full_int_reg ( .ip(n11873), .ck(PCLK_pclk), .q(
        i_ssi_tx_full) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_rd_addr_int_reg_1_ ( .ip(
        i_ssi_U_fifo_U_tx_fifo_N45), .ck(PCLK_pclk), .q(i_ssi_tx_rd_addr[1])
         );
  dp_1 i_ssi_U_fifo_U_rx_fifo_wr_addr_at_max_reg ( .ip(
        i_ssi_U_fifo_U_rx_fifo_N40), .ck(PCLK_pclk), .q(
        i_ssi_U_fifo_U_rx_fifo_wr_addr_at_max) );
  dp_1 i_ssi_U_fifo_U_rx_fifo_wr_addr_int_reg_1_ ( .ip(
        i_ssi_U_fifo_U_rx_fifo_N42), .ck(PCLK_pclk), .q(i_ssi_rx_wr_addr[1])
         );
  dp_1 i_ssi_U_fifo_U_rx_fifo_word_count_reg_2_ ( .ip(n11850), .ck(PCLK_pclk), 
        .q(i_ssi_U_fifo_unconnected_rx_wrd_count[2]) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_wr_addr_int_reg_1_ ( .ip(
        i_ssi_U_fifo_U_tx_fifo_N42), .ck(PCLK_pclk), .q(i_ssi_tx_wr_addr[1])
         );
  dp_1 i_ssi_U_fifo_U_tx_fifo_wr_addr_int_reg_0_ ( .ip(n11848), .ck(PCLK_pclk), 
        .q(i_ssi_tx_wr_addr[0]) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_word_count_reg_0_ ( .ip(n11853), .ck(PCLK_pclk), 
        .q(i_ssi_U_fifo_unconnected_tx_wrd_count[0]) );
  dp_1 i_ssi_U_fifo_U_tx_fifo_word_count_reg_1_ ( .ip(n11872), .ck(PCLK_pclk), 
        .q(i_ssi_U_fifo_unconnected_tx_wrd_count[1]) );
  drsp_1 i_ssi_U_regfile_ctrlr0_ir_reg_0_ ( .ip(n4581), .ck(PCLK_pclk), .rb(
        1'b1), .s(n11845), .q(i_ssi_dfs[0]) );
  drp_2 i_ssi_U_regfile_baudr_reg_7_ ( .ip(n4620), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[7]) );
  drp_2 i_ssi_U_shift_ss_n_reg_0_ ( .ip(n11838), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(n11816) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda_r_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda), .ck(i_i2c_ic_clk), .rb(1'b1), .s(n11843), .q(i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda_r) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_start_sda_reg ( .ip(n4956), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11843), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_start_sda) );
  drsp_1 i_i2c_U_DW_apb_i2c_sync_tx_empty_sync_r_reg ( .ip(n11861), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11843), .q(
        i_i2c_U_DW_apb_i2c_sync_tx_empty_sync_r) );
  drsp_1 i_i2c_U_DW_apb_i2c_clk_gen_count_en_reg ( .ip(n4118), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11843), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_count_en) );
  drsp_1 i_i2c_U_DW_apb_i2c_rx_filter_scl_int_q_reg ( .ip(n6352), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11842), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_scl_int_q) );
  drsp_1 i_i2c_U_DW_apb_i2c_rx_filter_sda_data_int_reg ( .ip(n5129), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11842), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_sda_data_int) );
  drsp_1 i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt_reg_1_ ( .ip(n5088), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11843), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt[1]) );
  drsp_1 i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt_reg_0_ ( .ip(n5087), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11843), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt[0]) );
  drsp_1 i_i2c_U_DW_apb_i2c_rx_filter_sda_int_q_reg ( .ip(n11833), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11842), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_sda_int_q) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_stop_sda_reg ( .ip(n5042), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11843), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_stop_sda) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_stop_scl_reg ( .ip(n5043), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11842), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_stop_scl) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda_reg ( .ip(n4953), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11843), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl_reg ( .ip(n4954), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11843), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_slv_data_sda_reg ( .ip(n5103), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11842), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_data_sda) );
  drsp_1 i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_data_scl_reg ( .ip(n4930), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11842), .q(i_i2c_mst_rx_data_scl) );
  drsp_1 i_i2c_U_DW_apb_i2c_rx_filter_sda_post_hold_done_reg ( .ip(n5097), 
        .ck(i_i2c_ic_clk), .rb(1'b1), .s(n11842), .q(
        i_i2c_U_DW_apb_i2c_rx_filter_sda_post_hold_done) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_data_scl_reg ( .ip(n4117), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11842), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_data_scl) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_data_sda_reg ( .ip(n4116), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11842), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_data_sda) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_stop_sda_gate_r_reg ( .ip(
        i_i2c_U_DW_apb_i2c_tx_shift_N281), .ck(i_i2c_ic_clk), .rb(1'b1), .s(
        n11843), .q(i_i2c_U_DW_apb_i2c_tx_shift_stop_sda_gate_r) );
  drsp_1 i_i2c_U_DW_apb_i2c_tx_shift_data_sda_prev_r_reg ( .ip(n4934), .ck(
        i_i2c_ic_clk), .rb(1'b1), .s(n11843), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_data_sda_prev_r) );
  drp_2 i_ssi_U_mstfsm_ssi_oe_n_reg ( .ip(n11794), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(n11795) );
  dtrsp_2 i_ssi_U_mstfsm_frame_cnt_reg_10_ ( .ip(n5607), .sip(1'b0), .sm(
        n11836), .ck(i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .s(1'b0), .q(
        i_ssi_U_mstfsm_frame_cnt[10]) );
  drp_2 i_ssi_U_mstfsm_fsm_multi_mst_reg ( .ip(n4241), .ck(i_ssi_ssi_clk), 
        .rb(i_ssi_ssi_rst_n), .q(i_ssi_fsm_multi_mst) );
  drp_2 i_ssi_U_sclkgen_sclk_out_reg ( .ip(n4242), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_sclk_out) );
  dtrsp_2 i_ssi_U_mstfsm_frame_cnt_reg_16_ ( .ip(n5603), .sip(1'b0), .sm(
        n11836), .ck(i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .s(1'b0), .q(
        i_ssi_U_mstfsm_frame_cnt[16]) );
  drp_2 i_ssi_U_sclkgen_ssi_cnt_reg_0_ ( .ip(n11855), .ck(i_ssi_ssi_clk), .rb(
        i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[0]) );
  drp_2 i_ssi_U_sclkgen_ssi_cnt_reg_3_ ( .ip(i_ssi_U_sclkgen_N43), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[3])
         );
  drp_2 i_ssi_U_sclkgen_ssi_cnt_reg_4_ ( .ip(i_ssi_U_sclkgen_N44), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[4])
         );
  drp_2 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_5_ ( .ip(n4945), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[5]) );
  drp_2 i_ssi_U_regfile_baudr_reg_2_ ( .ip(n4625), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[2]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_9_ ( .ip(n4941), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[9]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr_reg_10_ ( .ip(n5152), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N84), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[2])
         );
  drp_1 i_i2c_U_DW_apb_i2c_mstfsm_mst_current_state_reg_1_ ( .ip(
        i_i2c_U_DW_apb_i2c_mstfsm_N73), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_mst_debug_cstate[1]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr_reg_9_ ( .ip(n5137), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[9]) );
  drp_1 i_ssi_U_shift_U_rx_shifter_rx_buffer_reg_15_ ( .ip(n4423), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_rx_push_data[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_14_ ( .ip(n4144), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_12_ ( .ip(n4938), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_15_ ( .ip(n4935), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_13_ ( .ip(n4937), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[13]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_10_ ( .ip(n4940), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[10]) );
  drp_1 i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r_reg_11_ ( .ip(n4939), 
        .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[11]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_6_ ( .ip(n5121), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_14_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N76), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[14]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_3_ ( .ip(n4155), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr_reg_12_ ( .ip(
        i_i2c_U_DW_apb_i2c_clk_gen_N74), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[12]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_6_ ( .ip(n4152), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[6]) );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr_reg_15_ ( .ip(n4143), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[15]) );
  drp_1 i_i2c_U_DW_apb_i2c_sync_U_ic_ss_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_ss_sync_next_sample_syncm1_0_), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(i_i2c_ic_ss_sync) );
  drp_4 i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r_reg ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_hs), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r) );
  drp_2 i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt_reg_4_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N86), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[4])
         );
  drp_4 i_ahb_U_mux_hsel_prev_reg_4_ ( .ip(n4852), .ck(HCLK_hclk), .rb(
        HRESETn_hresetn), .q(i_ahb_U_mux_hsel_prev[4]) );
  drp_2 i_ssi_U_sclkgen_sclk_re_ir_reg ( .ip(i_ssi_U_sclkgen_N74), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_sclk_re) );
  drp_2 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_9_ ( .ip(n4394), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[9]) );
  drp_2 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_5_ ( .ip(n4398), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[5]) );
  drp_2 i_i2c_U_DW_apb_i2c_mstfsm_mst_current_state_reg_2_ ( .ip(
        i_i2c_U_DW_apb_i2c_mstfsm_N74), .ck(i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), 
        .q(i_i2c_mst_debug_cstate[2]) );
  drp_2 i_i2c_U_DW_apb_i2c_sync_U_ic_hs_sync_sample_syncl_reg_0_ ( .ip(
        i_i2c_U_DW_apb_i2c_sync_U_ic_hs_sync_next_sample_syncm1_0_), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv) );
  drp_2 i_ssi_U_regfile_ctrlr1_reg_9_ ( .ip(n4610), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[9]) );
  drp_1 i_ssi_U_regfile_start_xfer_reg ( .ip(i_ssi_U_regfile_N452), .ck(
        PCLK_pclk), .rb(PRESETn_presetn), .q(i_ssi_start_xfer) );
  drp_2 i_ssi_U_shift_U_tx_shifter_txd_reg ( .ip(n4388), .ck(i_ssi_ssi_clk), 
        .rb(i_ssi_ssi_rst_n), .q(i_ssi_txd) );
  drp_1 i_ssi_U_regfile_baud2_reg ( .ip(n5234), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baud2) );
  drp_2 i_ssi_U_regfile_ctrlr1_reg_15_ ( .ip(n4604), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[15]) );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_11_ ( .ip(n4608), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[11]) );
  drp_2 i_ssi_U_regfile_ctrlr1_reg_8_ ( .ip(n4611), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[8]) );
  drp_4 i_ssi_U_sclkgen_ssi_cnt_reg_2_ ( .ip(i_ssi_U_sclkgen_N42), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[2])
         );
  drp_1 i_ssi_U_regfile_ctrlr1_reg_3_ ( .ip(n4600), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[3]) );
  drp_2 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_15_ ( .ip(n4389), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[15]) );
  drp_2 i_ssi_U_sclkgen_ssi_cnt_reg_9_ ( .ip(i_ssi_U_sclkgen_N49), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[9])
         );
  drp_4 i_ssi_U_sclkgen_ssi_cnt_reg_1_ ( .ip(i_ssi_U_sclkgen_N41), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(i_ssi_U_sclkgen_ssi_cnt[1])
         );
  drp_2 i_ssi_U_regfile_ctrlr1_reg_10_ ( .ip(n4609), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[10]) );
  drp_2 i_ssi_U_regfile_ctrlr1_reg_6_ ( .ip(n4597), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[6]) );
  drsp_1 i_ssi_U_regfile_ctrlr0_ir_reg_2_ ( .ip(n4583), .ck(PCLK_pclk), .rb(
        1'b1), .s(n11845), .q(i_ssi_dfs[2]) );
  drsp_1 i_ssi_U_regfile_ctrlr0_ir_reg_1_ ( .ip(n4582), .ck(PCLK_pclk), .rb(
        1'b1), .s(n11845), .q(i_ssi_dfs[1]) );
  drp_2 i_ssi_U_regfile_baudr_reg_1_ ( .ip(n4626), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[1]) );
  drp_2 i_ssi_U_shift_U_tx_shifter_tx_shift_reg_reg_11_ ( .ip(n4392), .ck(
        i_ssi_ssi_clk), .rb(i_ssi_ssi_rst_n), .q(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[11]) );
  drp_2 i_ssi_U_regfile_ctrlr1_reg_7_ ( .ip(n4596), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_U_regfile_ctrlr1_int[7]) );
  drsp_1 i_ssi_U_regfile_ctrlr0_ir_reg_3_ ( .ip(n4584), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .s(1'b0), .q(i_ssi_dfs[3]) );
  drp_1 i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt_reg_6_ ( .ip(
        i_i2c_U_DW_apb_i2c_rx_filter_N88), .ck(i_i2c_ic_clk), .rb(
        i_i2c_ic_rst_n), .q(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[6])
         );
  drp_1 i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr_reg_0_ ( .ip(n5127), .ck(
        i_i2c_ic_clk), .rb(i_i2c_ic_rst_n), .q(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[0]) );
  drp_1 i_ssi_U_regfile_baudr_reg_3_ ( .ip(n4624), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[3]) );
  drp_2 i_ssi_U_regfile_baudr_reg_6_ ( .ip(n4621), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[6]) );
  drp_2 i_ssi_U_regfile_baudr_reg_5_ ( .ip(n4622), .ck(PCLK_pclk), .rb(
        PRESETn_presetn), .q(i_ssi_baudr[5]) );
  buf_2 U5559 ( .ip(n11121), .op(n11107) );
  inv_1 U5560 ( .ip(n10229), .op(n5286) );
  nor2_2 U5561 ( .ip1(n6861), .ip2(n6858), .op(n5249) );
  nor2_2 U5562 ( .ip1(n7176), .ip2(n7177), .op(n7201) );
  and3_1 U5563 ( .ip1(n10239), .ip2(i_ssi_tx_rd_addr[2]), .ip3(n10233), .op(
        n10402) );
  and2_1 U5564 ( .ip1(n10240), .ip2(i_ssi_tx_rd_addr[1]), .op(n10400) );
  nor2_2 U5565 ( .ip1(i_ssi_tx_rd_addr[1]), .ip2(n10234), .op(n10389) );
  nand2_2 U5566 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[0]), .ip2(
        n8730), .op(n8688) );
  nor2_2 U5567 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(n6510), .op(n11153) );
  nand2_1 U5568 ( .ip1(n7073), .ip2(n7069), .op(n7070) );
  mux2_1 U5569 ( .ip1(i_i2c_ic_fs_hcnt[2]), .ip2(i_i2c_ic_hcnt[2]), .s(n6060), 
        .op(n8223) );
  mux2_1 U5570 ( .ip1(i_i2c_ic_fs_lcnt[2]), .ip2(i_i2c_ic_lcnt[2]), .s(n6060), 
        .op(n7116) );
  mux2_4 U5571 ( .ip1(i_apb_pwdata_int[5]), .ip2(i_ssi_baudr[5]), .s(n9746), 
        .op(n4622) );
  mux2_4 U5572 ( .ip1(i_apb_pwdata_int[6]), .ip2(i_ssi_baudr[6]), .s(n9746), 
        .op(n4621) );
  nor2_1 U5573 ( .ip1(n9161), .ip2(n9124), .op(n9123) );
  nand2_1 U5574 ( .ip1(n6066), .ip2(n6065), .op(n5464) );
  nand2_1 U5575 ( .ip1(i_i2c_ic_hcnt[1]), .ip2(n6041), .op(n6065) );
  mux2_2 U5576 ( .ip1(n5456), .ip2(n5457), .s(n6060), .op(n5455) );
  inv_1 U5577 ( .ip(n6160), .op(n6190) );
  nand2_1 U5578 ( .ip1(n6073), .ip2(n6072), .op(n6160) );
  mux2_2 U5579 ( .ip1(i_i2c_ic_fs_hcnt[5]), .ip2(i_i2c_ic_hcnt[5]), .s(n6060), 
        .op(n8211) );
  nor2_1 U5580 ( .ip1(n9189), .ip2(n9188), .op(n9246) );
  inv_1 U5581 ( .ip(n5427), .op(n5270) );
  mux2_2 U5582 ( .ip1(i_i2c_ic_fs_hcnt[4]), .ip2(i_i2c_ic_hcnt[4]), .s(n6060), 
        .op(n8215) );
  nor2_1 U5583 ( .ip1(n9163), .ip2(n9162), .op(n9172) );
  nor2_1 U5584 ( .ip1(n7072), .ip2(n7021), .op(n7063) );
  nor3_1 U5585 ( .ip1(n8240), .ip2(n8239), .ip3(n8238), .op(n8216) );
  nor2_1 U5586 ( .ip1(n9233), .ip2(n9234), .op(n9238) );
  nand2_1 U5587 ( .ip1(n5261), .ip2(n8166), .op(n8208) );
  buf_1 U5588 ( .ip(n6041), .op(n5458) );
  inv_1 U5589 ( .ip(n8571), .op(n5266) );
  inv_1 U5590 ( .ip(n8536), .op(n5268) );
  or2_1 U5591 ( .ip1(n8271), .ip2(n8270), .op(n5465) );
  inv_1 U5592 ( .ip(n8208), .op(n5267) );
  inv_1 U5593 ( .ip(n5567), .op(n9282) );
  inv_1 U5594 ( .ip(n8530), .op(n5277) );
  or2_1 U5595 ( .ip1(n9201), .ip2(n9282), .op(n5579) );
  nor3_1 U5596 ( .ip1(n5916), .ip2(n6476), .ip3(n5917), .op(n5946) );
  nand2_1 U5597 ( .ip1(n9212), .ip2(n9211), .op(n5567) );
  nor2_1 U5598 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[9]), .ip2(n5532), .op(n5971) );
  nor4_1 U5599 ( .ip1(n10919), .ip2(n7834), .ip3(n10930), .ip4(n7833), .op(
        n7836) );
  buf_1 U5600 ( .ip(i_i2c_ic_ss_sync), .op(n5907) );
  inv_1 U5601 ( .ip(i_ssi_baudr[3]), .op(n6432) );
  nor2_1 U5602 ( .ip1(n9607), .ip2(i_apb_U_DW_apb_ahbsif_nextstate[0]), .op(
        n7406) );
  inv_1 U5603 ( .ip(i_i2c_mst_debug_cstate[2]), .op(n6351) );
  nand2_1 U5604 ( .ip1(n11854), .ip2(n6309), .op(n10199) );
  inv_1 U5605 ( .ip(n5613), .op(n5617) );
  nor2_1 U5606 ( .ip1(n10713), .ip2(n10712), .op(n10720) );
  inv_1 U5607 ( .ip(n5476), .op(n8327) );
  nand2_1 U5608 ( .ip1(n9449), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[5]), .op(n9452) );
  nand4_1 U5609 ( .ip1(n8117), .ip2(n8116), .ip3(n8115), .ip4(n11093), .op(
        n8118) );
  inv_1 U5610 ( .ip(n7721), .op(n7699) );
  inv_2 U5611 ( .ip(n10453), .op(n5271) );
  inv_1 U5612 ( .ip(n5613), .op(n5616) );
  nand2_1 U5613 ( .ip1(i_apb_U_DW_apb_ahbsif_nextstate[0]), .ip2(n10087), .op(
        n10095) );
  nor3_1 U5614 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(i_ahb_U_mux_hsel_prev[3]), .ip3(n6516), .op(n6676) );
  inv_1 U5615 ( .ip(n11837), .op(n10713) );
  nand4_1 U5616 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[0]), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[1]), .ip3(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[2]), .ip4(n11182), .op(n11135)
         );
  xor2_1 U5617 ( .ip1(n8317), .ip2(n8316), .op(n8318) );
  buf_1 U5618 ( .ip(n11401), .op(n11839) );
  nor3_1 U5619 ( .ip1(i_apb_paddr[12]), .ip2(n11152), .ip3(n6025), .op(n11401)
         );
  nor2_1 U5620 ( .ip1(n9432), .ip2(n9452), .op(n9454) );
  xor2_1 U5621 ( .ip1(n7754), .ip2(n7753), .op(n7755) );
  nand3_1 U5622 ( .ip1(n7566), .ip2(n7587), .ip3(n7565), .op(n7585) );
  nor4_1 U5623 ( .ip1(i_i2c_tx_wr_addr[2]), .ip2(i_i2c_tx_wr_addr[1]), .ip3(
        i_i2c_tx_wr_addr[0]), .ip4(n11325), .op(n11333) );
  and2_1 U5624 ( .ip1(n10705), .ip2(n10802), .op(n10865) );
  and2_1 U5625 ( .ip1(n5616), .ip2(n6686), .op(n6687) );
  nor2_1 U5626 ( .ip1(n9683), .ip2(n10095), .op(n11121) );
  nor2_1 U5627 ( .ip1(n6848), .ip2(n6847), .op(n10084) );
  nor2_1 U5628 ( .ip1(n6827), .ip2(n11158), .op(n11162) );
  nor2_1 U5629 ( .ip1(n9335), .ip2(n8315), .op(n4151) );
  nor2_1 U5630 ( .ip1(n7774), .ip2(n7741), .op(n5124) );
  nor2_1 U5631 ( .ip1(n7667), .ip2(n7661), .op(n5092) );
  xor2_1 U5632 ( .ip1(i_ssi_U_fifo_tx_pop_edge), .ip2(i_ssi_tx_pop), .op(
        i_ssi_tx_pop_sync) );
  or2_1 U5633 ( .ip1(n11348), .ip2(n6683), .op(ex_i_ahb_AHB_Slave_PID_hready)
         );
  inv_1 U5634 ( .ip(n9662), .op(ex_i_ahb_AHB_MASTER_CORTEXM0_hready) );
  xor2_1 U5635 ( .ip1(n7121), .ip2(n7122), .op(n5245) );
  and2_1 U5636 ( .ip1(n5914), .ip2(n5530), .op(n5246) );
  and2_2 U5637 ( .ip1(n5813), .ip2(n5812), .op(n5247) );
  ab_or_c_or_d U5638 ( .ip1(n7881), .ip2(n8111), .ip3(n7880), .ip4(n7879), 
        .op(n5248) );
  ab_or_c_or_d U5639 ( .ip1(i_ssi_U_mstfsm_c_state[1]), .ip2(
        i_ssi_U_mstfsm_abort_ir), .ip3(n10421), .ip4(n10422), .op(n5250) );
  or2_1 U5640 ( .ip1(n5621), .ip2(n5626), .op(n5251) );
  nor2_2 U5641 ( .ip1(i_ssi_tx_rd_addr[2]), .ip2(n10244), .op(n5252) );
  nand2_2 U5642 ( .ip1(n10226), .ip2(n10223), .op(n5253) );
  nand2_2 U5643 ( .ip1(n10226), .ip2(n10227), .op(n5254) );
  nand2_2 U5644 ( .ip1(n10226), .ip2(n10222), .op(n5255) );
  nand2_2 U5645 ( .ip1(n10226), .ip2(n10225), .op(n5256) );
  and2_1 U5646 ( .ip1(n5586), .ip2(n5587), .op(n5257) );
  and2_1 U5647 ( .ip1(n9247), .ip2(n9250), .op(n5258) );
  nand2_1 U5648 ( .ip1(n5257), .ip2(n9193), .op(n9212) );
  xnor2_2 U5649 ( .ip1(n7073), .ip2(n7072), .op(n5259) );
  and2_1 U5650 ( .ip1(n6057), .ip2(n6056), .op(n5260) );
  and2_1 U5651 ( .ip1(n8167), .ip2(n8217), .op(n5261) );
  inv_1 U5652 ( .ip(n8764), .op(n5265) );
  xor2_1 U5653 ( .ip1(n8692), .ip2(n8693), .op(n5262) );
  xor2_1 U5654 ( .ip1(n8923), .ip2(n8924), .op(n5263) );
  xor2_1 U5655 ( .ip1(n6132), .ip2(n6131), .op(n5264) );
  nand2_2 U5656 ( .ip1(n9972), .ip2(n5748), .op(n10703) );
  nand2_2 U5657 ( .ip1(n5505), .ip2(n5504), .op(n5329) );
  inv_1 U5658 ( .ip(n10440), .op(n10415) );
  nand2_2 U5659 ( .ip1(n5360), .ip2(n5357), .op(n5514) );
  nor2_4 U5660 ( .ip1(n5360), .ip2(n5281), .op(n10672) );
  nand2_2 U5661 ( .ip1(n10439), .ip2(n10479), .op(n10488) );
  inv_4 U5662 ( .ip(n9913), .op(n10479) );
  nand2_2 U5663 ( .ip1(n10981), .ip2(n10980), .op(n10990) );
  nand2_4 U5664 ( .ip1(n10987), .ip2(n10979), .op(n10980) );
  mux2_2 U5665 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[8]), .ip2(n10483), .s(n10516), .op(n4395) );
  nand2_1 U5666 ( .ip1(n10516), .ip2(n5298), .op(n5297) );
  inv_2 U5667 ( .ip(n5446), .op(n5450) );
  nand2_1 U5668 ( .ip1(n5281), .ip2(n5360), .op(n5310) );
  or2_2 U5669 ( .ip1(n5360), .ip2(n5357), .op(n5424) );
  nand2_2 U5670 ( .ip1(n10681), .ip2(n10662), .op(n10663) );
  xor2_1 U5671 ( .ip1(i_ssi_U_mstfsm_frame_cnt[15]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[15]), .op(n5645) );
  nand2_4 U5672 ( .ip1(n10442), .ip2(n10743), .op(n5410) );
  nor2_2 U5673 ( .ip1(n9469), .ip2(n5601), .op(n4938) );
  nor2_2 U5674 ( .ip1(n9331), .ip2(n8686), .op(n5161) );
  nor2_2 U5675 ( .ip1(n7729), .ip2(n7726), .op(i_i2c_U_DW_apb_i2c_clk_gen_N71)
         );
  and2_1 U5676 ( .ip1(n9405), .ip2(n9349), .op(n9350) );
  xnor2_1 U5677 ( .ip1(n5583), .ip2(n5584), .op(n5582) );
  nor2_1 U5678 ( .ip1(n8754), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[15]), .op(n8612) );
  and3_1 U5679 ( .ip1(n5558), .ip2(n5551), .ip3(n5560), .op(n5429) );
  nor2_1 U5680 ( .ip1(n6099), .ip2(n6098), .op(n6100) );
  xnor2_1 U5681 ( .ip1(n6943), .ip2(n6942), .op(n8754) );
  nor2_1 U5682 ( .ip1(n8216), .ip2(n5595), .op(n8242) );
  nor2_1 U5683 ( .ip1(n8268), .ip2(n5465), .op(n5460) );
  nor2_1 U5684 ( .ip1(n6117), .ip2(n6116), .op(n6119) );
  nor2_1 U5685 ( .ip1(n6102), .ip2(n6095), .op(n6099) );
  or2_1 U5686 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[9]), .ip2(n5474), 
        .op(n5551) );
  and2_1 U5687 ( .ip1(n5470), .ip2(n8187), .op(n8268) );
  and3_1 U5688 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[8]), .ip2(n5554), .ip3(n5475), .op(n5552) );
  xnor2_1 U5689 ( .ip1(n8186), .ip2(n8185), .op(n8187) );
  nor2_1 U5690 ( .ip1(n6075), .ip2(n6190), .op(n6182) );
  inv_1 U5691 ( .ip(n6990), .op(n5274) );
  and2_1 U5692 ( .ip1(n5545), .ip2(n8214), .op(n8238) );
  nand2_1 U5693 ( .ip1(n6160), .ip2(n6078), .op(n6086) );
  nor2_1 U5694 ( .ip1(n8188), .ip2(n8189), .op(n8184) );
  inv_2 U5695 ( .ip(n8548), .op(n5269) );
  nand2_1 U5696 ( .ip1(n8168), .ip2(n8260), .op(n8189) );
  xnor2_1 U5697 ( .ip1(n7115), .ip2(n7114), .op(n8442) );
  inv_1 U5698 ( .ip(n8443), .op(n5280) );
  and2_1 U5699 ( .ip1(n8165), .ip2(n8247), .op(n8166) );
  nor2_1 U5700 ( .ip1(n7121), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[0]), .op(n8889) );
  nor2_1 U5701 ( .ip1(n8207), .ip2(n8258), .op(n8260) );
  nor2_1 U5702 ( .ip1(n7121), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[0]), .op(n8586) );
  nand2_1 U5703 ( .ip1(n7025), .ip2(n7113), .op(n7090) );
  mux2_1 U5704 ( .ip1(i_i2c_ic_fs_hcnt[10]), .ip2(i_i2c_ic_hcnt[10]), .s(n5458), .op(n8262) );
  buf_4 U5705 ( .ip(n6857), .op(n11117) );
  nand2_4 U5706 ( .ip1(n8219), .ip2(n6061), .op(n6062) );
  nand4_2 U5707 ( .ip1(n11833), .ip2(n6352), .ip3(i_i2c_ic_enable_sync), .ip4(
        n9583), .op(n7729) );
  nor2_2 U5708 ( .ip1(n7667), .ip2(n7658), .op(n5093) );
  inv_1 U5709 ( .ip(n5461), .op(n5282) );
  inv_1 U5710 ( .ip(n7021), .op(n7071) );
  nor2_1 U5711 ( .ip1(n8223), .ip2(n8219), .op(n8167) );
  inv_1 U5712 ( .ip(n7121), .op(n7123) );
  nor2_1 U5713 ( .ip1(n7122), .ip2(n7121), .op(n7113) );
  inv_2 U5714 ( .ip(n5455), .op(n8219) );
  nor2_2 U5715 ( .ip1(n8215), .ip2(n6074), .op(n6075) );
  mux2_1 U5716 ( .ip1(i_i2c_ic_fs_hcnt[2]), .ip2(i_i2c_ic_hcnt[2]), .s(n6270), 
        .op(n5469) );
  mux2_1 U5717 ( .ip1(n5463), .ip2(n5462), .s(n6043), .op(n5461) );
  nor2_2 U5718 ( .ip1(n8215), .ip2(n8211), .op(n8247) );
  mux2_1 U5719 ( .ip1(i_i2c_ic_fs_lcnt[1]), .ip2(i_i2c_ic_lcnt[1]), .s(n6270), 
        .op(n7122) );
  mux2_1 U5720 ( .ip1(i_i2c_ic_fs_hcnt[2]), .ip2(i_i2c_ic_hcnt[2]), .s(n6041), 
        .op(n5468) );
  mux2_1 U5721 ( .ip1(i_i2c_ic_fs_lcnt[4]), .ip2(i_i2c_ic_lcnt[4]), .s(n6270), 
        .op(n7105) );
  mux2_1 U5722 ( .ip1(i_i2c_ic_fs_lcnt[5]), .ip2(i_i2c_ic_lcnt[5]), .s(n6270), 
        .op(n7026) );
  mux2_1 U5723 ( .ip1(i_i2c_ic_fs_lcnt[10]), .ip2(i_i2c_ic_lcnt[10]), .s(n6270), .op(n8550) );
  mux2_2 U5724 ( .ip1(i_i2c_ic_fs_lcnt[9]), .ip2(i_i2c_ic_lcnt[9]), .s(n6270), 
        .op(n7021) );
  mux2_1 U5725 ( .ip1(i_i2c_ic_fs_hcnt[9]), .ip2(i_i2c_ic_hcnt[9]), .s(n6270), 
        .op(n5454) );
  buf_2 U5726 ( .ip(n7266), .op(n7239) );
  mux2_1 U5727 ( .ip1(i_i2c_ic_fs_hcnt[9]), .ip2(i_i2c_ic_hcnt[9]), .s(n6270), 
        .op(n8207) );
  nor2_2 U5728 ( .ip1(n6853), .ip2(i_apb_U_DW_apb_ahbsif_nextstate[0]), .op(
        n10091) );
  nand2_1 U5729 ( .ip1(n5860), .ip2(n7644), .op(n5905) );
  nor2_2 U5730 ( .ip1(n10105), .ip2(n7415), .op(n9690) );
  or2_1 U5731 ( .ip1(n10203), .ip2(i_ssi_tx_wr_addr[2]), .op(n6337) );
  nand2_1 U5732 ( .ip1(n5473), .ip2(n5843), .op(n5857) );
  and2_1 U5733 ( .ip1(n10228), .ip2(n10227), .op(n10229) );
  nor2_2 U5734 ( .ip1(i_ssi_tx_wr_addr[0]), .ip2(n10199), .op(n10226) );
  and2_1 U5735 ( .ip1(i_ssi_U_mstfsm_tx_load_en_int), .ip2(n5308), .op(n5307)
         );
  nor2_2 U5736 ( .ip1(n9883), .ip2(n5638), .op(n9889) );
  inv_1 U5737 ( .ip(n5855), .op(n5856) );
  nor2_1 U5738 ( .ip1(n7378), .ip2(n5364), .op(n5482) );
  xor2_1 U5739 ( .ip1(n7644), .ip2(n7668), .op(n7645) );
  nand4_1 U5740 ( .ip1(n6635), .ip2(n6634), .ip3(n6633), .ip4(n6632), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[23]) );
  nand4_1 U5741 ( .ip1(n6520), .ip2(n6519), .ip3(n6518), .ip4(n6517), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[31]) );
  nand4_1 U5742 ( .ip1(n6650), .ip2(n6649), .ip3(n6648), .ip4(n6647), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[10]) );
  nand4_1 U5743 ( .ip1(n6625), .ip2(n6624), .ip3(n6623), .ip4(n6622), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[25]) );
  nand4_1 U5744 ( .ip1(n6615), .ip2(n6614), .ip3(n6613), .ip4(n6612), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[7]) );
  nor4_2 U5745 ( .ip1(i_i2c_tx_wr_addr[2]), .ip2(i_i2c_tx_wr_addr[0]), .ip3(
        n11323), .ip4(n11325), .op(n11331) );
  nand4_1 U5746 ( .ip1(n6620), .ip2(n6619), .ip3(n6618), .ip4(n6617), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[26]) );
  nand4_1 U5747 ( .ip1(n6525), .ip2(n6524), .ip3(n6523), .ip4(n6522), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[27]) );
  nor4_2 U5748 ( .ip1(i_i2c_tx_wr_addr[0]), .ip2(i_i2c_tx_wr_addr[1]), .ip3(
        n11321), .ip4(n11325), .op(n11329) );
  nand4_1 U5749 ( .ip1(n6560), .ip2(n6559), .ip3(n6558), .ip4(n6557), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[24]) );
  nand4_1 U5750 ( .ip1(n6575), .ip2(n6574), .ip3(n6573), .ip4(n6572), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[28]) );
  nand4_1 U5751 ( .ip1(n6540), .ip2(n6539), .ip3(n6538), .ip4(n6537), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[17]) );
  nand4_1 U5752 ( .ip1(n6670), .ip2(n6669), .ip3(n6668), .ip4(n6667), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[9]) );
  nand4_1 U5753 ( .ip1(n6545), .ip2(n6544), .ip3(n6543), .ip4(n6542), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[29]) );
  nand4_1 U5754 ( .ip1(n6600), .ip2(n6599), .ip3(n6598), .ip4(n6597), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[6]) );
  nand4_1 U5755 ( .ip1(n6660), .ip2(n6659), .ip3(n6658), .ip4(n6657), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[30]) );
  nand4_1 U5756 ( .ip1(n6590), .ip2(n6589), .ip3(n6588), .ip4(n6587), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[19]) );
  nand4_1 U5757 ( .ip1(n6535), .ip2(n6534), .ip3(n6533), .ip4(n6532), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[21]) );
  nand4_1 U5758 ( .ip1(n6565), .ip2(n6564), .ip3(n6563), .ip4(n6562), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[2]) );
  nand4_1 U5759 ( .ip1(n6605), .ip2(n6604), .ip3(n6603), .ip4(n6602), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[11]) );
  nand4_1 U5760 ( .ip1(n6585), .ip2(n6584), .ip3(n6583), .ip4(n6582), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[4]) );
  nand4_1 U5761 ( .ip1(n6640), .ip2(n6639), .ip3(n6638), .ip4(n6637), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[14]) );
  nand4_1 U5762 ( .ip1(n6645), .ip2(n6644), .ip3(n6643), .ip4(n6642), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[20]) );
  nand4_1 U5763 ( .ip1(n6570), .ip2(n6569), .ip3(n6568), .ip4(n6567), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[12]) );
  nand4_1 U5764 ( .ip1(n6610), .ip2(n6609), .ip3(n6608), .ip4(n6607), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[3]) );
  nand4_1 U5765 ( .ip1(n6675), .ip2(n6674), .ip3(n6673), .ip4(n6672), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[13]) );
  nand4_1 U5766 ( .ip1(n6550), .ip2(n6549), .ip3(n6548), .ip4(n6547), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[0]) );
  nand4_1 U5767 ( .ip1(n6530), .ip2(n6529), .ip3(n6528), .ip4(n6527), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[8]) );
  nand4_1 U5768 ( .ip1(n6655), .ip2(n6654), .ip3(n6653), .ip4(n6652), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[1]) );
  nand4_1 U5769 ( .ip1(n6555), .ip2(n6554), .ip3(n6553), .ip4(n6552), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[18]) );
  inv_2 U5770 ( .ip(n6688), .op(n6937) );
  nand4_1 U5771 ( .ip1(n6630), .ip2(n6629), .ip3(n6628), .ip4(n6627), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[16]) );
  nand4_1 U5772 ( .ip1(n6580), .ip2(n6579), .ip3(n6578), .ip4(n6577), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[22]) );
  nand4_1 U5773 ( .ip1(n6595), .ip2(n6594), .ip3(n6593), .ip4(n6592), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[5]) );
  nand4_1 U5774 ( .ip1(n6665), .ip2(n6664), .ip3(n6663), .ip4(n6662), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hrdata[15]) );
  inv_2 U5775 ( .ip(ex_i_ahb_AHB_Slave_PID_hready), .op(n9662) );
  and2_1 U5776 ( .ip1(n5949), .ip2(n5950), .op(n5555) );
  and2_1 U5777 ( .ip1(n5735), .ip2(n5736), .op(n5340) );
  or2_1 U5778 ( .ip1(n5798), .ip2(n5312), .op(n5715) );
  xor2_2 U5779 ( .ip1(n10996), .ip2(n6406), .op(n5515) );
  nand2_1 U5780 ( .ip1(n9123), .ip2(n9129), .op(n9132) );
  and3_1 U5781 ( .ip1(n5289), .ip2(n5426), .ip3(n5425), .op(n5354) );
  nand4_2 U5782 ( .ip1(n6682), .ip2(n6681), .ip3(n6680), .ip4(n6679), .op(
        n11348) );
  inv_1 U5783 ( .ip(n5730), .op(n5289) );
  nor2_2 U5784 ( .ip1(i_i2c_mst_debug_cstate[4]), .ip2(n7779), .op(n7873) );
  inv_1 U5785 ( .ip(n5510), .op(n5290) );
  inv_1 U5786 ( .ip(n5759), .op(n5303) );
  xnor2_2 U5787 ( .ip1(n6897), .ip2(i_ssi_rx_push), .op(n11837) );
  nand2_1 U5788 ( .ip1(n5760), .ip2(n5758), .op(n5302) );
  and2_1 U5789 ( .ip1(n5710), .ip2(i_ssi_U_mstfsm_frame_cnt[15]), .op(n5321)
         );
  mux2_1 U5790 ( .ip1(n9754), .ip2(n7349), .s(i_ssi_baudr[1]), .op(n7350) );
  xor2_1 U5791 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_sda_data_int), .ip2(n7590), 
        .op(n7565) );
  xor2_1 U5792 ( .ip1(n6419), .ip2(i_ssi_baudr[4]), .op(n6421) );
  inv_2 U5793 ( .ip(n10802), .op(n5291) );
  nor2_1 U5794 ( .ip1(i_ssi_tx_rd_addr[0]), .ip2(i_ssi_tx_rd_addr[2]), .op(
        n10240) );
  nor2_1 U5795 ( .ip1(i_ssi_baudr[2]), .ip2(i_ssi_baudr[3]), .op(n5356) );
  inv_1 U5796 ( .ip(i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv), .op(n5851) );
  and2_1 U5797 ( .ip1(i_i2c_mst_debug_cstate[1]), .ip2(
        i_i2c_mst_debug_cstate[2]), .op(n5846) );
  inv_1 U5798 ( .ip(i_ssi_cfs[0]), .op(n10437) );
  inv_1 U5799 ( .ip(i_ssi_U_mstfsm_last_frame), .op(n5336) );
  buf_1 U5800 ( .ip(i_ssi_U_regfile_ctrlr1_int[11]), .op(n5391) );
  inv_2 U5801 ( .ip(n10429), .op(n5272) );
  inv_1 U5802 ( .ip(i_ssi_cfs[2]), .op(n10441) );
  xnor2_1 U5803 ( .ip1(i_ssi_U_mstfsm_bit_cnt[2]), .ip2(i_ssi_dfs[2]), .op(
        n5759) );
  xor2_2 U5804 ( .ip1(n8960), .ip2(n8959), .op(n8961) );
  xor2_2 U5805 ( .ip1(n6249), .ip2(n7769), .op(n7770) );
  nor2_1 U5806 ( .ip1(n9469), .ip2(n5605), .op(n4939) );
  and2_1 U5807 ( .ip1(i_i2c_scl_s_setup_en), .ip2(n7159), .op(n7160) );
  xor2_1 U5808 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[10]), .ip2(
        n8713), .op(n5538) );
  nor2_1 U5809 ( .ip1(n8965), .ip2(n8934), .op(n5052) );
  nor2_1 U5810 ( .ip1(n9331), .ip2(n8703), .op(n5155) );
  xor2_1 U5811 ( .ip1(n8270), .ip2(n8321), .op(n8322) );
  xor2_1 U5812 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[10]), .ip2(
        n8319), .op(n8320) );
  nand2_2 U5813 ( .ip1(n9444), .ip2(n9424), .op(n9447) );
  nor2_1 U5814 ( .ip1(n7774), .ip2(n7735), .op(n5126) );
  nor2_1 U5815 ( .ip1(n9335), .ip2(n8311), .op(n4154) );
  nor2_1 U5816 ( .ip1(n8518), .ip2(n8511), .op(n5166) );
  nand2_1 U5817 ( .ip1(n9422), .ip2(n9423), .op(n9442) );
  and3_1 U5818 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[13]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[12]), .ip3(n7688), .op(n7689)
         );
  nor2_1 U5819 ( .ip1(n8518), .ip2(n8506), .op(n5169) );
  and2_1 U5820 ( .ip1(n8330), .ip2(n8329), .op(n8331) );
  nand2_1 U5821 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[3]), .ip2(
        n8308), .op(n8310) );
  and2_1 U5822 ( .ip1(n7696), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[11]), .op(n7688) );
  xnor2_1 U5823 ( .ip1(n7719), .ip2(n7718), .op(n7720) );
  and2_1 U5824 ( .ip1(n8522), .ip2(n8521), .op(n8523) );
  and2_1 U5825 ( .ip1(n9394), .ip2(n9393), .op(n5569) );
  nand2_1 U5826 ( .ip1(n9406), .ip2(n9441), .op(n9403) );
  nor2_1 U5827 ( .ip1(n8613), .ip2(n8612), .op(n8623) );
  nor2_1 U5828 ( .ip1(n6963), .ip2(n6962), .op(n6975) );
  xnor2_1 U5829 ( .ip1(n5579), .ip2(i_i2c_ic_sda_tx_hold_sync[13]), .op(n9406)
         );
  xnor2_1 U5830 ( .ip1(n5580), .ip2(i_i2c_ic_sda_tx_hold_sync[11]), .op(n9398)
         );
  and2_1 U5831 ( .ip1(n8626), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[11]), .op(n8627) );
  xnor2_1 U5832 ( .ip1(n5526), .ip2(n5525), .op(n5524) );
  nor4_1 U5833 ( .ip1(n6298), .ip2(n6297), .ip3(n6296), .ip4(n6295), .op(n6299) );
  inv_2 U5834 ( .ip(n8757), .op(n5273) );
  xnor2_1 U5835 ( .ip1(n5518), .ip2(n9231), .op(n9375) );
  nor2_1 U5836 ( .ip1(n6083), .ip2(n6082), .op(n6085) );
  nand4_1 U5837 ( .ip1(n10628), .ip2(n10627), .ip3(n10626), .ip4(n10625), .op(
        n10632) );
  nor3_2 U5838 ( .ip1(n10545), .ip2(n10544), .ip3(n5349), .op(n10587) );
  xnor2_1 U5839 ( .ip1(n8211), .ip2(n8213), .op(n8214) );
  nor2_1 U5840 ( .ip1(n6994), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[0]), 
        .op(n6218) );
  xnor2_1 U5841 ( .ip1(n6207), .ip2(n6206), .op(n8807) );
  nor2_1 U5842 ( .ip1(n6994), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[0]), .op(n8661) );
  and2_1 U5843 ( .ip1(n5944), .ip2(n5943), .op(n5945) );
  nand3_1 U5844 ( .ip1(n8222), .ip2(n8221), .ip3(n8220), .op(n8225) );
  xor2_1 U5845 ( .ip1(n8550), .ip2(n8549), .op(n8408) );
  nand2_2 U5846 ( .ip1(n7180), .ip2(n7179), .op(n9691) );
  and2_1 U5847 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[9]), .ip2(n10489), .op(n5296) );
  inv_2 U5848 ( .ip(n8537), .op(n5275) );
  and2_1 U5849 ( .ip1(n9209), .ip2(n9203), .op(n9204) );
  inv_2 U5850 ( .ip(n8392), .op(n5276) );
  inv_2 U5851 ( .ip(n5310), .op(n10678) );
  and2_1 U5852 ( .ip1(n9197), .ip2(n9152), .op(n9195) );
  inv_2 U5853 ( .ip(n8429), .op(n5278) );
  nand2_1 U5854 ( .ip1(n10672), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[9]), .op(n10549) );
  xnor2_1 U5855 ( .ip1(n6216), .ip2(n6215), .op(n8811) );
  and2_1 U5856 ( .ip1(n9236), .ip2(n9235), .op(n9237) );
  inv_4 U5857 ( .ip(n5443), .op(n5279) );
  nand2_2 U5858 ( .ip1(n6863), .ip2(n6862), .op(n7265) );
  inv_2 U5859 ( .ip(n9686), .op(n11122) );
  and2_1 U5860 ( .ip1(n9281), .ip2(n9280), .op(n9283) );
  buf_1 U5861 ( .ip(n6054), .op(n6158) );
  nand2_1 U5862 ( .ip1(n6052), .ip2(n6184), .op(n6172) );
  nor2_1 U5863 ( .ip1(n8262), .ip2(n8265), .op(n8168) );
  buf_1 U5864 ( .ip(n6214), .op(n6215) );
  inv_1 U5865 ( .ip(n10539), .op(n10551) );
  nand2_1 U5866 ( .ip1(n7027), .ip2(n7094), .op(n7028) );
  nand2_1 U5867 ( .ip1(n6183), .ip2(n6185), .op(n6052) );
  inv_4 U5868 ( .ip(n10538), .op(n5281) );
  nand2_1 U5869 ( .ip1(n5949), .ip2(n5948), .op(n5534) );
  inv_1 U5870 ( .ip(n6076), .op(n6185) );
  nand2_2 U5871 ( .ip1(n5431), .ip2(n5432), .op(n8229) );
  mux2_2 U5872 ( .ip1(i_i2c_ic_fs_lcnt[0]), .ip2(i_i2c_ic_lcnt[0]), .s(n6041), 
        .op(n7121) );
  inv_1 U5873 ( .ip(n5947), .op(n5948) );
  inv_1 U5874 ( .ip(n7391), .op(n11855) );
  nand2_1 U5875 ( .ip1(i_i2c_ic_fs_hcnt[0]), .ip2(n5430), .op(n5431) );
  nor2_1 U5876 ( .ip1(n11836), .ip2(n6035), .op(n6036) );
  nand2_2 U5877 ( .ip1(n10084), .ip2(n6852), .op(
        i_apb_U_DW_apb_ahbsif_nextstate[0]) );
  inv_2 U5878 ( .ip(n10479), .op(n5283) );
  and2_1 U5879 ( .ip1(n11835), .ip2(n9562), .op(n9563) );
  and2_1 U5880 ( .ip1(i_i2c_scl_lcnt_cmplt), .ip2(n5591), .op(n7776) );
  and2_1 U5881 ( .ip1(n11835), .ip2(n8090), .op(n8091) );
  inv_2 U5882 ( .ip(n7386), .op(n5284) );
  nand2_2 U5883 ( .ip1(n5857), .ip2(n5856), .op(i_i2c_hs_mcode_en) );
  inv_4 U5884 ( .ip(n6454), .op(n5285) );
  nor2_1 U5885 ( .ip1(n5531), .ip2(n5528), .op(n5530) );
  and2_1 U5886 ( .ip1(n11335), .ip2(i_i2c_rx_wr_addr[1]), .op(n11167) );
  nand2_1 U5887 ( .ip1(n5471), .ip2(n5859), .op(n5473) );
  and2_1 U5888 ( .ip1(n9948), .ip2(n10802), .op(n9941) );
  and2_1 U5889 ( .ip1(n9602), .ip2(n9601), .op(n9603) );
  mux2_1 U5890 ( .ip1(i_apb_pwdata_int[1]), .ip2(i_ssi_baudr[1]), .s(n9746), 
        .op(n4626) );
  mux2_1 U5891 ( .ip1(i_apb_pwdata_int[8]), .ip2(i_ssi_U_regfile_ctrlr1_int[8]), .s(n9903), .op(n4611) );
  mux2_1 U5892 ( .ip1(i_apb_pwdata_int[7]), .ip2(i_ssi_U_regfile_ctrlr1_int[7]), .s(n9903), .op(n4596) );
  mux2_1 U5893 ( .ip1(i_apb_pwdata_int[6]), .ip2(i_ssi_U_regfile_ctrlr1_int[6]), .s(n9903), .op(n4597) );
  nand2_2 U5894 ( .ip1(n11162), .ip2(n6828), .op(n7413) );
  inv_1 U5895 ( .ip(n5858), .op(n5859) );
  and2_1 U5896 ( .ip1(n5375), .ip2(n5376), .op(n5378) );
  nand2_2 U5897 ( .ip1(n5377), .ip2(n5375), .op(n9883) );
  nand2_1 U5898 ( .ip1(n5250), .ip2(n9857), .op(n5308) );
  nand2_1 U5899 ( .ip1(n9128), .ip2(n9127), .op(n9134) );
  nor2_1 U5900 ( .ip1(n7352), .ip2(n7348), .op(n5366) );
  nor2_1 U5901 ( .ip1(n6431), .ip2(n6430), .op(n6442) );
  nor2_1 U5902 ( .ip1(n5757), .ip2(n10118), .op(n5762) );
  inv_1 U5903 ( .ip(n9879), .op(n5375) );
  inv_1 U5904 ( .ip(n10682), .op(n5328) );
  nand2_1 U5905 ( .ip1(n9122), .ip2(n9121), .op(n9128) );
  inv_1 U5906 ( .ip(n10568), .op(n5287) );
  nor2_1 U5907 ( .ip1(n5755), .ip2(i_ssi_mwcr[0]), .op(n5756) );
  nor2_1 U5908 ( .ip1(n6426), .ip2(n6425), .op(n6427) );
  and4_1 U5909 ( .ip1(n5251), .ip2(n5379), .ip3(n5381), .ip4(n5380), .op(n5636) );
  or2_1 U5910 ( .ip1(n5715), .ip2(n5713), .op(n5505) );
  inv_1 U5911 ( .ip(n5951), .op(n5528) );
  nor2_1 U5912 ( .ip1(n5800), .ip2(n5439), .op(n5714) );
  nand2_1 U5913 ( .ip1(n7356), .ip2(n5606), .op(n7378) );
  and2_1 U5914 ( .ip1(n11638), .ip2(n11637), .op(n11639) );
  and2_1 U5915 ( .ip1(n10926), .ip2(n8328), .op(n5843) );
  inv_1 U5916 ( .ip(n5624), .op(n5379) );
  inv_1 U5917 ( .ip(n10430), .op(n5380) );
  nand2_1 U5918 ( .ip1(n5702), .ip2(n5701), .op(n5800) );
  and2_1 U5919 ( .ip1(n7152), .ip2(n7153), .op(n7154) );
  mux2_2 U5920 ( .ip1(i_i2c_ic_fs_lcnt[6]), .ip2(i_i2c_ic_lcnt[6]), .s(n5907), 
        .op(n5915) );
  inv_1 U5921 ( .ip(n10701), .op(n5339) );
  mux2_2 U5922 ( .ip1(i_i2c_ic_fs_lcnt[8]), .ip2(i_i2c_ic_lcnt[8]), .s(n5907), 
        .op(n5949) );
  xor2_1 U5923 ( .ip1(i_ssi_baudr[15]), .ip2(n6393), .op(n6394) );
  and2_1 U5924 ( .ip1(n7164), .ip2(n7165), .op(n7161) );
  nor2_1 U5925 ( .ip1(n5700), .ip2(n10429), .op(n5389) );
  inv_1 U5926 ( .ip(n5648), .op(n5417) );
  and2_1 U5927 ( .ip1(n9853), .ip2(n6031), .op(n5727) );
  nor2_2 U5928 ( .ip1(n5303), .ip2(n5302), .op(n5761) );
  inv_1 U5929 ( .ip(n6353), .op(n5471) );
  inv_1 U5930 ( .ip(n5335), .op(n9851) );
  xor2_2 U5931 ( .ip1(n5667), .ip2(n5658), .op(n5659) );
  and2_1 U5932 ( .ip1(n8350), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[3]), .op(n7152) );
  inv_1 U5933 ( .ip(n5513), .op(n5718) );
  xnor2_1 U5934 ( .ip1(n5680), .ip2(n5679), .op(n5692) );
  or2_1 U5935 ( .ip1(n5335), .ip2(i_ssi_U_mstfsm_abort_ir), .op(n5798) );
  and2_1 U5936 ( .ip1(n7481), .ip2(n7480), .op(n7482) );
  inv_1 U5937 ( .ip(n10418), .op(n5288) );
  xnor2_1 U5938 ( .ip1(n5682), .ip2(n5681), .op(n5691) );
  xor2_2 U5939 ( .ip1(n5642), .ip2(n5641), .op(n5649) );
  xor2_2 U5940 ( .ip1(n5640), .ip2(n5639), .op(n5650) );
  xor2_2 U5941 ( .ip1(n5646), .ip2(n5645), .op(n5647) );
  nand2_1 U5942 ( .ip1(n5318), .ip2(n9902), .op(n5709) );
  nor2_1 U5943 ( .ip1(n5299), .ip2(i_ssi_ssi_en_int), .op(n5777) );
  nor4_4 U5944 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(i_ahb_U_mux_hsel_prev[3]), .ip3(i_ahb_U_mux_hsel_prev[2]), .ip4(n6511), .op(n11154) );
  and2_1 U5945 ( .ip1(n10802), .ip2(n10801), .op(n10803) );
  nand2_1 U5946 ( .ip1(n5316), .ip2(n5315), .op(n9854) );
  inv_1 U5947 ( .ip(n10029), .op(n5395) );
  inv_1 U5948 ( .ip(n6069), .op(n5412) );
  nand2_1 U5949 ( .ip1(n7329), .ip2(n6383), .op(n6423) );
  xor2_2 U5950 ( .ip1(i_i2c_U_DW_apb_i2c_intctl_slv_clr_leftover_flg_sync), 
        .ip2(i_i2c_U_DW_apb_i2c_intctl_slv_clr_leftover_flg_sync_q), .op(n7398) );
  inv_1 U5951 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[13]), .op(n5470)
         );
  and2_1 U5952 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[4]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[5]), .op(n7153) );
  xor2_2 U5953 ( .ip1(i_ssi_cfs[1]), .ip2(i_ssi_U_mstfsm_ctrl_cnt[1]), .op(
        n6928) );
  xnor2_1 U5954 ( .ip1(i_ssi_U_mstfsm_bit_cnt[3]), .ip2(i_ssi_dfs[3]), .op(
        n5602) );
  nand2_1 U5955 ( .ip1(i_ssi_tx_rd_addr[0]), .ip2(i_ssi_tx_rd_addr[2]), .op(
        n10234) );
  inv_1 U5956 ( .ip(i_ssi_cfs[3]), .op(n5311) );
  inv_1 U5957 ( .ip(i_ssi_cfs[1]), .op(n10438) );
  and2_1 U5958 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[6]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[7]), .op(n6007) );
  and2_1 U5959 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[4]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[3]), .op(n6006) );
  buf_1 U5960 ( .ip(i_ssi_U_mstfsm_frame_cnt[16]), .op(n5320) );
  nand3_1 U5961 ( .ip1(i_ssi_U_mstfsm_c_state[3]), .ip2(
        i_ssi_U_mstfsm_c_state[1]), .ip3(i_ssi_U_mstfsm_c_state[0]), .op(n5299) );
  inv_1 U5962 ( .ip(i_ssi_U_shift_U_tx_shifter_tx_buffer[15]), .op(n5331) );
  and2_1 U5963 ( .ip1(ex_i_ahb_AHB_Slave_PID_hready_resp), .ip2(
        i_ahb_U_mux_hsel_prev[4]), .op(n6683) );
  inv_1 U5964 ( .ip(i_i2c_ic_sda_tx_hold_sync[10]), .op(n5525) );
  inv_1 U5965 ( .ip(i_ssi_sclk_fe), .op(n5315) );
  inv_1 U5966 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_scl_clk_int), .op(n5472) );
  and3_1 U5967 ( .ip1(n6824), .ip2(n6823), .ip3(n6822), .op(n6825) );
  nand3_2 U5968 ( .ip1(n10420), .ip2(n10419), .ip3(n5292), .op(n10424) );
  nand2_1 U5969 ( .ip1(n10424), .ip2(n10423), .op(n10589) );
  and2_1 U5970 ( .ip1(n10589), .ip2(n10416), .op(n5333) );
  inv_1 U5971 ( .ip(n9846), .op(n10419) );
  nor2_2 U5972 ( .ip1(n9849), .ip2(n9848), .op(n10420) );
  nor2_2 U5973 ( .ip1(n10418), .ip2(n10417), .op(n5292) );
  nand2_4 U5974 ( .ip1(n10443), .ip2(n5309), .op(n5360) );
  nand2_2 U5975 ( .ip1(n5323), .ip2(n10860), .op(n5309) );
  nand2_1 U5976 ( .ip1(n5294), .ip2(n5293), .op(n4394) );
  nand2_1 U5977 ( .ip1(n5296), .ip2(n5297), .op(n5293) );
  nand2_1 U5978 ( .ip1(n5295), .ip2(n10490), .op(n5294) );
  nand2_1 U5979 ( .ip1(n10489), .ip2(n5297), .op(n5295) );
  nand2_1 U5980 ( .ip1(n5423), .ip2(n10487), .op(n5298) );
  nand2_4 U5981 ( .ip1(n10460), .ip2(n10459), .op(n10516) );
  inv_1 U5982 ( .ip(n5300), .op(n5781) );
  nand2_1 U5983 ( .ip1(n5761), .ip2(n5301), .op(n5300) );
  inv_1 U5984 ( .ip(n5768), .op(n5301) );
  inv_1 U5985 ( .ip(n5508), .op(n5304) );
  nand2_4 U5986 ( .ip1(n5409), .ip2(n5410), .op(n10538) );
  nand2_4 U5987 ( .ip1(n5408), .ip2(n10441), .op(n5409) );
  nand2_1 U5988 ( .ip1(n5497), .ip2(n5796), .op(n5323) );
  nand2_2 U5989 ( .ip1(n5304), .ip2(n5311), .op(n10443) );
  nand2_1 U5990 ( .ip1(n5305), .ip2(n9857), .op(n5306) );
  inv_1 U5991 ( .ip(n9852), .op(n5305) );
  nand2_2 U5992 ( .ip1(n5307), .ip2(n5306), .op(n10440) );
  inv_1 U5993 ( .ip(n5444), .op(n5498) );
  nand2_2 U5994 ( .ip1(n5804), .ip2(n5444), .op(n5312) );
  nand2_4 U5995 ( .ip1(n5787), .ip2(n5512), .op(n5444) );
  nand2_1 U5996 ( .ip1(n5402), .ip2(n10737), .op(n5313) );
  nand2_2 U5997 ( .ip1(n5511), .ip2(n10438), .op(n5314) );
  inv_1 U5998 ( .ip(n5387), .op(n5422) );
  or2_1 U5999 ( .ip1(n10550), .ip2(n5325), .op(n5387) );
  nand2_1 U6000 ( .ip1(n5448), .ip2(n5449), .op(n5325) );
  nand2_1 U6001 ( .ip1(n5402), .ip2(n11471), .op(n5449) );
  nand2_1 U6002 ( .ip1(n5447), .ip2(n10437), .op(n5448) );
  nand2_4 U6003 ( .ip1(n5314), .ip2(n5313), .op(n10550) );
  inv_1 U6004 ( .ip(i_ssi_baud2), .op(n5316) );
  not_ab_or_c_or_d U6005 ( .ip1(n5319), .ip2(i_ssi_U_regfile_ctrlr1_int[15]), 
        .ip3(n5321), .ip4(n5317), .op(n5711) );
  nor2_2 U6006 ( .ip1(n5320), .ip2(i_ssi_U_regfile_ctrlr1_int[15]), .op(n5317)
         );
  buf_1 U6007 ( .ip(i_ssi_U_regfile_ctrlr1_int[15]), .op(n5318) );
  nor2_1 U6008 ( .ip1(n5710), .ip2(i_ssi_U_mstfsm_frame_cnt[15]), .op(n5319)
         );
  nand2_1 U6009 ( .ip1(n10424), .ip2(n10423), .op(n5322) );
  and2_1 U6010 ( .ip1(n10443), .ip2(n5309), .op(n5324) );
  nor2_2 U6011 ( .ip1(n5405), .ip2(n5503), .op(n5497) );
  nand2_2 U6012 ( .ip1(n10678), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[4]), .op(n10600) );
  nor2_2 U6013 ( .ip1(i_ssi_U_shift_U_tx_shifter_load_start_bit_ir), .ip2(
        n10479), .op(n10677) );
  nand2_1 U6014 ( .ip1(n5448), .ip2(n5449), .op(n10539) );
  inv_1 U6015 ( .ip(i_ssi_dfs[3]), .op(n5326) );
  inv_1 U6016 ( .ip(n5326), .op(n5327) );
  or2_1 U6017 ( .ip1(n10609), .ip2(n5328), .op(n10684) );
  inv_1 U6018 ( .ip(n5440), .op(n10683) );
  nand2_1 U6019 ( .ip1(n5505), .ip2(n5504), .op(n5503) );
  inv_1 U6020 ( .ip(n5502), .op(n5330) );
  or2_2 U6021 ( .ip1(n10703), .ip2(n5742), .op(n5743) );
  inv_2 U6022 ( .ip(n5445), .op(n5748) );
  or2_1 U6023 ( .ip1(n10609), .ip2(n5331), .op(n10627) );
  inv_1 U6024 ( .ip(n10609), .op(n10660) );
  and2_1 U6025 ( .ip1(n10614), .ip2(n10689), .op(n10621) );
  or2_1 U6026 ( .ip1(n5337), .ip2(n5332), .op(n10547) );
  inv_1 U6027 ( .ip(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[5]), .op(n5332) );
  inv_2 U6028 ( .ip(n5493), .op(n5796) );
  nand2_2 U6029 ( .ip1(n10689), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[14]), 
        .op(n10626) );
  and2_1 U6030 ( .ip1(n10416), .ip2(n5322), .op(n5487) );
  nor2_2 U6031 ( .ip1(n5739), .ip2(n5740), .op(n5334) );
  nor2_1 U6032 ( .ip1(n5739), .ip2(n5740), .op(n5744) );
  nor2_1 U6033 ( .ip1(n10588), .ip2(n10587), .op(n10606) );
  nor2_2 U6034 ( .ip1(i_ssi_tmod[1]), .ip2(n5336), .op(n5335) );
  inv_1 U6035 ( .ip(i_ssi_tmod[1]), .op(n10429) );
  nand2_1 U6036 ( .ip1(n5360), .ip2(n5281), .op(n5337) );
  nand2_2 U6037 ( .ip1(n5718), .ip2(n5339), .op(n5338) );
  inv_1 U6038 ( .ip(n5338), .op(n5809) );
  nand2_1 U6039 ( .ip1(n5734), .ip2(n5340), .op(n5737) );
  or2_1 U6040 ( .ip1(i_ssi_load_start_bit), .ip2(n5287), .op(n5342) );
  inv_1 U6041 ( .ip(n5322), .op(n5341) );
  or2_1 U6042 ( .ip1(n5341), .ip2(n5287), .op(n10591) );
  mux2_1 U6043 ( .ip1(i_apb_pwdata_int[9]), .ip2(n5383), .s(n9903), .op(n4610)
         );
  xor2_2 U6044 ( .ip1(i_ssi_U_mstfsm_frame_cnt[7]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[7]), .op(n5687) );
  inv_1 U6045 ( .ip(n5486), .op(n5478) );
  inv_1 U6046 ( .ip(n11471), .op(n5343) );
  nand2_1 U6047 ( .ip1(n5334), .ip2(n5743), .op(n5344) );
  nand3_1 U6048 ( .ip1(n5754), .ip2(n9853), .ip3(n5388), .op(n5764) );
  xnor2_2 U6049 ( .ip1(i_ssi_dfs[0]), .ip2(i_ssi_U_mstfsm_bit_cnt[0]), .op(
        n5760) );
  nand2_1 U6050 ( .ip1(n5744), .ip2(n5743), .op(n5405) );
  inv_1 U6051 ( .ip(n5491), .op(n5345) );
  inv_1 U6052 ( .ip(n5499), .op(n5500) );
  nand2_1 U6053 ( .ip1(n5797), .ip2(n5722), .op(n5346) );
  inv_1 U6054 ( .ip(n5346), .op(n5813) );
  nor2_4 U6055 ( .ip1(n7164), .ip2(n9890), .op(n9898) );
  nand3_4 U6056 ( .ip1(n9898), .ip2(i_ssi_U_mstfsm_frame_cnt[15]), .ip3(
        i_ssi_U_mstfsm_frame_cnt[14]), .op(n9899) );
  inv_1 U6057 ( .ip(n5401), .op(n5347) );
  nor2_1 U6058 ( .ip1(n10540), .ip2(n5348), .op(n10457) );
  nand2_1 U6059 ( .ip1(n5398), .ip2(n5287), .op(n5348) );
  nand2_1 U6060 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[1]), .ip2(
        n10633), .op(n10548) );
  inv_2 U6061 ( .ip(n5424), .op(n5362) );
  nor2_2 U6062 ( .ip1(n5793), .ip2(n5329), .op(n5384) );
  nor2_2 U6063 ( .ip1(i_ssi_baudr[1]), .ip2(i_ssi_baudr[2]), .op(n7329) );
  nor2_1 U6064 ( .ip1(n5424), .ip2(n5350), .op(n5349) );
  inv_1 U6065 ( .ip(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[14]), .op(n5350)
         );
  inv_1 U6066 ( .ip(n10737), .op(n5351) );
  inv_1 U6067 ( .ip(i_ssi_dfs[2]), .op(n5352) );
  inv_1 U6068 ( .ip(n5352), .op(n5353) );
  nand2_2 U6069 ( .ip1(n5750), .ip2(n5507), .op(n5740) );
  nand2_1 U6070 ( .ip1(n5512), .ip2(n5354), .op(n5488) );
  inv_1 U6071 ( .ip(i_ssi_U_mstfsm_c_state[2]), .op(n5425) );
  inv_1 U6072 ( .ip(i_ssi_sclk_re), .op(n5426) );
  or4_1 U6073 ( .ip1(n5792), .ip2(n5323), .ip3(n5346), .ip4(n10988), .op(n5355) );
  inv_1 U6074 ( .ip(i_ssi_baudr[2]), .op(n6433) );
  nand2_4 U6075 ( .ip1(n5410), .ip2(n5409), .op(n5357) );
  xor2_2 U6076 ( .ip1(i_ssi_U_mstfsm_frame_cnt[6]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[6]), .op(n5679) );
  inv_1 U6077 ( .ip(n10425), .op(n5358) );
  xor2_2 U6078 ( .ip1(i_ssi_U_mstfsm_frame_cnt[10]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[10]), .op(n5698) );
  nand4_1 U6079 ( .ip1(n10548), .ip2(n10549), .ip3(n10547), .ip4(n10546), .op(
        n5359) );
  nand4_1 U6080 ( .ip1(n10548), .ip2(n10549), .ip3(n10547), .ip4(n10546), .op(
        n10607) );
  or2_1 U6081 ( .ip1(n5424), .ip2(n5361), .op(n10599) );
  inv_1 U6082 ( .ip(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[12]), .op(n5361)
         );
  mux2_1 U6083 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[15]), .ip2(
        n10533), .s(n5363), .op(n4389) );
  or2_1 U6084 ( .ip1(n10531), .ip2(n10532), .op(n5363) );
  nand2_1 U6085 ( .ip1(n5365), .ip2(n5366), .op(n5364) );
  and2_1 U6086 ( .ip1(n7346), .ip2(n7347), .op(n5365) );
  inv_1 U6087 ( .ip(n10550), .op(n5367) );
  inv_1 U6088 ( .ip(n10550), .op(n10540) );
  nand2_1 U6089 ( .ip1(n10437), .ip2(n5447), .op(n5368) );
  inv_1 U6090 ( .ip(n10419), .op(n5369) );
  inv_1 U6091 ( .ip(n5369), .op(n5370) );
  nand2_1 U6092 ( .ip1(n10672), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[10]), .op(n10542) );
  nand2_1 U6093 ( .ip1(n5796), .ip2(n5767), .op(n5371) );
  nand2_1 U6094 ( .ip1(n5796), .ip2(n5767), .op(n10442) );
  not_ab_or_c_or_d U6095 ( .ip1(n5675), .ip2(n5674), .ip3(n5673), .ip4(n5672), 
        .op(n5372) );
  nor2_2 U6096 ( .ip1(n7370), .ip2(i_ssi_baudr[9]), .op(n7371) );
  nand2_2 U6097 ( .ip1(n10550), .ip2(n5398), .op(n5373) );
  nand2_2 U6098 ( .ip1(n10550), .ip2(n5398), .op(n10638) );
  inv_1 U6099 ( .ip(n10629), .op(n5374) );
  and2_1 U6100 ( .ip1(n9886), .ip2(n5376), .op(n5377) );
  inv_1 U6101 ( .ip(n9874), .op(n5376) );
  or2_1 U6102 ( .ip1(n10737), .ip2(n5759), .op(n5381) );
  nand2_1 U6103 ( .ip1(n5635), .ip2(n5636), .op(n9879) );
  inv_1 U6104 ( .ip(i_ssi_U_regfile_ctrlr1_int[9]), .op(n5382) );
  inv_1 U6105 ( .ip(n5382), .op(n5383) );
  xor2_2 U6106 ( .ip1(i_ssi_U_mstfsm_frame_cnt[8]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[8]), .op(n5684) );
  xor2_2 U6107 ( .ip1(i_ssi_U_regfile_ctrlr1_int[9]), .ip2(
        i_ssi_U_mstfsm_frame_cnt[9]), .op(n5681) );
  nand2_1 U6108 ( .ip1(n5387), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[15]), 
        .op(n5385) );
  nand2_1 U6109 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_buffer[3]), .ip2(n5422), 
        .op(n5386) );
  nand2_1 U6110 ( .ip1(n5386), .ip2(n5385), .op(n10595) );
  or2_1 U6111 ( .ip1(n9907), .ip2(n5500), .op(n5388) );
  inv_1 U6112 ( .ip(n5388), .op(n5776) );
  and2_1 U6113 ( .ip1(n5389), .ip2(n5702), .op(n5801) );
  xnor2_1 U6114 ( .ip1(i_ssi_U_regfile_ctrlr1_int[11]), .ip2(n5390), .op(n5695) );
  inv_1 U6115 ( .ip(i_ssi_U_mstfsm_frame_cnt[11]), .op(n5390) );
  or2_1 U6116 ( .ip1(n5392), .ip2(n5424), .op(n10546) );
  inv_1 U6117 ( .ip(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[13]), .op(n5392)
         );
  inv_1 U6118 ( .ip(n5514), .op(n5393) );
  nor2_1 U6119 ( .ip1(n7361), .ip2(n5395), .op(n5394) );
  inv_1 U6120 ( .ip(n5394), .op(n7370) );
  xnor2_1 U6121 ( .ip1(n6424), .ip2(n6397), .op(n6425) );
  and2_1 U6122 ( .ip1(n7320), .ip2(n5355), .op(n11851) );
  nand2_1 U6123 ( .ip1(n5677), .ip2(n5372), .op(n5396) );
  nor2_2 U6124 ( .ip1(n5666), .ip2(n5665), .op(n5677) );
  mux2_2 U6125 ( .ip1(i_apb_pwdata_int[3]), .ip2(i_ssi_U_regfile_ctrlr1_int[3]), .s(n9903), .op(n4600) );
  nand2_2 U6126 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[2]), .ip2(
        n10633), .op(n10543) );
  inv_1 U6127 ( .ip(n5279), .op(n5397) );
  nand2_2 U6128 ( .ip1(n5449), .ip2(n5368), .op(n5398) );
  inv_2 U6129 ( .ip(n10440), .op(n9913) );
  and4_1 U6130 ( .ip1(n7377), .ip2(n7376), .ip3(n7375), .ip4(n7374), .op(n5481) );
  inv_1 U6131 ( .ip(n10118), .op(n5399) );
  inv_1 U6132 ( .ip(n5399), .op(n5400) );
  nand2_2 U6133 ( .ip1(n5367), .ip2(n5398), .op(n5401) );
  inv_4 U6134 ( .ip(n5401), .op(n10689) );
  xor2_2 U6135 ( .ip1(i_ssi_U_mstfsm_frame_cnt[3]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[3]), .op(n5658) );
  nand2_1 U6136 ( .ip1(n5384), .ip2(n5450), .op(n5402) );
  nand2_1 U6137 ( .ip1(n5450), .ip2(n5384), .op(n5509) );
  xnor2_2 U6138 ( .ip1(i_ssi_U_mstfsm_bit_cnt[1]), .ip2(i_ssi_dfs[1]), .op(
        n5758) );
  inv_1 U6139 ( .ip(i_ssi_dfs[1]), .op(n10737) );
  nand4_2 U6140 ( .ip1(n10665), .ip2(n10666), .ip3(n10664), .ip4(n10663), .op(
        n10667) );
  nand2_2 U6141 ( .ip1(n10689), .ip2(n10661), .op(n10664) );
  or2_2 U6142 ( .ip1(n5404), .ip2(n5403), .op(n5750) );
  inv_1 U6143 ( .ip(n5729), .op(n5403) );
  ab_or_c_or_d U6144 ( .ip1(i_ssi_sclk_fe), .ip2(n10977), .ip3(
        i_ssi_U_mstfsm_c_state[0]), .ip4(n10111), .op(n5404) );
  nand2_1 U6145 ( .ip1(n5289), .ip2(n5425), .op(n5406) );
  nand2_1 U6146 ( .ip1(n5335), .ip2(n5407), .op(n5724) );
  inv_1 U6147 ( .ip(n5406), .op(n5407) );
  inv_2 U6148 ( .ip(n5371), .op(n5408) );
  nand2_1 U6149 ( .ip1(n5334), .ip2(n5743), .op(n5793) );
  nand2_1 U6150 ( .ip1(n5360), .ip2(n5357), .op(n10648) );
  nor2_2 U6151 ( .ip1(n6158), .ip2(n6055), .op(n6077) );
  nor2_4 U6152 ( .ip1(n8211), .ip2(n6051), .op(n6076) );
  nand2_1 U6153 ( .ip1(n5469), .ip2(n5411), .op(n6063) );
  nor2_1 U6154 ( .ip1(n5412), .ip2(n6070), .op(n5411) );
  xnor2_2 U6155 ( .ip1(n6093), .ip2(n6091), .op(n8778) );
  nand2_1 U6156 ( .ip1(n5469), .ip2(n6069), .op(n5413) );
  nor3_2 U6157 ( .ip1(n5972), .ip2(n5971), .ip3(n6487), .op(n5973) );
  nor2_2 U6158 ( .ip1(n7729), .ip2(n7727), .op(i_i2c_U_DW_apb_i2c_clk_gen_N74)
         );
  xnor2_2 U6159 ( .ip1(n6100), .ip2(n8173), .op(n8773) );
  xor2_1 U6160 ( .ip1(n5414), .ip2(n7373), .op(n7374) );
  xor2_1 U6161 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[12]), .ip2(i_ssi_baudr[12]), 
        .op(n5414) );
  nand2_1 U6162 ( .ip1(n10487), .ip2(n5423), .op(n5415) );
  nand2_4 U6163 ( .ip1(n5814), .ip2(n5247), .op(n10987) );
  inv_2 U6164 ( .ip(n7319), .op(n5814) );
  nand2_1 U6165 ( .ip1(n5487), .ip2(n10440), .op(n5416) );
  nand2_1 U6166 ( .ip1(n5333), .ip2(n10440), .op(n10467) );
  nand4_2 U6167 ( .ip1(n5650), .ip2(n5649), .ip3(n5417), .ip4(n5647), .op(
        n9848) );
  inv_1 U6168 ( .ip(i_ssi_U_regfile_ctrlr1_int[5]), .op(n5418) );
  inv_1 U6169 ( .ip(n5418), .op(n5419) );
  nor2_1 U6170 ( .ip1(n10541), .ip2(n5337), .op(n10545) );
  nand2_1 U6171 ( .ip1(n10672), .ip2(n10673), .op(n5420) );
  nand2_1 U6172 ( .ip1(n5421), .ip2(n10674), .op(n10675) );
  inv_1 U6173 ( .ip(n5420), .op(n5421) );
  nor2_2 U6174 ( .ip1(n5325), .ip2(n10550), .op(n10590) );
  inv_1 U6175 ( .ip(n10540), .op(n5423) );
  nand2_1 U6176 ( .ip1(i_ssi_baud2), .ip2(n10114), .op(n5734) );
  mux2_2 U6177 ( .ip1(n5428), .ip2(n6044), .s(n6043), .op(n5427) );
  inv_1 U6178 ( .ip(i_i2c_ic_hcnt[7]), .op(n5428) );
  nor2_1 U6179 ( .ip1(n8205), .ip2(n8206), .op(n8210) );
  nand2_1 U6180 ( .ip1(n5559), .ip2(n5429), .op(n8272) );
  nand2_1 U6181 ( .ip1(i_i2c_ic_hcnt[0]), .ip2(n6060), .op(n5432) );
  inv_1 U6182 ( .ip(n6060), .op(n5430) );
  nand2_1 U6183 ( .ip1(n8229), .ip2(i_i2c_ic_fs_spklen[0]), .op(n6214) );
  nor2_1 U6184 ( .ip1(n8204), .ip2(n8208), .op(n8205) );
  inv_1 U6185 ( .ip(i_ssi_U_regfile_ctrlr1_int[15]), .op(n5433) );
  inv_1 U6186 ( .ip(n5433), .op(n5434) );
  nor2_1 U6187 ( .ip1(n7397), .ip2(n5291), .op(n5435) );
  nand2_2 U6188 ( .ip1(n5483), .ip2(n10458), .op(n10501) );
  nor2_4 U6189 ( .ip1(n10446), .ip2(n10469), .op(n10447) );
  nand2_2 U6190 ( .ip1(n10503), .ip2(n10504), .op(n5436) );
  nand2_1 U6191 ( .ip1(n10504), .ip2(n10503), .op(n5437) );
  inv_1 U6192 ( .ip(n5324), .op(n5438) );
  nand2_4 U6193 ( .ip1(n9889), .ip2(i_ssi_U_mstfsm_frame_cnt[9]), .op(n9890)
         );
  inv_2 U6194 ( .ip(n10501), .op(n10459) );
  mux2_1 U6195 ( .ip1(i_apb_pwdata_int[11]), .ip2(n5391), .s(n9903), .op(n4608) );
  mux2_1 U6196 ( .ip1(i_apb_pwdata_int[5]), .ip2(n5419), .s(n9903), .op(n4598)
         );
  or4_1 U6197 ( .ip1(n5692), .ip2(n5691), .ip3(n5690), .ip4(n5689), .op(n5439)
         );
  inv_1 U6198 ( .ip(n10590), .op(n5440) );
  inv_1 U6199 ( .ip(n10590), .op(n10609) );
  nand2_1 U6200 ( .ip1(n5324), .ip2(n5357), .op(n5441) );
  nand2_2 U6201 ( .ip1(n5442), .ip2(n10579), .op(n10502) );
  inv_1 U6202 ( .ip(n5441), .op(n5442) );
  inv_1 U6203 ( .ip(n10467), .op(n10579) );
  nand2_2 U6204 ( .ip1(n10550), .ip2(n10551), .op(n5443) );
  inv_2 U6205 ( .ip(n9847), .op(n9849) );
  nand2_2 U6206 ( .ip1(i_ssi_mwcr[1]), .ip2(n5444), .op(n5445) );
  nand2_1 U6207 ( .ip1(n5765), .ip2(n5766), .op(n5446) );
  nand2_1 U6208 ( .ip1(n5766), .ip2(n5765), .op(n5493) );
  nor2_2 U6209 ( .ip1(n5329), .ip2(n5344), .op(n5767) );
  inv_1 U6210 ( .ip(n5509), .op(n5447) );
  inv_1 U6211 ( .ip(n5450), .op(n5451) );
  inv_1 U6212 ( .ip(n5451), .op(n5452) );
  inv_1 U6213 ( .ip(n10860), .op(n5453) );
  nor2_1 U6214 ( .ip1(n5737), .ip2(n5490), .op(n5489) );
  inv_1 U6215 ( .ip(n5500), .op(n10118) );
  inv_1 U6216 ( .ip(i_i2c_ic_fs_hcnt[3]), .op(n5456) );
  inv_1 U6217 ( .ip(i_i2c_ic_hcnt[3]), .op(n5457) );
  inv_1 U6218 ( .ip(n5454), .op(n6129) );
  inv_1 U6219 ( .ip(n5461), .op(n5459) );
  nor2_1 U6220 ( .ip1(n5465), .ip2(n8268), .op(n8193) );
  nor2_2 U6221 ( .ip1(n8388), .ip2(n8370), .op(n5137) );
  nand2_4 U6222 ( .ip1(n7630), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[2]), .op(n7628) );
  inv_1 U6223 ( .ip(i_i2c_ic_fs_hcnt[6]), .op(n5462) );
  inv_1 U6224 ( .ip(i_i2c_ic_hcnt[6]), .op(n5463) );
  inv_2 U6225 ( .ip(n6060), .op(n6043) );
  nor2_1 U6226 ( .ip1(n8205), .ip2(n8206), .op(n5466) );
  nand2_1 U6227 ( .ip1(n5467), .ip2(n8210), .op(n5475) );
  and2_1 U6228 ( .ip1(n8317), .ip2(n8209), .op(n5467) );
  inv_1 U6229 ( .ip(n8258), .op(n8203) );
  xnor2_2 U6230 ( .ip1(n7071), .ip2(n7070), .op(n8858) );
  xor2_2 U6231 ( .ip1(n8505), .ip2(n8504), .op(n8506) );
  inv_1 U6232 ( .ip(n8187), .op(n8192) );
  or2_1 U6233 ( .ip1(n5472), .ip2(n5840), .op(n5842) );
  and2_2 U6234 ( .ip1(n5844), .ip2(i_i2c_mst_debug_cstate[0]), .op(n7685) );
  nand2_1 U6235 ( .ip1(n8209), .ip2(n5466), .op(n5474) );
  nor2_2 U6236 ( .ip1(n5270), .ip2(n5282), .op(n8165) );
  nand2_1 U6237 ( .ip1(n5427), .ip2(n6046), .op(n6167) );
  or2_1 U6238 ( .ip1(n8287), .ip2(n8288), .op(n5476) );
  nand2_1 U6239 ( .ip1(n8201), .ip2(n8202), .op(n8288) );
  nor2_1 U6240 ( .ip1(n9428), .ip2(n9447), .op(n9449) );
  nor2_1 U6241 ( .ip1(n9469), .ip2(n9451), .op(n4945) );
  nor2_1 U6242 ( .ip1(n8288), .ip2(n8287), .op(n8304) );
  nand2_2 U6243 ( .ip1(n6351), .ip2(i_i2c_mst_debug_cstate[1]), .op(n7779) );
  xnor2_1 U6244 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[11]), 
        .ip2(n9460), .op(n5605) );
  inv_1 U6245 ( .ip(n9796), .op(n5477) );
  nor2_2 U6246 ( .ip1(n5514), .ip2(n5373), .op(n10553) );
  inv_2 U6247 ( .ip(n5485), .op(n5486) );
  inv_1 U6248 ( .ip(n9876), .op(n5479) );
  nand2_2 U6249 ( .ip1(n10445), .ip2(n5486), .op(n5480) );
  inv_4 U6250 ( .ip(n5480), .op(n10469) );
  nand2_2 U6251 ( .ip1(n5481), .ip2(n5482), .op(n9795) );
  inv_1 U6252 ( .ip(n10467), .op(n5483) );
  nor2_2 U6253 ( .ip1(n9794), .ip2(n9795), .op(n7397) );
  nor2_2 U6254 ( .ip1(n5436), .ip2(n10505), .op(n10506) );
  inv_1 U6255 ( .ip(n5751), .op(n5495) );
  or2_1 U6256 ( .ip1(n5727), .ip2(n5345), .op(n5738) );
  nand2_1 U6257 ( .ip1(n10516), .ip2(n5415), .op(n10494) );
  inv_1 U6258 ( .ip(n5284), .op(n5484) );
  or2_1 U6259 ( .ip1(n5288), .ip2(n5499), .op(n5754) );
  inv_1 U6260 ( .ip(n10488), .op(n5485) );
  nand2_1 U6261 ( .ip1(n10231), .ip2(n5488), .op(n5490) );
  inv_1 U6262 ( .ip(n9854), .op(n5491) );
  inv_1 U6263 ( .ip(n9854), .op(n5499) );
  inv_1 U6264 ( .ip(n5290), .op(n5492) );
  inv_1 U6265 ( .ip(i_ssi_start_xfer), .op(n10977) );
  inv_1 U6266 ( .ip(n5752), .op(n5494) );
  nor2_2 U6267 ( .ip1(n5495), .ip2(n5496), .op(n5766) );
  nand2_1 U6268 ( .ip1(n5750), .ip2(n5494), .op(n5496) );
  inv_2 U6269 ( .ip(i_ssi_baud2), .op(n5512) );
  inv_1 U6270 ( .ip(n5498), .op(n9815) );
  inv_1 U6271 ( .ip(n5330), .op(n5501) );
  inv_1 U6272 ( .ip(n5491), .op(n5502) );
  inv_1 U6273 ( .ip(n5503), .op(n5745) );
  or2_2 U6274 ( .ip1(n5708), .ip2(n5747), .op(n5504) );
  nand2_1 U6275 ( .ip1(n5724), .ip2(n5723), .op(n5506) );
  inv_1 U6276 ( .ip(n5506), .op(n5507) );
  xnor2_1 U6277 ( .ip1(n6432), .ip2(n6428), .op(n6429) );
  nand2_1 U6278 ( .ip1(n5497), .ip2(n5796), .op(n5508) );
  inv_1 U6279 ( .ip(i_ssi_start_xfer), .op(n5510) );
  inv_4 U6280 ( .ip(n10638), .op(n10681) );
  inv_1 U6281 ( .ip(n5509), .op(n5511) );
  xor2_2 U6282 ( .ip1(n9791), .ip2(n6394), .op(n6446) );
  inv_1 U6283 ( .ip(n5512), .op(n5513) );
  nor2_2 U6284 ( .ip1(n5416), .ip2(n10553), .op(n10530) );
  xor2_2 U6285 ( .ip1(n6034), .ip2(n9895), .op(n6035) );
  inv_4 U6286 ( .ip(n6337), .op(n10354) );
  xnor2_2 U6287 ( .ip1(n5579), .ip2(i_i2c_ic_sda_tx_hold_sync[13]), .op(n5516)
         );
  nand2_1 U6288 ( .ip1(n9383), .ip2(n9382), .op(n5517) );
  or2_1 U6289 ( .ip1(n9228), .ip2(n9227), .op(n5518) );
  and2_1 U6290 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[10]), .ip2(
        n5524), .op(n5519) );
  nand2_1 U6291 ( .ip1(n9178), .ip2(n5522), .op(n5520) );
  nand2_1 U6292 ( .ip1(n5520), .ip2(n5521), .op(n9255) );
  or2_1 U6293 ( .ip1(i_i2c_ic_sda_tx_hold_sync[1]), .ip2(n9179), .op(n5521) );
  and2_1 U6294 ( .ip1(n9177), .ip2(n5539), .op(n5522) );
  nor4_2 U6295 ( .ip1(n5831), .ip2(n5830), .ip3(n5829), .ip4(n5828), .op(n5837) );
  nand2_1 U6296 ( .ip1(n9204), .ip2(n5567), .op(n5584) );
  nand2_1 U6297 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[12]), 
        .ip2(n5582), .op(n5523) );
  nor2_1 U6298 ( .ip1(n9232), .ip2(n9239), .op(n9233) );
  nor4_2 U6299 ( .ip1(n7454), .ip2(n5822), .ip3(n5821), .ip4(n7457), .op(n5826) );
  inv_1 U6300 ( .ip(n5524), .op(n9396) );
  nand2_1 U6301 ( .ip1(n9283), .ip2(n5567), .op(n5526) );
  xnor2_2 U6302 ( .ip1(n9237), .ip2(n9238), .op(n9374) );
  nand2_1 U6303 ( .ip1(n9195), .ip2(n5567), .op(n9196) );
  or2_1 U6304 ( .ip1(n9165), .ip2(n9186), .op(n9174) );
  mux2_2 U6305 ( .ip1(i_i2c_ic_fs_spklen[2]), .ip2(i_i2c_ic_hs_spklen[2]), .s(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r), .op(n9106) );
  nand2_1 U6306 ( .ip1(n9190), .ip2(n9252), .op(n9191) );
  or2_1 U6307 ( .ip1(n9172), .ip2(n9240), .op(n9166) );
  inv_1 U6308 ( .ip(n9172), .op(n9236) );
  nor2_1 U6309 ( .ip1(n9443), .ip2(n9442), .op(n9444) );
  nor2_1 U6310 ( .ip1(n8290), .ip2(n8310), .op(n8312) );
  xnor2_2 U6311 ( .ip1(n6085), .ip2(n6084), .op(n8620) );
  nor2_2 U6312 ( .ip1(n5459), .ip2(n6053), .op(n6054) );
  nor2_1 U6313 ( .ip1(n7743), .ip2(n6303), .op(n7747) );
  nand2_2 U6314 ( .ip1(n9185), .ip2(n9256), .op(n9252) );
  nor2_2 U6315 ( .ip1(n9154), .ip2(n9132), .op(n9138) );
  and2_2 U6316 ( .ip1(n5927), .ip2(n6466), .op(n5590) );
  xor2_2 U6317 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[6]), .ip2(n7721), .op(n7722) );
  or2_1 U6318 ( .ip1(n7716), .ip2(n6010), .op(n7725) );
  inv_1 U6319 ( .ip(n8226), .op(n8232) );
  inv_1 U6320 ( .ip(i_i2c_ic_fs_hcnt[7]), .op(n6044) );
  xnor2_1 U6321 ( .ip1(n9213), .ip2(n9212), .op(n9388) );
  inv_1 U6322 ( .ip(n6115), .op(n6116) );
  nand2_1 U6323 ( .ip1(n8711), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[9]), .op(n8713) );
  nand2_1 U6324 ( .ip1(n8231), .ip2(n8233), .op(n5548) );
  nand2_1 U6325 ( .ip1(n8217), .ip2(n8218), .op(n8222) );
  nor2_1 U6326 ( .ip1(n8229), .ip2(n8227), .op(n8217) );
  xnor2_1 U6327 ( .ip1(i_i2c_ic_sda_tx_hold_sync[5]), .ip2(n9160), .op(n9163)
         );
  inv_1 U6328 ( .ip(i_i2c_ic_sda_tx_hold_sync[1]), .op(n5539) );
  nand2_1 U6329 ( .ip1(n6205), .ip2(n6071), .op(n6072) );
  nor2_1 U6330 ( .ip1(n7116), .ip2(n7114), .op(n7025) );
  nor2_2 U6331 ( .ip1(n7105), .ip2(n7026), .op(n7094) );
  nor2_1 U6332 ( .ip1(n8251), .ip2(n5589), .op(n8249) );
  nand2_1 U6333 ( .ip1(n8266), .ip2(n5547), .op(n5546) );
  inv_1 U6334 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[11]), .op(n5547)
         );
  nor2_1 U6335 ( .ip1(n5597), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[7]), .op(n8650) );
  nand2_1 U6336 ( .ip1(n5288), .ip2(n9843), .op(n5755) );
  nor2_1 U6337 ( .ip1(n9385), .ip2(n9390), .op(n9386) );
  and2_1 U6338 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[8]), .ip2(
        n9389), .op(n5581) );
  nor2_1 U6339 ( .ip1(n8761), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[10]), .op(n6963) );
  nor2_1 U6340 ( .ip1(n8773), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[14]), .op(n8613) );
  inv_1 U6341 ( .ip(n5950), .op(n5533) );
  or2_1 U6342 ( .ip1(n8200), .ip2(n8269), .op(n8201) );
  nor4_1 U6343 ( .ip1(n9299), .ip2(n9298), .ip3(n9297), .ip4(n9296), .op(n9300) );
  xnor2_1 U6344 ( .ip1(n5568), .ip2(i_i2c_ic_sda_tx_hold_sync[14]), .op(n9402)
         );
  nand2_1 U6345 ( .ip1(n6355), .ip2(n10926), .op(n5853) );
  nand2_1 U6346 ( .ip1(n5489), .ip2(n5738), .op(n5739) );
  nand2_1 U6347 ( .ip1(n5764), .ip2(n5763), .op(n5765) );
  nor4_1 U6348 ( .ip1(n10999), .ip2(n10998), .ip3(n10997), .ip4(n10996), .op(
        n11009) );
  or2_1 U6349 ( .ip1(n9419), .ip2(n9418), .op(n9420) );
  and2_1 U6350 ( .ip1(n9417), .ip2(n9416), .op(n9418) );
  nand2_1 U6351 ( .ip1(n5842), .ip2(n5841), .op(n5858) );
  inv_1 U6352 ( .ip(n9436), .op(n5570) );
  nand2_1 U6353 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[9]), .ip2(
        n8316), .op(n8319) );
  nor2_1 U6354 ( .ip1(n8706), .ip2(n8705), .op(n8711) );
  nand2_1 U6355 ( .ip1(n8702), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[6]), .op(n8705) );
  nor2_1 U6356 ( .ip1(n8689), .ip2(n8688), .op(n8693) );
  nand2_1 U6357 ( .ip1(n8933), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[6]), .op(n8936) );
  nor2_1 U6358 ( .ip1(n6011), .ip2(n7725), .op(n7696) );
  nor4_1 U6359 ( .ip1(n7913), .ip2(n7912), .ip3(n7911), .ip4(n7910), .op(n8987) );
  nor4_1 U6360 ( .ip1(n7843), .ip2(n7842), .ip3(n7841), .ip4(n7840), .op(n7863) );
  inv_1 U6361 ( .ip(i_i2c_ic_sda_tx_hold_sync[6]), .op(n5573) );
  nand2_1 U6362 ( .ip1(i_i2c_ic_sda_tx_hold_sync[7]), .ip2(n9103), .op(n5574)
         );
  nand2_1 U6363 ( .ip1(n9149), .ip2(n9138), .op(n9103) );
  mux2_2 U6364 ( .ip1(i_i2c_ic_fs_spklen[7]), .ip2(i_i2c_ic_hs_spklen[7]), .s(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r), .op(n9101) );
  inv_1 U6365 ( .ip(n6167), .op(n6055) );
  nand2_1 U6366 ( .ip1(n6066), .ip2(n6065), .op(n8227) );
  inv_1 U6367 ( .ip(n9101), .op(n9149) );
  nor2_1 U6368 ( .ip1(n5464), .ip2(n6067), .op(n6211) );
  nand2_1 U6369 ( .ip1(n5464), .ip2(n6067), .op(n6212) );
  and4_1 U6370 ( .ip1(n5548), .ip2(n8226), .ip3(n5549), .ip4(n5550), .op(n8235) );
  inv_1 U6371 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[5]), .op(n5545)
         );
  xnor2_2 U6372 ( .ip1(n9249), .ip2(n9248), .op(n9365) );
  nor2_1 U6373 ( .ip1(n6080), .ip2(n6079), .op(n6108) );
  nor2_1 U6374 ( .ip1(n8258), .ip2(n6125), .op(n6079) );
  nand2_1 U6375 ( .ip1(n6068), .ip2(n6212), .op(n6205) );
  or2_1 U6376 ( .ip1(n6214), .ip2(n6211), .op(n6068) );
  nor2_1 U6377 ( .ip1(n7117), .ip2(n7116), .op(n7115) );
  xnor2_1 U6378 ( .ip1(n5267), .ip2(n8258), .op(n5554) );
  nor4_1 U6379 ( .ip1(n6253), .ip2(n6254), .ip3(n6252), .ip4(n6251), .op(n6257) );
  inv_1 U6380 ( .ip(n7026), .op(n7104) );
  nor2_1 U6381 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[5]), .ip2(n5285), .op(n5939) );
  xnor2_1 U6382 ( .ip1(n6129), .ip2(n6128), .op(n8764) );
  xnor2_1 U6383 ( .ip1(n7062), .ip2(n7061), .op(n8548) );
  xnor2_1 U6384 ( .ip1(n7044), .ip2(n7043), .op(n8536) );
  xnor2_1 U6385 ( .ip1(n7093), .ip2(n7092), .op(n8571) );
  nor2_1 U6386 ( .ip1(n5266), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[7]), .op(n8575) );
  inv_1 U6387 ( .ip(n8435), .op(n8457) );
  xnor2_1 U6388 ( .ip1(n6187), .ip2(n6186), .op(n8800) );
  nor2_1 U6389 ( .ip1(n8800), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[5]), .op(n8671) );
  nor2_1 U6390 ( .ip1(n8651), .ip2(n8650), .op(n8673) );
  nor2_1 U6391 ( .ip1(n8255), .ip2(n5596), .op(n8256) );
  nand2_1 U6392 ( .ip1(n8249), .ip2(n8250), .op(n8257) );
  inv_1 U6393 ( .ip(n5546), .op(n8277) );
  xnor2_1 U6394 ( .ip1(n8265), .ip2(n8264), .op(n8266) );
  nand2_1 U6395 ( .ip1(n9402), .ip2(n9466), .op(n9404) );
  inv_1 U6396 ( .ip(i_i2c_ic_sda_tx_hold_sync[12]), .op(n5583) );
  nor2_1 U6397 ( .ip1(n5268), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[13]), .op(n8404) );
  nor2_1 U6398 ( .ip1(n8858), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[9]), 
        .op(n8423) );
  nor2_1 U6399 ( .ip1(n6941), .ip2(n6940), .op(n6942) );
  mux2_1 U6400 ( .ip1(i_i2c_ic_fs_lcnt[8]), .ip2(i_i2c_ic_lcnt[8]), .s(n6270), 
        .op(n7072) );
  xnor2_1 U6401 ( .ip1(n6119), .ip2(n6118), .op(n8761) );
  inv_1 U6402 ( .ip(n7005), .op(n8822) );
  xnor2_1 U6403 ( .ip1(n6192), .ip2(n6191), .op(n7005) );
  xor2_1 U6404 ( .ip1(i_i2c_ic_fs_spklen[2]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[2]), .op(n5821) );
  nor2_1 U6405 ( .ip1(n5862), .ip2(n5824), .op(n5825) );
  xor2_1 U6406 ( .ip1(i_i2c_ic_hs_spklen[6]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[6]), .op(n5828) );
  xnor2_1 U6407 ( .ip1(n6169), .ip2(n6168), .op(n5597) );
  nor2_1 U6408 ( .ip1(n6165), .ip2(n6164), .op(n6169) );
  nor2_1 U6409 ( .ip1(n7870), .ip2(n7869), .op(n7896) );
  nor2_1 U6410 ( .ip1(n5269), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[11]), .op(n8554) );
  nor2_1 U6411 ( .ip1(n5268), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[13]), .op(n8544) );
  nor2_1 U6412 ( .ip1(n8778), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[13]), .op(n8621) );
  nand2_1 U6413 ( .ip1(n5535), .ip2(n5915), .op(n5531) );
  nand2_1 U6414 ( .ip1(n5761), .ip2(n5762), .op(n5763) );
  nand2_1 U6415 ( .ip1(n5602), .ip2(n5756), .op(n5757) );
  xor2_1 U6416 ( .ip1(n6422), .ip2(i_ssi_baudr[5]), .op(n6424) );
  nor4_1 U6417 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[7]), .ip2(
        i_ssi_U_sclkgen_ssi_cnt[10]), .ip3(i_ssi_U_sclkgen_ssi_cnt[14]), .ip4(
        i_ssi_U_sclkgen_ssi_cnt[12]), .op(n10970) );
  nand2_1 U6418 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[9]), .ip2(
        n9353), .op(n9392) );
  nand2_1 U6419 ( .ip1(n9348), .ip2(n9347), .op(n9405) );
  xnor2_1 U6420 ( .ip1(n6943), .ip2(n6104), .op(n8772) );
  xnor2_1 U6421 ( .ip1(n5912), .ip2(n5911), .op(n5527) );
  nor3_1 U6422 ( .ip1(n5996), .ip2(n6453), .ip3(n5995), .op(n5997) );
  mux2_2 U6423 ( .ip1(n7831), .ip2(n7873), .s(n7830), .op(n7832) );
  nand4_1 U6424 ( .ip1(n5893), .ip2(n5892), .ip3(n5891), .ip4(n7528), .op(
        n5894) );
  inv_1 U6425 ( .ip(n7460), .op(n7562) );
  nand2_1 U6426 ( .ip1(n10216), .ip2(i_ssi_tx_full), .op(n6309) );
  nand2_1 U6427 ( .ip1(i_ssi_tx_pop_sync), .ip2(i_ssi_U_fifo_U_tx_fifo_empty_n), .op(n10216) );
  nor2_1 U6428 ( .ip1(n8183), .ip2(n8182), .op(n8202) );
  nor4_1 U6429 ( .ip1(i_apb_paddr[26]), .ip2(i_apb_paddr[25]), .ip3(
        i_apb_paddr[23]), .ip4(i_apb_paddr[22]), .op(n6022) );
  nor4_1 U6430 ( .ip1(i_apb_paddr[19]), .ip2(i_apb_paddr[21]), .ip3(
        i_apb_paddr[20]), .ip4(i_apb_paddr[18]), .op(n6021) );
  nor4_1 U6431 ( .ip1(i_apb_paddr[17]), .ip2(i_apb_paddr[15]), .ip3(
        i_apb_paddr[14]), .ip4(i_apb_paddr[13]), .op(n6020) );
  nor4_1 U6432 ( .ip1(n9303), .ip2(n9302), .ip3(n9301), .ip4(n9300), .op(n9306) );
  nor2_1 U6433 ( .ip1(n8469), .ip2(n8468), .op(n8490) );
  nor2_1 U6434 ( .ip1(n7779), .ip2(n7778), .op(n7808) );
  nor2_1 U6435 ( .ip1(i_i2c_mst_debug_cstate[0]), .ip2(n11023), .op(n10919) );
  or2_1 U6436 ( .ip1(n6354), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_hcnt_cmplt_int), .op(n5591) );
  nor2_1 U6437 ( .ip1(n6351), .ip2(n7778), .op(n7917) );
  inv_1 U6438 ( .ip(n6502), .op(n5988) );
  xnor2_1 U6439 ( .ip1(n5956), .ip2(n5246), .op(n6498) );
  inv_1 U6440 ( .ip(n6423), .op(n6397) );
  nand2_1 U6441 ( .ip1(n5612), .ip2(n6427), .op(n6431) );
  nor2_1 U6442 ( .ip1(n9436), .ip2(n9458), .op(n9460) );
  inv_1 U6443 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[14]), .op(n8196)
         );
  inv_1 U6444 ( .ip(i_ssi_U_sclkgen_ssi_cnt[3]), .op(n6419) );
  inv_1 U6445 ( .ip(i_ssi_U_sclkgen_ssi_cnt[0]), .op(n9764) );
  nor4_1 U6446 ( .ip1(n10995), .ip2(n10994), .ip3(n10993), .ip4(n10992), .op(
        n11010) );
  nor4_1 U6447 ( .ip1(n11003), .ip2(n11002), .ip3(n11001), .ip4(n11000), .op(
        n11008) );
  nor4_1 U6448 ( .ip1(n9753), .ip2(n9752), .ip3(n9751), .ip4(n9750), .op(
        n10972) );
  nand2_1 U6449 ( .ip1(n10228), .ip2(i_ssi_tx_wr_addr[1]), .op(n10203) );
  nor2_1 U6450 ( .ip1(n8314), .ip2(n8291), .op(n8316) );
  nand2_1 U6451 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[6]), .ip2(
        n8312), .op(n8314) );
  inv_1 U6452 ( .ip(n8330), .op(n9335) );
  inv_1 U6453 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_hcnt_cmplt_int), .op(n8328)
         );
  nor2_1 U6454 ( .ip1(n8697), .ip2(n8696), .op(n8702) );
  nand2_1 U6455 ( .ip1(n8693), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[3]), .op(n8696) );
  and2_1 U6456 ( .ip1(n8385), .ip2(n7154), .op(n5594) );
  nor2_1 U6457 ( .ip1(i_i2c_mst_debug_cstate[3]), .ip2(n8746), .op(n10942) );
  nor2_1 U6458 ( .ip1(n8928), .ip2(n8927), .op(n8933) );
  nor2_1 U6459 ( .ip1(n8920), .ip2(n8919), .op(n8924) );
  nor2_1 U6460 ( .ip1(n7754), .ip2(n6039), .op(n6305) );
  nand2_1 U6461 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[12]), .ip2(
        n7760), .op(n6039) );
  and2_1 U6462 ( .ip1(n7760), .ip2(n7759), .op(n7763) );
  nor2_1 U6463 ( .ip1(n7736), .ip2(n6302), .op(n7739) );
  nand2_1 U6464 ( .ip1(n7771), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[0]), .op(n7736) );
  inv_1 U6465 ( .ip(n7504), .op(n7501) );
  nand2_1 U6466 ( .ip1(n8914), .ip2(n8913), .op(n8962) );
  nand2_1 U6467 ( .ip1(n5591), .ip2(n6356), .op(n9473) );
  inv_1 U6468 ( .ip(n6355), .op(n6356) );
  nand2_1 U6469 ( .ip1(n8683), .ip2(n8682), .op(n8730) );
  nor4_1 U6470 ( .ip1(n8058), .ip2(n8989), .ip3(n8053), .ip4(n8987), .op(n7914) );
  nor4_1 U6471 ( .ip1(n11859), .ip2(n9338), .ip3(n9337), .ip4(n9336), .op(
        n9480) );
  inv_1 U6472 ( .ip(n10122), .op(n10868) );
  nand4_1 U6473 ( .ip1(n10277), .ip2(n10276), .ip3(n10275), .ip4(n10274), .op(
        n10283) );
  nand4_1 U6474 ( .ip1(n10281), .ip2(n10280), .ip3(n10279), .ip4(n10278), .op(
        n10282) );
  nand4_1 U6475 ( .ip1(n10287), .ip2(n10286), .ip3(n10285), .ip4(n10284), .op(
        n10293) );
  nand4_1 U6476 ( .ip1(n10291), .ip2(n10290), .ip3(n10289), .ip4(n10288), .op(
        n10292) );
  nand4_1 U6477 ( .ip1(n10297), .ip2(n10296), .ip3(n10295), .ip4(n10294), .op(
        n10303) );
  nand4_1 U6478 ( .ip1(n10301), .ip2(n10300), .ip3(n10299), .ip4(n10298), .op(
        n10302) );
  nand4_1 U6479 ( .ip1(n10307), .ip2(n10306), .ip3(n10305), .ip4(n10304), .op(
        n10313) );
  nand4_1 U6480 ( .ip1(n10311), .ip2(n10310), .ip3(n10309), .ip4(n10308), .op(
        n10312) );
  nand4_1 U6481 ( .ip1(n10317), .ip2(n10316), .ip3(n10315), .ip4(n10314), .op(
        n10323) );
  nand4_1 U6482 ( .ip1(n10321), .ip2(n10320), .ip3(n10319), .ip4(n10318), .op(
        n10322) );
  nand4_1 U6483 ( .ip1(n10327), .ip2(n10326), .ip3(n10325), .ip4(n10324), .op(
        n10333) );
  nand4_1 U6484 ( .ip1(n10331), .ip2(n10330), .ip3(n10329), .ip4(n10328), .op(
        n10332) );
  nand4_1 U6485 ( .ip1(n10337), .ip2(n10336), .ip3(n10335), .ip4(n10334), .op(
        n10343) );
  nand4_1 U6486 ( .ip1(n10341), .ip2(n10340), .ip3(n10339), .ip4(n10338), .op(
        n10342) );
  nand4_1 U6487 ( .ip1(n10347), .ip2(n10346), .ip3(n10345), .ip4(n10344), .op(
        n10353) );
  nand4_1 U6488 ( .ip1(n10351), .ip2(n10350), .ip3(n10349), .ip4(n10348), .op(
        n10352) );
  nand4_1 U6489 ( .ip1(n10358), .ip2(n10357), .ip3(n10356), .ip4(n10355), .op(
        n10364) );
  nand4_1 U6490 ( .ip1(n10362), .ip2(n10361), .ip3(n10360), .ip4(n10359), .op(
        n10363) );
  nand4_1 U6491 ( .ip1(n10369), .ip2(n10368), .ip3(n10367), .ip4(n10366), .op(
        n10376) );
  nand4_1 U6492 ( .ip1(n10374), .ip2(n10373), .ip3(n10372), .ip4(n10371), .op(
        n10375) );
  nand4_1 U6493 ( .ip1(n10381), .ip2(n10380), .ip3(n10379), .ip4(n10378), .op(
        n10387) );
  nand4_1 U6494 ( .ip1(n10385), .ip2(n10384), .ip3(n10383), .ip4(n10382), .op(
        n10386) );
  nand4_1 U6495 ( .ip1(n10393), .ip2(n10392), .ip3(n10391), .ip4(n10390), .op(
        n10399) );
  nand4_1 U6496 ( .ip1(n10397), .ip2(n10396), .ip3(n10395), .ip4(n10394), .op(
        n10398) );
  nand4_1 U6497 ( .ip1(n10406), .ip2(n10405), .ip3(n10404), .ip4(n10403), .op(
        n10414) );
  nand4_1 U6498 ( .ip1(n10412), .ip2(n10411), .ip3(n10410), .ip4(n10409), .op(
        n10413) );
  nand4_1 U6499 ( .ip1(n10238), .ip2(n10237), .ip3(n10236), .ip4(n10235), .op(
        n10250) );
  nand4_1 U6500 ( .ip1(n10248), .ip2(n10247), .ip3(n10246), .ip4(n10245), .op(
        n10249) );
  inv_1 U6501 ( .ip(n7177), .op(n7180) );
  inv_1 U6502 ( .ip(n11795), .op(i_ssi_ssi_oe_n) );
  inv_1 U6503 ( .ip(n11816), .op(i_ssi_ss_0_n) );
  nor2_1 U6504 ( .ip1(n9335), .ip2(n8313), .op(n4152) );
  nor2_1 U6505 ( .ip1(n9335), .ip2(n8309), .op(n4155) );
  nor2_1 U6506 ( .ip1(n7774), .ip2(n7748), .op(n5121) );
  xor2_1 U6507 ( .ip1(n9463), .ip2(n9462), .op(n5601) );
  xnor2_1 U6508 ( .ip1(i_ssi_U_mstfsm_frame_cnt[16]), .ip2(n9899), .op(n5603)
         );
  xor2_1 U6509 ( .ip1(n8369), .ip2(n8368), .op(n8370) );
  nor2_1 U6510 ( .ip1(n9469), .ip2(n9453), .op(n4944) );
  inv_1 U6511 ( .ip(n5540), .op(n9453) );
  xnor2_1 U6512 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[6]), .ip2(
        n9452), .op(n5540) );
  nor2_1 U6513 ( .ip1(n7774), .ip2(n6308), .op(n5115) );
  nand2_1 U6514 ( .ip1(n6307), .ip2(n6306), .op(n6308) );
  nor2_1 U6515 ( .ip1(n5615), .ip2(n5593), .op(n6307) );
  nand2_1 U6516 ( .ip1(n6277), .ip2(n7758), .op(n6306) );
  inv_1 U6517 ( .ip(n7725), .op(n7695) );
  xor2_1 U6518 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[3]), .ip2(n7716), .op(n7717) );
  nor4_1 U6519 ( .ip1(n6509), .ip2(n6508), .ip3(n6507), .ip4(n11018), .op(
        i_i2c_U_DW_apb_i2c_clk_gen_N51) );
  nor4_1 U6520 ( .ip1(n6506), .ip2(n6505), .ip3(n6504), .ip4(n6503), .op(n6507) );
  xor2_1 U6521 ( .ip1(i_i2c_ic_fs_spklen[5]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[5]), .op(n5822) );
  xor2_1 U6522 ( .ip1(i_i2c_ic_hs_spklen[5]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[5]), .op(n5830) );
  nor2_1 U6523 ( .ip1(n7712), .ip2(n6005), .op(n7714) );
  nor2_2 U6524 ( .ip1(n7729), .ip2(n7728), .op(i_i2c_U_DW_apb_i2c_clk_gen_N76)
         );
  nand2_1 U6525 ( .ip1(n8224), .ip2(n8225), .op(n8226) );
  nor2_2 U6526 ( .ip1(n9331), .ip2(n8701), .op(n5156) );
  xor2_2 U6527 ( .ip1(i_i2c_tx_abrt_flg), .ip2(n11292), .op(n5196) );
  nand2_1 U6528 ( .ip1(n9454), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[8]), .op(n9458) );
  nor2_1 U6529 ( .ip1(n9469), .ip2(n9459), .op(n4941) );
  inv_1 U6530 ( .ip(n5527), .op(n6480) );
  xor2_2 U6531 ( .ip1(n8495), .ip2(n8494), .op(n8496) );
  inv_1 U6532 ( .ip(n5531), .op(n5529) );
  and2_1 U6533 ( .ip1(n5529), .ip2(n5914), .op(n5536) );
  nand2_1 U6534 ( .ip1(n5920), .ip2(n5919), .op(n5913) );
  xor2_2 U6535 ( .ip1(n8915), .ip2(n8962), .op(n8916) );
  xor2_1 U6536 ( .ip1(n6266), .ip2(n7747), .op(n7748) );
  xnor2_2 U6537 ( .ip1(n5533), .ip2(n5534), .op(n5532) );
  inv_1 U6538 ( .ip(n5532), .op(n6488) );
  xor2_1 U6539 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[9]), .ip2(
        n9458), .op(n9459) );
  xor2_2 U6540 ( .ip1(n8510), .ip2(n8509), .op(n8511) );
  xor2_2 U6541 ( .ip1(n8940), .ip2(n8942), .op(n8941) );
  and2_1 U6542 ( .ip1(n5555), .ip2(n5912), .op(n5535) );
  nor2_4 U6543 ( .ip1(n9469), .ip2(n9448), .op(n4947) );
  nor2_2 U6544 ( .ip1(n7774), .ip2(n7734), .op(n5127) );
  nand2_1 U6545 ( .ip1(n6451), .ip2(n5965), .op(n5537) );
  nand2_1 U6546 ( .ip1(n6451), .ip2(n5965), .op(n5994) );
  nor2_2 U6547 ( .ip1(n8388), .ip2(n8378), .op(n5134) );
  xor2_2 U6548 ( .ip1(n8500), .ip2(n8499), .op(n8501) );
  xnor2_2 U6549 ( .ip1(n5964), .ip2(n5963), .op(n6451) );
  nor2_2 U6550 ( .ip1(n8965), .ip2(n8932), .op(n5053) );
  inv_1 U6551 ( .ip(n9181), .op(n9184) );
  nand2_1 U6552 ( .ip1(n5541), .ip2(n5542), .op(n8276) );
  or2_1 U6553 ( .ip1(n5474), .ip2(n5552), .op(n5541) );
  or2_1 U6554 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[9]), .ip2(n5552), 
        .op(n5542) );
  or2_1 U6555 ( .ip1(n8681), .ip2(n5543), .op(n8682) );
  nand2_1 U6556 ( .ip1(n5544), .ip2(n8835), .op(n5543) );
  nand2_1 U6557 ( .ip1(n8680), .ip2(n8679), .op(n5544) );
  ab_or_c_or_d U6558 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[1]), 
        .ip2(n8230), .ip3(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[0]), .ip4(
        n8229), .op(n5549) );
  or2_1 U6559 ( .ip1(n8230), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[1]), 
        .op(n5550) );
  inv_1 U6560 ( .ip(n8225), .op(n8236) );
  inv_1 U6561 ( .ip(n5554), .op(n8273) );
  inv_1 U6562 ( .ip(n8214), .op(n5553) );
  mux2_2 U6563 ( .ip1(i_i2c_ic_fs_hcnt[8]), .ip2(i_i2c_ic_hcnt[8]), .s(n5458), 
        .op(n8258) );
  inv_1 U6564 ( .ip(n8275), .op(n5558) );
  nand2_1 U6565 ( .ip1(n8242), .ip2(n8241), .op(n8250) );
  nand2_1 U6566 ( .ip1(n8257), .ip2(n8256), .op(n5559) );
  nor2_1 U6567 ( .ip1(n8272), .ip2(n8283), .op(n8286) );
  inv_1 U6568 ( .ip(n9398), .op(n5556) );
  nand3_1 U6569 ( .ip1(n9405), .ip2(n9404), .ip3(n9403), .op(n5557) );
  or2_1 U6570 ( .ip1(n9232), .ip2(n9192), .op(n9193) );
  nor2_2 U6571 ( .ip1(n9331), .ip2(n8710), .op(n5153) );
  nand2_1 U6572 ( .ip1(n6043), .ip2(i_i2c_ic_fs_hcnt[1]), .op(n6066) );
  nand2_1 U6573 ( .ip1(n8208), .ip2(n6129), .op(n8209) );
  nand2_1 U6574 ( .ip1(n8273), .ip2(n8274), .op(n5560) );
  nor2_1 U6575 ( .ip1(n8761), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[10]), .op(n8630) );
  buf_4 U6576 ( .ip(n6060), .op(n6041) );
  or2_1 U6577 ( .ip1(n8229), .ip2(n8227), .op(n5561) );
  inv_1 U6578 ( .ip(n9521), .op(n5562) );
  or2_1 U6579 ( .ip1(n8285), .ip2(n8286), .op(n8287) );
  xor2_2 U6580 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[0]), .ip2(n8519), 
        .op(n8491) );
  nor2_4 U6581 ( .ip1(n8388), .ip2(n8362), .op(n5140) );
  or2_1 U6582 ( .ip1(n9189), .ip2(n9188), .op(n5563) );
  nand2_2 U6583 ( .ip1(n9166), .ip2(n9235), .op(n9228) );
  or2_1 U6584 ( .ip1(n9175), .ip2(n9186), .op(n5564) );
  or2_1 U6585 ( .ip1(n9175), .ip2(n9186), .op(n9176) );
  xnor2_2 U6586 ( .ip1(i_i2c_ic_sda_tx_hold_sync[9]), .ip2(n5565), .op(n9383)
         );
  or2_1 U6587 ( .ip1(n9214), .ip2(n9282), .op(n5565) );
  and2_2 U6588 ( .ip1(n5258), .ip2(n9191), .op(n9232) );
  nand2_1 U6589 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[12]), 
        .ip2(n5582), .op(n9407) );
  xnor2_2 U6590 ( .ip1(i_i2c_ic_sda_tx_hold_sync[3]), .ip2(n9174), .op(n9188)
         );
  xnor2_1 U6591 ( .ip1(i_i2c_ic_sda_tx_hold_sync[2]), .ip2(n9176), .op(n5566)
         );
  inv_1 U6592 ( .ip(n9414), .op(n9419) );
  inv_1 U6593 ( .ip(n9169), .op(n5586) );
  or2_1 U6594 ( .ip1(n9198), .ip2(n9282), .op(n5568) );
  nand2_1 U6595 ( .ip1(n5569), .ip2(n9395), .op(n9413) );
  nor2_1 U6596 ( .ip1(n5571), .ip2(n9458), .op(n9462) );
  nand2_1 U6597 ( .ip1(n5570), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[11]), .op(n5571) );
  mux2_1 U6598 ( .ip1(i_i2c_ic_fs_spklen[1]), .ip2(i_i2c_ic_hs_spklen[1]), .s(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r), .op(n5572) );
  and2_1 U6599 ( .ip1(n9106), .ip2(i_i2c_ic_sda_tx_hold_sync[2]), .op(n9110)
         );
  nand2_1 U6600 ( .ip1(n5573), .ip2(n5574), .op(n5576) );
  or2_1 U6601 ( .ip1(n9138), .ip2(n5577), .op(n5575) );
  nand2_1 U6602 ( .ip1(n5575), .ip2(n5576), .op(n9104) );
  or2_1 U6603 ( .ip1(n9149), .ip2(i_i2c_ic_sda_tx_hold_sync[6]), .op(n5577) );
  and2_1 U6604 ( .ip1(n5578), .ip2(n9392), .op(n5585) );
  nand2_1 U6605 ( .ip1(n5517), .ip2(n5581), .op(n5578) );
  or2_1 U6606 ( .ip1(n9210), .ip2(n9282), .op(n5580) );
  inv_1 U6607 ( .ip(n9384), .op(n9390) );
  inv_1 U6608 ( .ip(n5582), .op(n9415) );
  nand2_1 U6609 ( .ip1(n9391), .ip2(n5585), .op(n9395) );
  nor2_1 U6610 ( .ip1(n9244), .ip2(n9246), .op(n9190) );
  nor2_1 U6611 ( .ip1(n9232), .ip2(n9226), .op(n9227) );
  nand2_1 U6612 ( .ip1(n9228), .ip2(n9173), .op(n5587) );
  xor2_2 U6613 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[0]), .ip2(n5476), .op(n8305) );
  and2_1 U6614 ( .ip1(n9375), .ip2(n9431), .op(n9372) );
  or2_1 U6615 ( .ip1(n5557), .ip2(n9410), .op(n9414) );
  nand2_1 U6616 ( .ip1(i_ssi_tx_pop_sync), .ip2(i_ssi_U_fifo_U_tx_fifo_empty_n), .op(n5588) );
  and2_4 U6617 ( .ip1(n10776), .ip2(i_ssi_rx_wr_addr[2]), .op(n10777) );
  nand2_2 U6618 ( .ip1(n10228), .ip2(n10223), .op(n10365) );
  and2_1 U6619 ( .ip1(n8252), .ip2(n8253), .op(n5589) );
  nor2_2 U6620 ( .ip1(n9685), .ip2(n11117), .op(n5592) );
  and2_1 U6621 ( .ip1(n6305), .ip2(n7753), .op(n5593) );
  and2_1 U6622 ( .ip1(n5553), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[5]), .op(n5595) );
  and2_1 U6623 ( .ip1(n8254), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[7]), .op(n5596) );
  xnor2_2 U6624 ( .ip1(n6176), .ip2(n6175), .op(n5598) );
  or2_1 U6625 ( .ip1(n8258), .ip2(n6125), .op(n5599) );
  nand2_1 U6626 ( .ip1(n6237), .ip2(n6236), .op(n5600) );
  and2_1 U6627 ( .ip1(n9098), .ip2(n9097), .op(n5604) );
  xor2_1 U6628 ( .ip1(n7355), .ip2(n7354), .op(n5606) );
  inv_2 U6629 ( .ip(i_ssi_load_start_bit), .op(n10416) );
  xnor2_2 U6630 ( .ip1(i_ssi_U_mstfsm_frame_cnt[10]), .ip2(n9890), .op(n5607)
         );
  nor2_4 U6631 ( .ip1(n10220), .ip2(n10203), .op(n5608) );
  and2_4 U6632 ( .ip1(n10776), .ip2(n10779), .op(n10721) );
  nor2_2 U6633 ( .ip1(n10243), .ip2(n10244), .op(n5609) );
  nor2_2 U6634 ( .ip1(n10784), .ip2(n10781), .op(n5610) );
  nor2_2 U6635 ( .ip1(n10782), .ip2(n10781), .op(n5611) );
  and4_1 U6636 ( .ip1(n6418), .ip2(n10802), .ip3(n11004), .ip4(n7394), .op(
        n5612) );
  nand2_1 U6637 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[9]), .ip2(n7753), .op(n7758) );
  or2_1 U6638 ( .ip1(n6029), .ip2(n11152), .op(n5613) );
  inv_1 U6639 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[3]), .op(n8224)
         );
  xor2_1 U6640 ( .ip1(i_ssi_rx_rd_addr[2]), .ip2(n10131), .op(n5614) );
  and2_1 U6641 ( .ip1(n7757), .ip2(n6277), .op(n5615) );
  inv_1 U6642 ( .ip(i_ahb_U_dfltslv_current_state), .op(n6677) );
  inv_1 U6643 ( .ip(i_ssi_U_sclkgen_ssi_cnt[4]), .op(n6422) );
  and2_1 U6644 ( .ip1(i_ssi_U_mstfsm_frame_cnt[12]), .ip2(
        i_ssi_U_mstfsm_frame_cnt[13]), .op(n5619) );
  nand2_1 U6645 ( .ip1(i_ssi_U_mstfsm_frame_cnt[11]), .ip2(
        i_ssi_U_mstfsm_frame_cnt[10]), .op(n6033) );
  inv_1 U6646 ( .ip(n6033), .op(n5618) );
  nand2_1 U6647 ( .ip1(n5619), .ip2(n5618), .op(n7164) );
  and2_1 U6648 ( .ip1(i_ssi_U_mstfsm_bit_cnt[3]), .ip2(
        i_ssi_U_mstfsm_bit_cnt[4]), .op(n5621) );
  inv_1 U6649 ( .ip(i_ssi_U_mstfsm_bit_cnt[3]), .op(n9838) );
  nor2_1 U6650 ( .ip1(n9838), .ip2(i_ssi_dfs[3]), .op(n5620) );
  nor2_1 U6651 ( .ip1(i_ssi_U_mstfsm_bit_cnt[4]), .ip2(n5620), .op(n5626) );
  nor2_1 U6652 ( .ip1(i_ssi_dfs[2]), .ip2(i_ssi_dfs[3]), .op(n10843) );
  inv_1 U6653 ( .ip(i_ssi_U_mstfsm_bit_cnt[1]), .op(n9827) );
  nor2_1 U6654 ( .ip1(i_ssi_U_mstfsm_bit_cnt[3]), .ip2(n9827), .op(n5622) );
  nand2_1 U6655 ( .ip1(n10843), .ip2(n5622), .op(n5623) );
  nand2_1 U6656 ( .ip1(n5623), .ip2(n5760), .op(n5624) );
  inv_1 U6657 ( .ip(i_ssi_U_mstfsm_c_state[3]), .op(n9974) );
  nand2_1 U6658 ( .ip1(n9974), .ip2(i_ssi_U_mstfsm_c_state[2]), .op(n5733) );
  nor2_1 U6659 ( .ip1(i_ssi_U_mstfsm_c_state[0]), .ip2(n5733), .op(n10699) );
  inv_1 U6660 ( .ip(i_ssi_U_mstfsm_c_state[1]), .op(n10111) );
  nand2_1 U6661 ( .ip1(n10111), .ip2(i_ssi_sclk_fe), .op(n10112) );
  inv_1 U6662 ( .ip(n10112), .op(n9975) );
  nand2_1 U6663 ( .ip1(n10699), .ip2(n9975), .op(n10430) );
  and2_1 U6664 ( .ip1(i_ssi_U_mstfsm_bit_cnt[2]), .ip2(
        i_ssi_U_mstfsm_bit_cnt[1]), .op(n5627) );
  inv_1 U6665 ( .ip(n5627), .op(n5634) );
  nand2_1 U6666 ( .ip1(n9838), .ip2(n5327), .op(n5625) );
  nand2_1 U6667 ( .ip1(n5626), .ip2(n5625), .op(n5768) );
  nand2_1 U6668 ( .ip1(n5627), .ip2(n5353), .op(n5629) );
  nand2_1 U6669 ( .ip1(n10737), .ip2(n9827), .op(n5628) );
  nand2_1 U6670 ( .ip1(n5629), .ip2(n5628), .op(n5633) );
  inv_1 U6671 ( .ip(i_ssi_dfs[2]), .op(n10743) );
  nand4_1 U6672 ( .ip1(n10743), .ip2(i_ssi_U_mstfsm_bit_cnt[3]), .ip3(n5327), 
        .ip4(i_ssi_U_mstfsm_bit_cnt[1]), .op(n5631) );
  nand3_1 U6673 ( .ip1(n5272), .ip2(i_ssi_tmod[0]), .ip3(
        i_ssi_U_mstfsm_spi0_control), .op(n5630) );
  nand2_1 U6674 ( .ip1(n5631), .ip2(n5630), .op(n5632) );
  not_ab_or_c_or_d U6675 ( .ip1(n5634), .ip2(n5768), .ip3(n5633), .ip4(n5632), 
        .op(n5635) );
  inv_1 U6676 ( .ip(i_ssi_U_mstfsm_frame_cnt[2]), .op(n5651) );
  nand2_1 U6677 ( .ip1(i_ssi_U_mstfsm_frame_cnt[1]), .ip2(
        i_ssi_U_mstfsm_frame_cnt[0]), .op(n9865) );
  nor2_1 U6678 ( .ip1(n5651), .ip2(n9865), .op(n9875) );
  and2_1 U6679 ( .ip1(i_ssi_U_mstfsm_frame_cnt[4]), .ip2(
        i_ssi_U_mstfsm_frame_cnt[3]), .op(n5637) );
  nand2_1 U6680 ( .ip1(n9875), .ip2(n5637), .op(n9874) );
  and2_1 U6681 ( .ip1(i_ssi_U_mstfsm_frame_cnt[5]), .ip2(
        i_ssi_U_mstfsm_frame_cnt[6]), .op(n9886) );
  nand2_1 U6682 ( .ip1(i_ssi_U_mstfsm_frame_cnt[8]), .ip2(
        i_ssi_U_mstfsm_frame_cnt[7]), .op(n5638) );
  inv_1 U6685 ( .ip(i_ssi_U_mstfsm_frame_cnt[13]), .op(n9897) );
  nand2_1 U6686 ( .ip1(n9897), .ip2(i_ssi_U_regfile_ctrlr1_int[13]), .op(n5640) );
  xor2_1 U6687 ( .ip1(i_ssi_U_mstfsm_frame_cnt[14]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[14]), .op(n5639) );
  nand2_1 U6688 ( .ip1(n5390), .ip2(i_ssi_U_regfile_ctrlr1_int[11]), .op(n5642) );
  xor2_1 U6689 ( .ip1(i_ssi_U_mstfsm_frame_cnt[12]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[12]), .op(n5641) );
  inv_1 U6690 ( .ip(i_ssi_U_mstfsm_frame_cnt[12]), .op(n6034) );
  nand2_1 U6691 ( .ip1(n6034), .ip2(i_ssi_U_regfile_ctrlr1_int[12]), .op(n5644) );
  xor2_1 U6692 ( .ip1(i_ssi_U_regfile_ctrlr1_int[13]), .ip2(
        i_ssi_U_mstfsm_frame_cnt[13]), .op(n5643) );
  xnor2_1 U6693 ( .ip1(n5644), .ip2(n5643), .op(n5648) );
  inv_1 U6694 ( .ip(i_ssi_U_mstfsm_frame_cnt[14]), .op(n7165) );
  nand2_1 U6695 ( .ip1(n7165), .ip2(i_ssi_U_regfile_ctrlr1_int[14]), .op(n5646) );
  nand2_1 U6696 ( .ip1(n5651), .ip2(i_ssi_U_regfile_ctrlr1_int[2]), .op(n5667)
         );
  inv_1 U6697 ( .ip(i_ssi_U_regfile_ctrlr1_int[2]), .op(n5652) );
  nand2_1 U6698 ( .ip1(n5652), .ip2(i_ssi_U_mstfsm_frame_cnt[2]), .op(n5675)
         );
  nand2_1 U6699 ( .ip1(n5667), .ip2(n5675), .op(n5654) );
  inv_1 U6700 ( .ip(i_ssi_U_mstfsm_frame_cnt[1]), .op(n5653) );
  nand2_1 U6701 ( .ip1(n5653), .ip2(i_ssi_U_regfile_ctrlr1_int[1]), .op(n5669)
         );
  nand2_1 U6702 ( .ip1(n5654), .ip2(n5669), .op(n5657) );
  xor2_1 U6703 ( .ip1(i_ssi_U_mstfsm_frame_cnt[1]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[0]), .op(n5655) );
  xnor2_1 U6704 ( .ip1(i_ssi_U_regfile_ctrlr1_int[1]), .ip2(n5655), .op(n5656)
         );
  nand2_1 U6705 ( .ip1(n5657), .ip2(n5656), .op(n5666) );
  inv_1 U6706 ( .ip(i_ssi_U_mstfsm_frame_cnt[4]), .op(n5660) );
  nand2_1 U6707 ( .ip1(n5660), .ip2(i_ssi_U_regfile_ctrlr1_int[4]), .op(n5662)
         );
  xor2_1 U6708 ( .ip1(i_ssi_U_mstfsm_frame_cnt[5]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[5]), .op(n5661) );
  xnor2_1 U6709 ( .ip1(n5662), .ip2(n5661), .op(n5663) );
  inv_1 U6710 ( .ip(n5663), .op(n5664) );
  nand2_1 U6711 ( .ip1(n5659), .ip2(n5664), .op(n5665) );
  inv_1 U6712 ( .ip(n5667), .op(n5668) );
  nor2_1 U6713 ( .ip1(n5669), .ip2(n5668), .op(n5674) );
  inv_1 U6714 ( .ip(i_ssi_U_mstfsm_frame_cnt[3]), .op(n9869) );
  nand2_1 U6715 ( .ip1(n9869), .ip2(i_ssi_U_regfile_ctrlr1_int[3]), .op(n5671)
         );
  xor2_1 U6716 ( .ip1(i_ssi_U_regfile_ctrlr1_int[4]), .ip2(
        i_ssi_U_mstfsm_frame_cnt[4]), .op(n5670) );
  xnor2_1 U6717 ( .ip1(n5671), .ip2(n5670), .op(n5673) );
  xnor2_1 U6718 ( .ip1(i_ssi_U_mstfsm_frame_cnt[0]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[0]), .op(n5672) );
  not_ab_or_c_or_d U6719 ( .ip1(n5675), .ip2(n5674), .ip3(n5673), .ip4(n5672), 
        .op(n5676) );
  nand2_1 U6720 ( .ip1(n5677), .ip2(n5676), .op(n10417) );
  nor2_1 U6721 ( .ip1(n9848), .ip2(n5396), .op(n5799) );
  inv_1 U6722 ( .ip(i_ssi_U_mstfsm_frame_cnt[5]), .op(n5678) );
  nand2_1 U6723 ( .ip1(n5678), .ip2(i_ssi_U_regfile_ctrlr1_int[5]), .op(n5680)
         );
  inv_1 U6724 ( .ip(i_ssi_U_mstfsm_frame_cnt[8]), .op(n9888) );
  nand2_1 U6725 ( .ip1(n9888), .ip2(i_ssi_U_regfile_ctrlr1_int[8]), .op(n5682)
         );
  inv_1 U6726 ( .ip(i_ssi_U_mstfsm_frame_cnt[7]), .op(n5683) );
  nand2_1 U6727 ( .ip1(n5683), .ip2(i_ssi_U_regfile_ctrlr1_int[7]), .op(n5685)
         );
  xnor2_1 U6728 ( .ip1(n5685), .ip2(n5684), .op(n5690) );
  inv_1 U6729 ( .ip(i_ssi_U_mstfsm_frame_cnt[6]), .op(n5686) );
  nand2_1 U6730 ( .ip1(n5686), .ip2(i_ssi_U_regfile_ctrlr1_int[6]), .op(n5688)
         );
  xnor2_1 U6731 ( .ip1(n5688), .ip2(n5687), .op(n5689) );
  nor4_2 U6732 ( .ip1(n5692), .ip2(n5690), .ip3(n5691), .ip4(n5689), .op(n5802) );
  nand2_1 U6733 ( .ip1(n5425), .ip2(i_ssi_U_mstfsm_c_state[3]), .op(n5712) );
  inv_1 U6734 ( .ip(n5712), .op(n5693) );
  inv_1 U6735 ( .ip(i_ssi_U_mstfsm_frame_cnt[15]), .op(n9902) );
  xor2_1 U6736 ( .ip1(i_ssi_U_mstfsm_frame_cnt[16]), .ip2(n5709), .op(n9847)
         );
  and4_1 U6737 ( .ip1(n10111), .ip2(n5693), .ip3(n5272), .ip4(n9847), .op(
        n5704) );
  inv_1 U6738 ( .ip(i_ssi_U_mstfsm_frame_cnt[10]), .op(n5694) );
  nand2_1 U6739 ( .ip1(n5694), .ip2(i_ssi_U_regfile_ctrlr1_int[10]), .op(n5696) );
  xnor2_1 U6740 ( .ip1(n5696), .ip2(n5695), .op(n5697) );
  inv_1 U6741 ( .ip(n5697), .op(n5702) );
  inv_1 U6742 ( .ip(i_ssi_U_mstfsm_frame_cnt[9]), .op(n9892) );
  nand2_1 U6743 ( .ip1(i_ssi_U_regfile_ctrlr1_int[9]), .ip2(n9892), .op(n5699)
         );
  xnor2_1 U6744 ( .ip1(n5699), .ip2(n5698), .op(n5700) );
  inv_1 U6745 ( .ip(n5700), .op(n5701) );
  inv_1 U6746 ( .ip(n5800), .op(n5703) );
  nand2_1 U6747 ( .ip1(n5704), .ip2(n5703), .op(n5705) );
  nor2_1 U6748 ( .ip1(n5439), .ip2(n5705), .op(n5706) );
  nand2_1 U6749 ( .ip1(n5799), .ip2(n5706), .op(n5795) );
  inv_1 U6750 ( .ip(n5795), .op(n5792) );
  inv_1 U6751 ( .ip(i_ssi_mwcr[1]), .op(n5741) );
  nand2_1 U6752 ( .ip1(n5502), .ip2(n5741), .op(n5708) );
  nand2_1 U6753 ( .ip1(n9974), .ip2(i_ssi_U_mstfsm_c_state[1]), .op(n5707) );
  nand2_1 U6754 ( .ip1(n5425), .ip2(i_ssi_U_mstfsm_c_state[0]), .op(n9973) );
  nor2_1 U6755 ( .ip1(n5707), .ip2(n9973), .op(n9972) );
  nand2_1 U6756 ( .ip1(n9972), .ip2(i_ssi_U_mstfsm_c_done_ir), .op(n5747) );
  inv_1 U6757 ( .ip(i_ssi_U_mstfsm_frame_cnt[16]), .op(n5710) );
  nor2_1 U6758 ( .ip1(n5711), .ip2(n10429), .op(n5713) );
  or2_1 U6759 ( .ip1(i_ssi_U_mstfsm_c_state[1]), .ip2(
        i_ssi_U_mstfsm_c_state[0]), .op(n5725) );
  nor2_1 U6760 ( .ip1(n5712), .ip2(n5725), .op(n5804) );
  nand3_1 U6761 ( .ip1(n5799), .ip2(n5745), .ip3(n5714), .op(n5717) );
  nand2_1 U6762 ( .ip1(n5745), .ip2(n5715), .op(n5716) );
  nand2_1 U6763 ( .ip1(n5716), .ip2(n5717), .op(n5797) );
  nor2_1 U6764 ( .ip1(i_ssi_U_mstfsm_c_state[0]), .ip2(n10111), .op(n5721) );
  nor3_1 U6765 ( .ip1(i_ssi_U_mstfsm_c_state[1]), .ip2(n5498), .ip3(n9973), 
        .op(n5720) );
  and2_1 U6766 ( .ip1(i_ssi_U_mstfsm_c_state[3]), .ip2(
        i_ssi_U_mstfsm_c_state[2]), .op(n5729) );
  not_ab_or_c_or_d U6767 ( .ip1(n5290), .ip2(i_ssi_sclk_re), .ip3(n5718), 
        .ip4(n5750), .op(n5719) );
  not_ab_or_c_or_d U6768 ( .ip1(n5400), .ip2(n5721), .ip3(n5720), .ip4(n5719), 
        .op(n5722) );
  nand2_1 U6769 ( .ip1(n10111), .ip2(i_ssi_U_mstfsm_c_state[3]), .op(n5730) );
  inv_1 U6770 ( .ip(n5777), .op(n5723) );
  inv_1 U6771 ( .ip(n5725), .op(n9802) );
  nand2_1 U6772 ( .ip1(n5729), .ip2(n9802), .op(n9853) );
  nor2_1 U6773 ( .ip1(i_ssi_U_mstfsm_c_state[2]), .ip2(
        i_ssi_U_mstfsm_c_state[0]), .op(n5753) );
  and2_1 U6774 ( .ip1(i_ssi_U_mstfsm_c_state[3]), .ip2(
        i_ssi_U_mstfsm_c_state[1]), .op(n5726) );
  nand2_1 U6775 ( .ip1(n5753), .ip2(n5726), .op(n6031) );
  inv_1 U6776 ( .ip(i_ssi_U_mstfsm_c_state[0]), .op(n9812) );
  nor2_1 U6777 ( .ip1(i_ssi_U_mstfsm_c_state[1]), .ip2(n9812), .op(n5728) );
  nand2_1 U6778 ( .ip1(n5729), .ip2(n5728), .op(n10231) );
  inv_1 U6779 ( .ip(n10231), .op(n10966) );
  nand2_1 U6780 ( .ip1(n5425), .ip2(i_ssi_U_mstfsm_abort_ir), .op(n5731) );
  nand2_1 U6781 ( .ip1(n9973), .ip2(n5731), .op(n5732) );
  nand2_1 U6782 ( .ip1(n5732), .ip2(n5289), .op(n5736) );
  inv_1 U6783 ( .ip(i_ssi_sclk_fe), .op(n10421) );
  nor2_1 U6784 ( .ip1(n9812), .ip2(n5733), .op(n10114) );
  nand2_1 U6785 ( .ip1(n10114), .ip2(i_ssi_U_mstfsm_c_state[1]), .op(n9907) );
  or2_1 U6786 ( .ip1(n10421), .ip2(n9907), .op(n5735) );
  nand2_1 U6787 ( .ip1(n5290), .ip2(i_ssi_U_mstfsm_c_done_ir), .op(n5742) );
  nand2_1 U6788 ( .ip1(n10114), .ip2(n10111), .op(n10701) );
  nor2_1 U6789 ( .ip1(n10966), .ip2(n10699), .op(n5746) );
  nand2_1 U6790 ( .ip1(n5338), .ip2(n5746), .op(n5752) );
  inv_1 U6791 ( .ip(n5747), .op(n5749) );
  nand2_1 U6792 ( .ip1(n5749), .ip2(n5748), .op(n5751) );
  nand2_1 U6793 ( .ip1(n5753), .ip2(n9974), .op(n9797) );
  nor2_1 U6794 ( .ip1(n10111), .ip2(n9797), .op(n10418) );
  nand2_1 U6795 ( .ip1(n5781), .ip2(n10699), .op(n5771) );
  inv_1 U6796 ( .ip(n9973), .op(n5769) );
  nand2_1 U6797 ( .ip1(n5769), .ip2(n5498), .op(n5770) );
  nand2_1 U6798 ( .ip1(n5771), .ip2(n5770), .op(n5785) );
  inv_1 U6799 ( .ip(i_ssi_U_mstfsm_ss_in_n_sync), .op(n9988) );
  nor4_1 U6800 ( .ip1(i_ssi_mst_contention), .ip2(n5492), .ip3(n9988), .ip4(
        n10112), .op(n5772) );
  inv_1 U6801 ( .ip(n9797), .op(n9817) );
  nand2_1 U6802 ( .ip1(n5772), .ip2(n9817), .op(n5773) );
  nand2_1 U6803 ( .ip1(n5338), .ip2(n5773), .op(n5784) );
  nor2_1 U6804 ( .ip1(n5492), .ip2(n5498), .op(n5774) );
  mux2_1 U6805 ( .ip1(n5501), .ip2(n5774), .s(i_ssi_mwcr[1]), .op(n5775) );
  nand2_1 U6806 ( .ip1(n5775), .ip2(i_ssi_U_mstfsm_c_done_ir), .op(n5778) );
  not_ab_or_c_or_d U6807 ( .ip1(n9972), .ip2(n5778), .ip3(n5777), .ip4(n5776), 
        .op(n5783) );
  inv_1 U6808 ( .ip(i_ssi_mwcr[0]), .op(n5786) );
  nand2_1 U6809 ( .ip1(n5502), .ip2(n5786), .op(n5779) );
  nor2_1 U6810 ( .ip1(n5779), .ip2(n9853), .op(n5780) );
  nand2_1 U6811 ( .ip1(n5781), .ip2(n5780), .op(n5782) );
  nand2_1 U6812 ( .ip1(n5783), .ip2(n5782), .op(n5808) );
  not_ab_or_c_or_d U6813 ( .ip1(n10111), .ip2(n5785), .ip3(n5784), .ip4(n5808), 
        .op(n5791) );
  nand2_1 U6814 ( .ip1(n5786), .ip2(n5290), .op(n10230) );
  nand2_1 U6815 ( .ip1(n9815), .ip2(n10230), .op(n5810) );
  inv_1 U6816 ( .ip(i_ssi_sclk_re), .op(n5787) );
  nand2_1 U6817 ( .ip1(n5810), .ip2(n5787), .op(n5788) );
  nand2_1 U6818 ( .ip1(i_ssi_rxd), .ip2(n5788), .op(n5789) );
  nand2_1 U6819 ( .ip1(n10966), .ip2(n5789), .op(n5790) );
  and2_1 U6820 ( .ip1(n5791), .ip2(n5790), .op(n10982) );
  inv_1 U6821 ( .ip(n10982), .op(n10988) );
  inv_1 U6822 ( .ip(n5405), .op(n5794) );
  and2_1 U6823 ( .ip1(n5795), .ip2(n5794), .op(n9989) );
  nand2_1 U6824 ( .ip1(n5797), .ip2(n5452), .op(n10981) );
  nor2_1 U6825 ( .ip1(n9989), .ip2(n10981), .op(n5815) );
  inv_1 U6826 ( .ip(n5798), .op(n5806) );
  nand2_1 U6827 ( .ip1(n5799), .ip2(n9847), .op(n9904) );
  inv_1 U6828 ( .ip(n9904), .op(n5803) );
  nand2_1 U6829 ( .ip1(n5802), .ip2(n5801), .op(n9846) );
  nand2_1 U6830 ( .ip1(n5803), .ip2(n5370), .op(n5805) );
  inv_1 U6831 ( .ip(n5804), .op(n9807) );
  not_ab_or_c_or_d U6832 ( .ip1(n5806), .ip2(n5805), .ip3(n5400), .ip4(n9807), 
        .op(n5807) );
  ab_or_c_or_d U6833 ( .ip1(n5809), .ip2(i_ssi_sclk_re), .ip3(n5808), .ip4(
        n5807), .op(n7319) );
  nor2_1 U6834 ( .ip1(n10231), .ip2(n5810), .op(n5811) );
  nand2_1 U6835 ( .ip1(i_ssi_rxd), .ip2(n5811), .op(n5812) );
  nand2_1 U6836 ( .ip1(n5815), .ip2(n10987), .op(n5816) );
  nand2_1 U6837 ( .ip1(n5355), .ip2(n5816), .op(n10952) );
  inv_1 U6838 ( .ip(n10952), .op(n11794) );
  inv_1 U6871 ( .ip(HRESETn_hresetn), .op(n11829) );
  inv_1 U6872 ( .ip(i_i2c_mst_debug_cstate[3]), .op(n5844) );
  and2_1 U6873 ( .ip1(n7873), .ip2(n7685), .op(n10926) );
  or2_1 U6874 ( .ip1(i_i2c_scl_hcnt_en), .ip2(i_i2c_rx_scl_hcnt_en), .op(n8330) );
  nand2_1 U6875 ( .ip1(n8330), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_int_d), 
        .op(n6353) );
  xor2_1 U6876 ( .ip1(i_i2c_ic_fs_spklen[6]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[6]), .op(n5820) );
  xor2_1 U6877 ( .ip1(i_i2c_ic_fs_spklen[0]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[0]), .op(n5819) );
  xor2_1 U6878 ( .ip1(i_i2c_ic_fs_spklen[4]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[4]), .op(n5818) );
  xor2_1 U6879 ( .ip1(i_i2c_ic_fs_spklen[3]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[3]), .op(n5817) );
  nor4_2 U6880 ( .ip1(n5820), .ip2(n5819), .ip3(n5818), .ip4(n5817), .op(n5827) );
  inv_1 U6881 ( .ip(i_i2c_ic_fs_spklen[7]), .op(n5861) );
  and2_1 U6882 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[7]), 
        .ip2(n5861), .op(n7454) );
  nor2_1 U6883 ( .ip1(n5861), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[7]), .op(n7457) );
  inv_1 U6884 ( .ip(i_i2c_ic_fs_sync), .op(n8072) );
  and3_1 U6885 ( .ip1(n8072), .ip2(i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r), 
        .ip3(n5851), .op(n5862) );
  inv_1 U6886 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[1]), .op(
        n5823) );
  nand2_1 U6887 ( .ip1(n5823), .ip2(i_i2c_ic_fs_spklen[1]), .op(n7443) );
  inv_1 U6888 ( .ip(i_i2c_ic_fs_spklen[1]), .op(n6067) );
  nand2_1 U6889 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[1]), 
        .ip2(n6067), .op(n7439) );
  nand2_1 U6890 ( .ip1(n7443), .ip2(n7439), .op(n5824) );
  nand3_1 U6891 ( .ip1(n5826), .ip2(n5827), .ip3(n5825), .op(n5839) );
  xor2_1 U6892 ( .ip1(i_i2c_ic_hs_spklen[4]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[4]), .op(n5831) );
  xor2_1 U6893 ( .ip1(i_i2c_ic_hs_spklen[0]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[0]), .op(n5829) );
  xor2_1 U6894 ( .ip1(i_i2c_ic_hs_spklen[3]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[3]), .op(n5832) );
  inv_1 U6895 ( .ip(i_i2c_ic_hs_spklen[1]), .op(n5881) );
  nor2_1 U6896 ( .ip1(n5881), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[1]), .op(n7466) );
  and2_1 U6897 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[1]), 
        .ip2(n5881), .op(n7469) );
  nor3_1 U6898 ( .ip1(n5832), .ip2(n7466), .ip3(n7469), .op(n5836) );
  xor2_1 U6899 ( .ip1(i_i2c_ic_hs_spklen[2]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[2]), .op(n5834) );
  inv_1 U6900 ( .ip(i_i2c_ic_hs_spklen[7]), .op(n5887) );
  nor2_1 U6901 ( .ip1(n5887), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[7]), .op(n7484) );
  nand2_1 U6902 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[7]), 
        .ip2(n5887), .op(n5833) );
  nand2_1 U6903 ( .ip1(n5833), .ip2(i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r), 
        .op(n7488) );
  nor3_1 U6904 ( .ip1(n5834), .ip2(n7484), .ip3(n7488), .op(n5835) );
  nand3_1 U6905 ( .ip1(n5837), .ip2(n5836), .ip3(n5835), .op(n5838) );
  nand2_1 U6906 ( .ip1(n5839), .ip2(n5838), .op(n5840) );
  inv_1 U6907 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_data_d_int_0_), 
        .op(n9530) );
  nand2_1 U6908 ( .ip1(n5840), .ip2(n9530), .op(n5841) );
  nand2_1 U6909 ( .ip1(n7873), .ip2(i_i2c_mst_debug_cstate[0]), .op(n8332) );
  nor2_1 U6910 ( .ip1(n5844), .ip2(n8332), .op(n6359) );
  inv_1 U6911 ( .ip(i_i2c_U_DW_apb_i2c_mstfsm_N252), .op(n5845) );
  nor2_1 U6912 ( .ip1(i_i2c_ic_tar[10]), .ip2(n5845), .op(n7829) );
  nand2_1 U6913 ( .ip1(n6359), .ip2(n7829), .op(n5850) );
  inv_1 U6914 ( .ip(i_i2c_mst_debug_cstate[4]), .op(n7684) );
  nand2_1 U6915 ( .ip1(n5846), .ip2(n7684), .op(n6358) );
  nor2_1 U6916 ( .ip1(i_i2c_mst_debug_cstate[0]), .ip2(n6358), .op(n5848) );
  inv_1 U6917 ( .ip(n7685), .op(n5847) );
  nor2_1 U6918 ( .ip1(i_i2c_mst_debug_cstate[1]), .ip2(
        i_i2c_mst_debug_cstate[2]), .op(n6448) );
  nand2_1 U6919 ( .ip1(n6448), .ip2(n7684), .op(n7869) );
  nor2_1 U6920 ( .ip1(n5847), .ip2(n7869), .op(n7895) );
  nor2_1 U6921 ( .ip1(n5848), .ip2(n7895), .op(n5849) );
  nand2_1 U6922 ( .ip1(n5850), .ip2(n5849), .op(n5852) );
  nand2_1 U6923 ( .ip1(n5852), .ip2(n5851), .op(n5854) );
  nand2_1 U6924 ( .ip1(i_i2c_scl_lcnt_cmplt), .ip2(i_i2c_mst_tx_ack_vld), .op(
        n6355) );
  nand2_1 U6925 ( .ip1(n5854), .ip2(n5853), .op(n5855) );
  or4_1 U6926 ( .ip1(i_i2c_ic_sda_rx_hold_sync[3]), .ip2(
        i_i2c_ic_sda_rx_hold_sync[2]), .ip3(i_i2c_ic_sda_rx_hold_sync[1]), 
        .ip4(i_i2c_ic_sda_rx_hold_sync[0]), .op(n7611) );
  or2_1 U6927 ( .ip1(i_i2c_ic_sda_rx_hold_sync[4]), .ip2(n7611), .op(n7613) );
  or2_1 U6928 ( .ip1(i_i2c_ic_sda_rx_hold_sync[5]), .ip2(n7613), .op(n7599) );
  nor2_1 U6929 ( .ip1(i_i2c_ic_sda_rx_hold_sync[6]), .ip2(n7599), .op(n7601)
         );
  inv_1 U6930 ( .ip(i_i2c_ic_sda_rx_hold_sync[7]), .op(n7591) );
  nand2_1 U6931 ( .ip1(n7601), .ip2(n7591), .op(n7640) );
  inv_1 U6932 ( .ip(n5859), .op(n6352) );
  and2_1 U6933 ( .ip1(n7640), .ip2(n6352), .op(n5860) );
  inv_1 U6934 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_sda_post_hold_done), .op(
        n7644) );
  inv_1 U6935 ( .ip(n5860), .op(n5903) );
  inv_1 U6936 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_sda_data_int), .op(n5902) );
  nor2_1 U6937 ( .ip1(n5861), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[7]), .op(n7556) );
  and2_1 U6938 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[7]), 
        .ip2(n5861), .op(n7561) );
  xor2_1 U6939 ( .ip1(i_i2c_ic_fs_spklen[5]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[5]), .op(n5863) );
  inv_1 U6940 ( .ip(n5862), .op(n7460) );
  nor4_1 U6941 ( .ip1(n7556), .ip2(n7561), .ip3(n5863), .ip4(n7562), .op(n5873) );
  inv_1 U6942 ( .ip(i_i2c_ic_fs_spklen[0]), .op(n5866) );
  and2_1 U6943 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[1]), 
        .ip2(n6067), .op(n7537) );
  inv_1 U6944 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[1]), .op(
        n7568) );
  nand2_1 U6945 ( .ip1(n7568), .ip2(i_i2c_ic_fs_spklen[1]), .op(n5865) );
  inv_1 U6946 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[0]), .op(
        n7567) );
  nand2_1 U6947 ( .ip1(n7567), .ip2(i_i2c_ic_fs_spklen[0]), .op(n5864) );
  nand2_1 U6948 ( .ip1(n5865), .ip2(n5864), .op(n7540) );
  not_ab_or_c_or_d U6949 ( .ip1(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[0]), .ip2(n5866), .ip3(
        n7537), .ip4(n7540), .op(n5872) );
  inv_1 U6950 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[6]), .op(
        n7583) );
  nand2_1 U6951 ( .ip1(n7583), .ip2(i_i2c_ic_fs_spklen[6]), .op(n7555) );
  inv_1 U6952 ( .ip(i_i2c_ic_fs_spklen[2]), .op(n7440) );
  nand2_1 U6953 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[2]), 
        .ip2(n7440), .op(n7538) );
  inv_1 U6954 ( .ip(i_i2c_ic_fs_spklen[4]), .op(n9095) );
  nand2_1 U6955 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[4]), 
        .ip2(n9095), .op(n7551) );
  inv_1 U6956 ( .ip(i_i2c_ic_fs_spklen[6]), .op(n9093) );
  nand2_1 U6957 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[6]), 
        .ip2(n9093), .op(n7559) );
  and4_1 U6958 ( .ip1(n7555), .ip2(n7538), .ip3(n7551), .ip4(n7559), .op(n5871) );
  inv_1 U6959 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[4]), .op(
        n7577) );
  nand2_1 U6960 ( .ip1(n7577), .ip2(i_i2c_ic_fs_spklen[4]), .op(n7541) );
  inv_1 U6961 ( .ip(i_i2c_ic_fs_spklen[3]), .op(n7438) );
  nand2_1 U6962 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[3]), 
        .ip2(n7438), .op(n7542) );
  nand2_1 U6963 ( .ip1(n7541), .ip2(n7542), .op(n5869) );
  inv_1 U6964 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[2]), .op(
        n7571) );
  nand2_1 U6965 ( .ip1(n7571), .ip2(i_i2c_ic_fs_spklen[2]), .op(n5868) );
  inv_1 U6966 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[3]), .op(
        n7574) );
  nand2_1 U6967 ( .ip1(n7574), .ip2(i_i2c_ic_fs_spklen[3]), .op(n5867) );
  nand2_1 U6968 ( .ip1(n5868), .ip2(n5867), .op(n7543) );
  nor2_1 U6969 ( .ip1(n5869), .ip2(n7543), .op(n5870) );
  nand4_1 U6970 ( .ip1(n5873), .ip2(n5872), .ip3(n5871), .ip4(n5870), .op(
        n5895) );
  inv_1 U6971 ( .ip(i_i2c_ic_hs_spklen[3]), .op(n7462) );
  nand2_1 U6972 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[3]), 
        .ip2(n7462), .op(n7523) );
  inv_1 U6973 ( .ip(i_i2c_ic_hs_spklen[2]), .op(n7470) );
  nand2_1 U6974 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[2]), 
        .ip2(n7470), .op(n5874) );
  nand2_1 U6975 ( .ip1(n7523), .ip2(n5874), .op(n7519) );
  or2_1 U6976 ( .ip1(n5887), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[7]), .op(n7530) );
  inv_1 U6977 ( .ip(i_i2c_ic_hs_spklen[5]), .op(n7479) );
  nor2_1 U6978 ( .ip1(n7479), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[5]), .op(n5876) );
  inv_1 U6979 ( .ip(i_i2c_ic_hs_spklen[6]), .op(n9092) );
  nor2_1 U6980 ( .ip1(n9092), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[6]), .op(n5875) );
  nor2_1 U6981 ( .ip1(n5876), .ip2(n5875), .op(n5877) );
  nand2_1 U6982 ( .ip1(n7530), .ip2(n5877), .op(n7533) );
  nor2_1 U6983 ( .ip1(n7519), .ip2(n7533), .op(n5893) );
  inv_1 U6984 ( .ip(i_i2c_ic_hs_spklen[0]), .op(n7465) );
  inv_1 U6985 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r), .op(n5880) );
  nand2_1 U6986 ( .ip1(n7574), .ip2(i_i2c_ic_hs_spklen[3]), .op(n5879) );
  nand2_1 U6987 ( .ip1(n7571), .ip2(i_i2c_ic_hs_spklen[2]), .op(n5878) );
  nand2_1 U6988 ( .ip1(n5879), .ip2(n5878), .op(n7524) );
  not_ab_or_c_or_d U6989 ( .ip1(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[0]), .ip2(n7465), .ip3(
        n5880), .ip4(n7524), .op(n5892) );
  nand2_1 U6990 ( .ip1(n7577), .ip2(i_i2c_ic_hs_spklen[4]), .op(n7526) );
  nand2_1 U6991 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[1]), 
        .ip2(n5881), .op(n7520) );
  nand2_1 U6992 ( .ip1(n7526), .ip2(n7520), .op(n5884) );
  nand2_1 U6993 ( .ip1(n7568), .ip2(i_i2c_ic_hs_spklen[1]), .op(n5883) );
  nand2_1 U6994 ( .ip1(n7567), .ip2(i_i2c_ic_hs_spklen[0]), .op(n5882) );
  nand2_1 U6995 ( .ip1(n5883), .ip2(n5882), .op(n7521) );
  nor2_1 U6996 ( .ip1(n5884), .ip2(n7521), .op(n5891) );
  inv_1 U6997 ( .ip(i_i2c_ic_hs_spklen[4]), .op(n9094) );
  nand2_1 U6998 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[4]), 
        .ip2(n9094), .op(n5886) );
  nand2_1 U6999 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[5]), 
        .ip2(n7479), .op(n5885) );
  nand2_1 U7000 ( .ip1(n5886), .ip2(n5885), .op(n5890) );
  nand2_1 U7001 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[7]), 
        .ip2(n5887), .op(n5889) );
  nand2_1 U7002 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[6]), 
        .ip2(n9092), .op(n5888) );
  nand2_1 U7003 ( .ip1(n5889), .ip2(n5888), .op(n7531) );
  nor2_1 U7004 ( .ip1(n5890), .ip2(n7531), .op(n7528) );
  nand2_1 U7005 ( .ip1(n5895), .ip2(n5894), .op(n5900) );
  nor4_1 U7006 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[0]), 
        .ip2(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[3]), .ip3(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[1]), .ip4(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[7]), .op(n5897) );
  inv_1 U7007 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[2]), .op(
        n7504) );
  nor4_1 U7008 ( .ip1(n7501), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[4]), .ip3(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[5]), .ip4(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[6]), .op(n5896) );
  nand2_1 U7009 ( .ip1(n5897), .ip2(n5896), .op(n5899) );
  nor2_1 U7010 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_data_d_int_0_), 
        .ip2(n5472), .op(n5898) );
  nand2_1 U7011 ( .ip1(n5899), .ip2(n5898), .op(n7587) );
  nand2_1 U7012 ( .ip1(n5900), .ip2(n7587), .op(n5901) );
  mux2_1 U7013 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_data_d_int_0_), 
        .ip2(n5902), .s(n5901), .op(n7668) );
  nand2_1 U7014 ( .ip1(n5903), .ip2(n7668), .op(n5904) );
  and2_1 U7015 ( .ip1(n5905), .ip2(n5904), .op(n11833) );
  inv_1 U7016 ( .ip(i_i2c_s_det), .op(n9583) );
  inv_1 U7017 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[11]), .op(n6012)
         );
  nand2_1 U7018 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[10]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[9]), .op(n6011) );
  buf_1 U7019 ( .ip(i_i2c_ic_ss_sync), .op(n5908) );
  mux2_1 U7020 ( .ip1(i_i2c_ic_fs_lcnt[9]), .ip2(i_i2c_ic_lcnt[9]), .s(n5908), 
        .op(n5950) );
  mux2_1 U7021 ( .ip1(i_i2c_ic_fs_lcnt[5]), .ip2(i_i2c_ic_lcnt[5]), .s(n5908), 
        .op(n5920) );
  mux2_1 U7022 ( .ip1(i_i2c_ic_fs_lcnt[0]), .ip2(i_i2c_ic_lcnt[0]), .s(
        i_i2c_ic_ss_sync), .op(n5929) );
  mux2_1 U7023 ( .ip1(i_i2c_ic_fs_lcnt[1]), .ip2(i_i2c_ic_lcnt[1]), .s(
        i_i2c_ic_ss_sync), .op(n5928) );
  nand2_1 U7024 ( .ip1(n5929), .ip2(n5928), .op(n5906) );
  inv_1 U7025 ( .ip(n5906), .op(n5925) );
  mux2_1 U7026 ( .ip1(i_i2c_ic_fs_lcnt[2]), .ip2(i_i2c_ic_lcnt[2]), .s(n5907), 
        .op(n5926) );
  and2_1 U7027 ( .ip1(n5925), .ip2(n5926), .op(n5923) );
  mux2_1 U7028 ( .ip1(i_i2c_ic_fs_lcnt[3]), .ip2(i_i2c_ic_lcnt[3]), .s(n5908), 
        .op(n5924) );
  and2_1 U7029 ( .ip1(n5923), .ip2(n5924), .op(n5921) );
  mux2_1 U7030 ( .ip1(i_i2c_ic_fs_lcnt[4]), .ip2(i_i2c_ic_lcnt[4]), .s(n5907), 
        .op(n5922) );
  nand2_1 U7031 ( .ip1(n5921), .ip2(n5922), .op(n5909) );
  inv_1 U7032 ( .ip(n5909), .op(n5919) );
  inv_1 U7033 ( .ip(n5915), .op(n5910) );
  nor2_1 U7034 ( .ip1(n5913), .ip2(n5910), .op(n5911) );
  mux2_1 U7035 ( .ip1(i_i2c_ic_fs_lcnt[7]), .ip2(i_i2c_ic_lcnt[7]), .s(n5908), 
        .op(n5912) );
  nand2_1 U7036 ( .ip1(n5911), .ip2(n5912), .op(n5947) );
  inv_1 U7037 ( .ip(n5913), .op(n5914) );
  xor2_1 U7038 ( .ip1(n5915), .ip2(n5914), .op(n6476) );
  nor2_1 U7039 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[7]), .ip2(n5527), .op(n5917) );
  inv_1 U7040 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[6]), .op(n5916)
         );
  nand2_1 U7041 ( .ip1(n6476), .ip2(n5916), .op(n6472) );
  inv_1 U7042 ( .ip(n6472), .op(n5918) );
  nor2_1 U7043 ( .ip1(n5918), .ip2(n5917), .op(n5944) );
  xor2_1 U7044 ( .ip1(n5920), .ip2(n5919), .op(n6454) );
  inv_1 U7045 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[4]), .op(n5940)
         );
  xor2_1 U7046 ( .ip1(n5922), .ip2(n5921), .op(n6455) );
  nor3_1 U7047 ( .ip1(n5940), .ip2(n5939), .ip3(n6455), .op(n5942) );
  xor2_1 U7048 ( .ip1(n5924), .ip2(n5923), .op(n6466) );
  inv_1 U7049 ( .ip(n6466), .op(n5937) );
  xor2_1 U7050 ( .ip1(n5926), .ip2(n5925), .op(n6465) );
  inv_1 U7051 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[2]), .op(n5934)
         );
  and2_1 U7052 ( .ip1(n6465), .ip2(n5934), .op(n5933) );
  inv_1 U7053 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[3]), .op(n5927)
         );
  xor2_1 U7054 ( .ip1(n5928), .ip2(n5929), .op(n6458) );
  inv_1 U7055 ( .ip(n6458), .op(n5930) );
  inv_1 U7056 ( .ip(n5929), .op(n6457) );
  not_ab_or_c_or_d U7057 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[1]), 
        .ip2(n5930), .ip3(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[0]), .ip4(
        n5929), .op(n5932) );
  nor2_1 U7058 ( .ip1(n5930), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[1]), .op(n5931) );
  nor4_1 U7059 ( .ip1(n5933), .ip2(n5590), .ip3(n5932), .ip4(n5931), .op(n5936) );
  nor3_1 U7060 ( .ip1(n5934), .ip2(n5590), .ip3(n6465), .op(n5935) );
  not_ab_or_c_or_d U7061 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[3]), 
        .ip2(n5937), .ip3(n5936), .ip4(n5935), .op(n5938) );
  not_ab_or_c_or_d U7062 ( .ip1(n6455), .ip2(n5940), .ip3(n5939), .ip4(n5938), 
        .op(n5941) );
  ab_or_c_or_d U7063 ( .ip1(n5285), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[5]), .ip3(n5942), .ip4(n5941), 
        .op(n5943) );
  not_ab_or_c_or_d U7064 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[7]), 
        .ip2(n5527), .ip3(n5946), .ip4(n5945), .op(n5955) );
  xor2_1 U7065 ( .ip1(n5949), .ip2(n5948), .op(n6487) );
  inv_1 U7066 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[8]), .op(n5972)
         );
  and2_1 U7067 ( .ip1(n6487), .ip2(n5972), .op(n5954) );
  mux2_1 U7068 ( .ip1(i_i2c_ic_fs_lcnt[10]), .ip2(i_i2c_ic_lcnt[10]), .s(n5907), .op(n5951) );
  xor2_1 U7069 ( .ip1(n5951), .ip2(n5536), .op(n6495) );
  inv_1 U7070 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[10]), .op(n5979)
         );
  nand2_1 U7071 ( .ip1(n6495), .ip2(n5979), .op(n5953) );
  mux2_1 U7072 ( .ip1(i_i2c_ic_fs_lcnt[11]), .ip2(i_i2c_ic_lcnt[11]), .s(n5908), .op(n5956) );
  nor2_1 U7073 ( .ip1(n6498), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[11]), .op(n5978) );
  inv_1 U7074 ( .ip(n5978), .op(n5952) );
  nand2_1 U7075 ( .ip1(n5953), .ip2(n5952), .op(n5976) );
  or4_1 U7076 ( .ip1(n5971), .ip2(n5955), .ip3(n5954), .ip4(n5976), .op(n5970)
         );
  mux2_1 U7077 ( .ip1(i_i2c_ic_fs_lcnt[12]), .ip2(i_i2c_ic_lcnt[12]), .s(n5907), .op(n5960) );
  nand2_1 U7078 ( .ip1(n5246), .ip2(n5956), .op(n5957) );
  inv_1 U7079 ( .ip(n5957), .op(n5959) );
  xor2_1 U7080 ( .ip1(n5960), .ip2(n5959), .op(n6501) );
  inv_1 U7081 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[12]), .op(n5987)
         );
  mux2_1 U7082 ( .ip1(i_i2c_ic_fs_lcnt[14]), .ip2(i_i2c_ic_lcnt[14]), .s(n5907), .op(n5962) );
  mux2_1 U7083 ( .ip1(i_i2c_ic_fs_lcnt[13]), .ip2(i_i2c_ic_lcnt[13]), .s(n5908), .op(n5958) );
  inv_1 U7084 ( .ip(n5958), .op(n5969) );
  nand2_1 U7085 ( .ip1(n5960), .ip2(n5959), .op(n5967) );
  nor2_1 U7086 ( .ip1(n5969), .ip2(n5967), .op(n5961) );
  xor2_1 U7087 ( .ip1(n5962), .ip2(n5961), .op(n6453) );
  inv_1 U7088 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[14]), .op(n5996)
         );
  nand2_1 U7089 ( .ip1(n6453), .ip2(n5996), .op(n5966) );
  mux2_1 U7090 ( .ip1(i_i2c_ic_fs_lcnt[15]), .ip2(i_i2c_ic_lcnt[15]), .s(n5908), .op(n5964) );
  nand2_1 U7091 ( .ip1(n5962), .ip2(n5961), .op(n5963) );
  inv_1 U7092 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[15]), .op(n5965)
         );
  nand2_1 U7093 ( .ip1(n5966), .ip2(n5537), .op(n5992) );
  inv_1 U7094 ( .ip(n5967), .op(n5968) );
  xnor2_1 U7095 ( .ip1(n5969), .ip2(n5968), .op(n6502) );
  nor2_1 U7096 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[13]), .ip2(
        n5988), .op(n5986) );
  ab_or_c_or_d U7097 ( .ip1(n6501), .ip2(n5987), .ip3(n5992), .ip4(n5986), 
        .op(n5982) );
  nor2_1 U7098 ( .ip1(n5970), .ip2(n5982), .op(n5985) );
  nor2_1 U7099 ( .ip1(n5532), .ip2(n5973), .op(n5975) );
  nor2_1 U7100 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[9]), .ip2(n5973), .op(n5974) );
  or2_1 U7101 ( .ip1(n5974), .ip2(n5975), .op(n5977) );
  nor2_1 U7102 ( .ip1(n5977), .ip2(n5976), .op(n5981) );
  nor3_1 U7103 ( .ip1(n5979), .ip2(n6495), .ip3(n5978), .op(n5980) );
  not_ab_or_c_or_d U7104 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[11]), 
        .ip2(n6498), .ip3(n5981), .ip4(n5980), .op(n5983) );
  nor2_1 U7105 ( .ip1(n5982), .ip2(n5983), .op(n5984) );
  nor2_1 U7106 ( .ip1(n5984), .ip2(n5985), .op(n6004) );
  nor3_1 U7107 ( .ip1(n5987), .ip2(n5986), .ip3(n6501), .op(n5989) );
  nor2_1 U7108 ( .ip1(n5988), .ip2(n5989), .op(n5991) );
  nor2_1 U7109 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[13]), .ip2(
        n5989), .op(n5990) );
  or2_1 U7110 ( .ip1(n5991), .ip2(n5990), .op(n5993) );
  or2_1 U7111 ( .ip1(n5993), .ip2(n5992), .op(n6001) );
  inv_1 U7112 ( .ip(n5994), .op(n5995) );
  nor2_1 U7113 ( .ip1(n6451), .ip2(n5965), .op(n6504) );
  nor2_1 U7114 ( .ip1(n5997), .ip2(n6504), .op(n5998) );
  nand2_1 U7115 ( .ip1(n5998), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_count_en), .op(
        n5999) );
  inv_1 U7116 ( .ip(n5999), .op(n6000) );
  nand2_1 U7117 ( .ip1(n6000), .ip2(n6001), .op(n6002) );
  inv_1 U7118 ( .ip(n6002), .op(n6003) );
  nand2_1 U7119 ( .ip1(n6003), .ip2(n6004), .op(n7712) );
  nand2_1 U7120 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[1]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[0]), .op(n6005) );
  nand2_1 U7121 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[2]), .ip2(
        n7714), .op(n7716) );
  nand2_1 U7122 ( .ip1(n6006), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[5]), .op(n7698) );
  inv_1 U7123 ( .ip(n7698), .op(n6008) );
  nand2_1 U7124 ( .ip1(n6008), .ip2(n6007), .op(n7700) );
  inv_1 U7125 ( .ip(n7700), .op(n6009) );
  nand2_1 U7126 ( .ip1(n6009), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[8]), .op(n6010) );
  xor2_1 U7127 ( .ip1(n6012), .ip2(n7696), .op(n6013) );
  nor2_2 U7128 ( .ip1(n7729), .ip2(n6013), .op(i_i2c_U_DW_apb_i2c_clk_gen_N73)
         );
  nor2_1 U7129 ( .ip1(i_apb_paddr[31]), .ip2(i_apb_paddr[29]), .op(n6015) );
  nor2_1 U7130 ( .ip1(i_apb_paddr[24]), .ip2(i_apb_paddr[30]), .op(n6014) );
  nand2_1 U7131 ( .ip1(n6015), .ip2(n6014), .op(n6018) );
  nor2_1 U7132 ( .ip1(i_apb_paddr[27]), .ip2(i_apb_paddr[28]), .op(n6016) );
  nand2_1 U7133 ( .ip1(n6016), .ip2(i_apb_paddr[16]), .op(n6017) );
  nor2_1 U7134 ( .ip1(n6018), .ip2(n6017), .op(n6019) );
  nand4_1 U7135 ( .ip1(n6022), .ip2(n6021), .ip3(n6020), .ip4(n6019), .op(
        n11152) );
  inv_1 U7136 ( .ip(i_apb_pwrite), .op(n6024) );
  inv_1 U7137 ( .ip(i_apb_penable), .op(n6023) );
  and3_1 U7138 ( .ip1(n6024), .ip2(i_apb_psel_en), .ip3(n6023), .op(n6686) );
  inv_1 U7139 ( .ip(n6686), .op(n6025) );
  nand4_1 U7140 ( .ip1(i_ssi_reg_addr[5]), .ip2(i_ssi_reg_addr[4]), .ip3(
        i_ssi_reg_addr[3]), .ip4(i_ssi_reg_addr[2]), .op(n6028) );
  nand2_1 U7141 ( .ip1(i_ssi_reg_addr[4]), .ip2(i_ssi_reg_addr[3]), .op(n6026)
         );
  inv_1 U7142 ( .ip(i_ssi_reg_addr[5]), .op(n6685) );
  nand2_1 U7143 ( .ip1(n6026), .ip2(n6685), .op(n6027) );
  and2_1 U7144 ( .ip1(n6028), .ip2(n6027), .op(n11632) );
  inv_1 U7145 ( .ip(n11632), .op(n11590) );
  inv_1 U7146 ( .ip(i_apb_paddr[12]), .op(n6029) );
  and3_1 U7147 ( .ip1(i_apb_pwrite), .ip2(i_apb_penable), .ip3(i_apb_psel_en), 
        .op(n6030) );
  nand2_1 U7148 ( .ip1(n5616), .ip2(n6030), .op(n10139) );
  nor2_1 U7149 ( .ip1(n11590), .ip2(n10139), .op(n11854) );
  nand2_1 U7150 ( .ip1(n9817), .ip2(n10111), .op(n6032) );
  nand2_1 U7151 ( .ip1(n6032), .ip2(n6031), .op(n11836) );
  nor2_1 U7152 ( .ip1(n6033), .ip2(n9890), .op(n9895) );
  nor2_1 U7153 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv), .ip2(
        i_i2c_p_det), .op(n6037) );
  nand2_1 U7154 ( .ip1(n6037), .ip2(i_i2c_ic_enable_sync), .op(n6038) );
  or2_1 U7155 ( .ip1(n11833), .ip2(n6038), .op(n7774) );
  nand2_1 U7156 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[10]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[11]), .op(n7757) );
  nand2_1 U7157 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[7]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[8]), .op(n6304) );
  nor2_1 U7158 ( .ip1(i_i2c_ic_ss_sync), .ip2(i_i2c_ic_fs_sync), .op(n6040) );
  nand2_4 U7159 ( .ip1(n6040), .ip2(i_i2c_hs_mcode_en), .op(n6060) );
  buf_4 U7160 ( .ip(n6060), .op(n6270) );
  mux2_1 U7161 ( .ip1(i_i2c_ic_fs_hcnt[11]), .ip2(i_i2c_ic_hcnt[11]), .s(n6270), .op(n8265) );
  inv_1 U7162 ( .ip(n8265), .op(n6107) );
  or2_1 U7163 ( .ip1(i_i2c_ic_fs_spklen[1]), .ip2(i_i2c_ic_fs_spklen[2]), .op(
        n6058) );
  and2_1 U7164 ( .ip1(n6058), .ip2(i_i2c_ic_fs_spklen[3]), .op(n6049) );
  and2_1 U7165 ( .ip1(n6049), .ip2(i_i2c_ic_fs_spklen[4]), .op(n6050) );
  and2_1 U7166 ( .ip1(n6050), .ip2(i_i2c_ic_fs_spklen[5]), .op(n6042) );
  and2_1 U7167 ( .ip1(n6042), .ip2(i_i2c_ic_fs_spklen[6]), .op(n6045) );
  and2_1 U7168 ( .ip1(n6045), .ip2(i_i2c_ic_fs_spklen[7]), .op(n6125) );
  nand2_1 U7169 ( .ip1(n8258), .ip2(n6125), .op(n6130) );
  nand2_1 U7170 ( .ip1(n5454), .ip2(n8262), .op(n6080) );
  nor2_1 U7171 ( .ip1(n6130), .ip2(n6080), .op(n6096) );
  inv_1 U7172 ( .ip(n6096), .op(n6109) );
  nor2_1 U7173 ( .ip1(n6107), .ip2(n6109), .op(n6083) );
  xor2_1 U7174 ( .ip1(i_i2c_ic_fs_spklen[6]), .ip2(n6042), .op(n6053) );
  nand2_2 U7175 ( .ip1(n5282), .ip2(n6053), .op(n6173) );
  xor2_1 U7176 ( .ip1(i_i2c_ic_fs_spklen[7]), .ip2(n6045), .op(n6047) );
  inv_1 U7177 ( .ip(n6047), .op(n6046) );
  or2_1 U7178 ( .ip1(n6173), .ip2(n6055), .op(n6048) );
  nand2_2 U7179 ( .ip1(n5270), .ip2(n6047), .op(n6166) );
  and2_1 U7180 ( .ip1(n6048), .ip2(n6166), .op(n6057) );
  xor2_1 U7181 ( .ip1(i_i2c_ic_fs_spklen[4]), .ip2(n6049), .op(n6074) );
  nand2_2 U7182 ( .ip1(n8215), .ip2(n6074), .op(n6188) );
  inv_1 U7183 ( .ip(n6188), .op(n6183) );
  xor2_1 U7184 ( .ip1(i_i2c_ic_fs_spklen[5]), .ip2(n6050), .op(n6051) );
  nand2_1 U7185 ( .ip1(n8211), .ip2(n6051), .op(n6184) );
  nand2_1 U7186 ( .ip1(n6172), .ip2(n6077), .op(n6056) );
  xor2_1 U7187 ( .ip1(i_i2c_ic_fs_spklen[3]), .ip2(n6058), .op(n6061) );
  inv_1 U7188 ( .ip(n6061), .op(n6059) );
  nand2_1 U7189 ( .ip1(n5455), .ip2(n6059), .op(n6199) );
  inv_1 U7190 ( .ip(n6199), .op(n6070) );
  xnor2_1 U7191 ( .ip1(i_i2c_ic_fs_spklen[1]), .ip2(i_i2c_ic_fs_spklen[2]), 
        .op(n6069) );
  nand2_1 U7192 ( .ip1(n6063), .ip2(n6062), .op(n6064) );
  inv_1 U7193 ( .ip(n6064), .op(n6073) );
  nor2_1 U7194 ( .ip1(n5468), .ip2(n6069), .op(n6200) );
  nor2_1 U7195 ( .ip1(n6200), .ip2(n6070), .op(n6071) );
  nor2_1 U7196 ( .ip1(n6075), .ip2(n6076), .op(n6161) );
  and2_1 U7197 ( .ip1(n6161), .ip2(n6077), .op(n6078) );
  nand2_2 U7198 ( .ip1(n5260), .ip2(n6086), .op(n6131) );
  inv_1 U7199 ( .ip(n6108), .op(n6087) );
  nor2_1 U7200 ( .ip1(n6087), .ip2(n6107), .op(n6081) );
  and2_1 U7201 ( .ip1(n6131), .ip2(n6081), .op(n6082) );
  mux2_2 U7202 ( .ip1(i_i2c_ic_fs_hcnt[12]), .ip2(i_i2c_ic_hcnt[12]), .s(n6270), .op(n8188) );
  inv_1 U7203 ( .ip(n8188), .op(n6084) );
  nor2_1 U7204 ( .ip1(n8620), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[12]), .op(n6092) );
  mux2_1 U7205 ( .ip1(i_i2c_ic_fs_hcnt[13]), .ip2(i_i2c_ic_hcnt[13]), .s(n6270), .op(n8186) );
  inv_1 U7206 ( .ip(n8186), .op(n6093) );
  nand2_1 U7207 ( .ip1(n8265), .ip2(n8188), .op(n6094) );
  nor2_1 U7208 ( .ip1(n6094), .ip2(n6109), .op(n6090) );
  nand2_1 U7209 ( .ip1(n5260), .ip2(n6086), .op(n6126) );
  nor2_1 U7210 ( .ip1(n6087), .ip2(n6094), .op(n6088) );
  and2_1 U7211 ( .ip1(n6126), .ip2(n6088), .op(n6089) );
  nor2_1 U7212 ( .ip1(n6090), .ip2(n6089), .op(n6091) );
  nor2_1 U7213 ( .ip1(n8778), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[13]), .op(n6145) );
  nor2_1 U7214 ( .ip1(n6092), .ip2(n6145), .op(n6106) );
  nor2_1 U7215 ( .ip1(n6094), .ip2(n6093), .op(n6097) );
  nand2_1 U7216 ( .ip1(n6108), .ip2(n6097), .op(n6102) );
  inv_1 U7217 ( .ip(n6131), .op(n6095) );
  nand2_1 U7218 ( .ip1(n6097), .ip2(n6096), .op(n6101) );
  inv_1 U7219 ( .ip(n6101), .op(n6098) );
  mux2_1 U7220 ( .ip1(i_i2c_ic_fs_hcnt[14]), .ip2(i_i2c_ic_hcnt[14]), .s(n6270), .op(n8172) );
  inv_1 U7221 ( .ip(n8172), .op(n8173) );
  nor2_1 U7222 ( .ip1(n8773), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[14]), .op(n6105) );
  mux2_1 U7223 ( .ip1(i_i2c_ic_fs_hcnt[15]), .ip2(i_i2c_ic_hcnt[15]), .s(n6270), .op(n8178) );
  inv_1 U7224 ( .ip(n8178), .op(n6943) );
  nor2_1 U7225 ( .ip1(n8173), .ip2(n6101), .op(n6941) );
  nor2_1 U7226 ( .ip1(n6102), .ip2(n8173), .op(n6103) );
  and2_1 U7227 ( .ip1(n6131), .ip2(n6103), .op(n6940) );
  nor2_1 U7228 ( .ip1(n6941), .ip2(n6940), .op(n6104) );
  nor2_1 U7229 ( .ip1(n8772), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[15]), .op(n6141) );
  nor2_1 U7230 ( .ip1(n6105), .ip2(n6141), .op(n6149) );
  nand2_1 U7231 ( .ip1(n6106), .ip2(n6149), .op(n6156) );
  nand2_1 U7232 ( .ip1(n6131), .ip2(n6108), .op(n6110) );
  nand2_1 U7233 ( .ip1(n6110), .ip2(n6109), .op(n6111) );
  xor2_1 U7234 ( .ip1(n8265), .ip2(n6111), .op(n8757) );
  inv_1 U7235 ( .ip(n8757), .op(n6112) );
  nand2_1 U7236 ( .ip1(n6112), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[11]), .op(n6122) );
  nor2_1 U7237 ( .ip1(n6112), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[11]), .op(n6123) );
  nor2_1 U7238 ( .ip1(n6129), .ip2(n6130), .op(n6117) );
  nor2_1 U7239 ( .ip1(n8258), .ip2(n6125), .op(n6113) );
  nor2_1 U7240 ( .ip1(n6113), .ip2(n6129), .op(n6114) );
  nand2_1 U7241 ( .ip1(n6131), .ip2(n6114), .op(n6115) );
  inv_1 U7242 ( .ip(n8262), .op(n6118) );
  nand2_1 U7243 ( .ip1(n8761), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[10]), .op(n6120) );
  or2_1 U7244 ( .ip1(n6123), .ip2(n6120), .op(n6121) );
  nand2_1 U7245 ( .ip1(n6122), .ip2(n6121), .op(n6138) );
  nor2_1 U7246 ( .ip1(n8761), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[10]), .op(n6124) );
  nor2_1 U7247 ( .ip1(n6124), .ip2(n6123), .op(n6154) );
  nand2_1 U7248 ( .ip1(n6126), .ip2(n5599), .op(n6127) );
  nand2_1 U7249 ( .ip1(n6130), .ip2(n6127), .op(n6128) );
  nand2_1 U7250 ( .ip1(n5265), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[9]), .op(n6135) );
  nor2_1 U7251 ( .ip1(n5265), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[9]), 
        .op(n6152) );
  nand2_1 U7252 ( .ip1(n5599), .ip2(n6130), .op(n6132) );
  nand2_1 U7253 ( .ip1(n5264), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[8]), .op(n6133) );
  or2_1 U7254 ( .ip1(n6152), .ip2(n6133), .op(n6134) );
  nand2_1 U7255 ( .ip1(n6135), .ip2(n6134), .op(n6136) );
  and2_1 U7256 ( .ip1(n6154), .ip2(n6136), .op(n6137) );
  nor2_1 U7257 ( .ip1(n6138), .ip2(n6137), .op(n6139) );
  or2_1 U7258 ( .ip1(n6156), .ip2(n6139), .op(n6239) );
  nand2_1 U7259 ( .ip1(n8772), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[15]), .op(n6143) );
  nand2_1 U7260 ( .ip1(n8773), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[14]), .op(n6140) );
  or2_1 U7261 ( .ip1(n6141), .ip2(n6140), .op(n6142) );
  nand2_1 U7262 ( .ip1(n6143), .ip2(n6142), .op(n6151) );
  nand2_1 U7263 ( .ip1(n8778), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[13]), .op(n6147) );
  nand2_1 U7264 ( .ip1(n8620), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[12]), .op(n6144) );
  or2_1 U7265 ( .ip1(n6145), .ip2(n6144), .op(n6146) );
  nand2_1 U7266 ( .ip1(n6147), .ip2(n6146), .op(n6148) );
  and2_1 U7267 ( .ip1(n6149), .ip2(n6148), .op(n6150) );
  nor2_1 U7268 ( .ip1(n6151), .ip2(n6150), .op(n6238) );
  nor2_1 U7269 ( .ip1(i_i2c_ic_fs_sync), .ip2(n5562), .op(n7018) );
  inv_1 U7270 ( .ip(n5907), .op(n7146) );
  nand2_1 U7271 ( .ip1(n7018), .ip2(n7146), .op(n8835) );
  nor2_1 U7272 ( .ip1(n5264), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[8]), 
        .op(n6153) );
  nor2_1 U7273 ( .ip1(n6153), .ip2(n6152), .op(n6155) );
  nand2_1 U7274 ( .ip1(n6155), .ip2(n6154), .op(n6157) );
  nor2_1 U7275 ( .ip1(n6157), .ip2(n6156), .op(n6237) );
  inv_1 U7276 ( .ip(n6158), .op(n6174) );
  nand2_1 U7277 ( .ip1(n6172), .ip2(n6174), .op(n6159) );
  nand2_1 U7278 ( .ip1(n6173), .ip2(n6159), .op(n6165) );
  inv_1 U7279 ( .ip(n6161), .op(n6170) );
  inv_1 U7280 ( .ip(n6174), .op(n6162) );
  or2_1 U7281 ( .ip1(n6170), .ip2(n6162), .op(n6163) );
  nor2_1 U7282 ( .ip1(n6190), .ip2(n6163), .op(n6164) );
  nand2_1 U7283 ( .ip1(n6167), .ip2(n6166), .op(n6168) );
  nand2_1 U7284 ( .ip1(n5597), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[7]), .op(n6179) );
  nor2_1 U7285 ( .ip1(n5597), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[7]), 
        .op(n6180) );
  nor2_1 U7286 ( .ip1(n6190), .ip2(n6170), .op(n6171) );
  nor2_1 U7287 ( .ip1(n6172), .ip2(n6171), .op(n6176) );
  nand2_1 U7288 ( .ip1(n6174), .ip2(n6173), .op(n6175) );
  nand2_1 U7289 ( .ip1(n5598), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[6]), .op(n6177) );
  or2_1 U7290 ( .ip1(n6180), .ip2(n6177), .op(n6178) );
  nand2_1 U7291 ( .ip1(n6179), .ip2(n6178), .op(n6198) );
  nor2_1 U7292 ( .ip1(n5598), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[6]), 
        .op(n6181) );
  nor2_1 U7293 ( .ip1(n6181), .ip2(n6180), .op(n6230) );
  nor2_1 U7294 ( .ip1(n6183), .ip2(n6182), .op(n6187) );
  nand2_1 U7295 ( .ip1(n6185), .ip2(n6184), .op(n6186) );
  nand2_1 U7296 ( .ip1(n8800), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[5]), .op(n6195) );
  nor2_1 U7297 ( .ip1(n8800), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[5]), 
        .op(n6228) );
  inv_1 U7298 ( .ip(n6075), .op(n6189) );
  nand2_1 U7299 ( .ip1(n6189), .ip2(n6188), .op(n6192) );
  inv_1 U7300 ( .ip(n6190), .op(n6191) );
  nand2_1 U7301 ( .ip1(n8822), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[4]), .op(n6193) );
  or2_1 U7302 ( .ip1(n6228), .ip2(n6193), .op(n6194) );
  nand2_1 U7303 ( .ip1(n6195), .ip2(n6194), .op(n6196) );
  and2_1 U7304 ( .ip1(n6230), .ip2(n6196), .op(n6197) );
  nor2_1 U7305 ( .ip1(n6198), .ip2(n6197), .op(n6235) );
  nand2_1 U7306 ( .ip1(n6199), .ip2(n6062), .op(n6203) );
  inv_1 U7307 ( .ip(n6200), .op(n6204) );
  nand2_1 U7308 ( .ip1(n6205), .ip2(n6204), .op(n6201) );
  nand2_1 U7309 ( .ip1(n5413), .ip2(n6201), .op(n6202) );
  xnor2_1 U7310 ( .ip1(n6203), .ip2(n6202), .op(n6990) );
  nand2_1 U7311 ( .ip1(n5274), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[3]), .op(n6210) );
  nor2_1 U7312 ( .ip1(n5274), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[3]), 
        .op(n6222) );
  nand2_1 U7313 ( .ip1(n6204), .ip2(n5413), .op(n6207) );
  inv_1 U7314 ( .ip(n6205), .op(n6206) );
  nand2_1 U7315 ( .ip1(n8807), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[2]), .op(n6208) );
  or2_1 U7316 ( .ip1(n6222), .ip2(n6208), .op(n6209) );
  nand2_1 U7317 ( .ip1(n6210), .ip2(n6209), .op(n6227) );
  inv_1 U7318 ( .ip(n6211), .op(n6213) );
  nand2_1 U7319 ( .ip1(n6213), .ip2(n6212), .op(n6216) );
  nand2_1 U7320 ( .ip1(n8811), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[1]), .op(n6221) );
  or2_1 U7321 ( .ip1(n8229), .ip2(i_i2c_ic_fs_spklen[0]), .op(n6217) );
  nand2_1 U7322 ( .ip1(n6217), .ip2(n6215), .op(n6994) );
  nor2_1 U7323 ( .ip1(n8811), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[1]), 
        .op(n6219) );
  or2_1 U7324 ( .ip1(n6218), .ip2(n6219), .op(n6220) );
  nand2_1 U7325 ( .ip1(n6221), .ip2(n6220), .op(n6225) );
  nor2_1 U7326 ( .ip1(n8807), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[2]), 
        .op(n6223) );
  nor2_1 U7327 ( .ip1(n6223), .ip2(n6222), .op(n6224) );
  and2_1 U7328 ( .ip1(n6225), .ip2(n6224), .op(n6226) );
  nor2_1 U7329 ( .ip1(n6227), .ip2(n6226), .op(n6233) );
  nor2_1 U7330 ( .ip1(n8822), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[4]), 
        .op(n6229) );
  nor2_1 U7331 ( .ip1(n6229), .ip2(n6228), .op(n6231) );
  nand2_1 U7332 ( .ip1(n6231), .ip2(n6230), .op(n6232) );
  or2_1 U7333 ( .ip1(n6233), .ip2(n6232), .op(n6234) );
  nand2_1 U7334 ( .ip1(n6235), .ip2(n6234), .op(n6236) );
  nand4_1 U7335 ( .ip1(n6239), .ip2(n6238), .ip3(n8835), .ip4(n5600), .op(
        n6301) );
  nor2_1 U7336 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv), .ip2(n5562), 
        .op(n8911) );
  mux2_1 U7337 ( .ip1(i_i2c_ic_fs_lcnt[13]), .ip2(i_i2c_ic_lcnt[13]), .s(n6270), .op(n7044) );
  inv_1 U7338 ( .ip(n7044), .op(n6240) );
  inv_1 U7339 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[12]), .op(n6277)
         );
  nor2_1 U7340 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[13]), .ip2(n6240), .op(n6275) );
  mux2_1 U7341 ( .ip1(i_i2c_ic_fs_lcnt[12]), .ip2(i_i2c_ic_lcnt[12]), .s(n6270), .op(n7048) );
  nor3_1 U7342 ( .ip1(n6277), .ip2(n6275), .ip3(n7048), .op(n6241) );
  nor2_1 U7343 ( .ip1(n6240), .ip2(n6241), .op(n6243) );
  nor2_1 U7344 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[13]), .ip2(n6241), .op(n6242) );
  or2_1 U7345 ( .ip1(n6243), .ip2(n6242), .op(n6245) );
  mux2_1 U7346 ( .ip1(i_i2c_ic_fs_lcnt[14]), .ip2(i_i2c_ic_lcnt[14]), .s(n6270), .op(n7036) );
  inv_1 U7347 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[14]), .op(n6248)
         );
  nand2_1 U7348 ( .ip1(n7036), .ip2(n6248), .op(n6244) );
  mux2_1 U7349 ( .ip1(i_i2c_ic_fs_lcnt[15]), .ip2(i_i2c_ic_lcnt[15]), .s(n6270), .op(n7031) );
  inv_1 U7350 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[15]), .op(n6249)
         );
  nand2_1 U7351 ( .ip1(n7031), .ip2(n6249), .op(n6246) );
  nand2_1 U7352 ( .ip1(n6244), .ip2(n6246), .op(n6276) );
  nor2_1 U7353 ( .ip1(n6245), .ip2(n6276), .op(n6298) );
  inv_1 U7354 ( .ip(n6246), .op(n6247) );
  nor3_1 U7355 ( .ip1(n6248), .ip2(n7036), .ip3(n6247), .op(n6297) );
  nor2_1 U7356 ( .ip1(n7031), .ip2(n6249), .op(n6296) );
  nor2_1 U7357 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[9]), .ip2(n7071), 
        .op(n6279) );
  mux2_1 U7358 ( .ip1(i_i2c_ic_fs_lcnt[7]), .ip2(i_i2c_ic_lcnt[7]), .s(n6270), 
        .op(n7093) );
  inv_1 U7359 ( .ip(n7093), .op(n6269) );
  inv_1 U7360 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[6]), .op(n6266) );
  mux2_1 U7361 ( .ip1(i_i2c_ic_fs_lcnt[6]), .ip2(i_i2c_ic_lcnt[6]), .s(n6270), 
        .op(n7096) );
  nor2_1 U7362 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[7]), .ip2(n6269), 
        .op(n6264) );
  nor3_1 U7363 ( .ip1(n6266), .ip2(n7096), .ip3(n6264), .op(n6268) );
  inv_1 U7364 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[4]), .op(n6261) );
  nor2_1 U7365 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[5]), .ip2(n7104), 
        .op(n6260) );
  nor3_1 U7366 ( .ip1(n6261), .ip2(n6260), .ip3(n7105), .op(n6263) );
  mux2_1 U7367 ( .ip1(i_i2c_ic_fs_lcnt[3]), .ip2(i_i2c_ic_lcnt[3]), .s(n6270), 
        .op(n7114) );
  inv_1 U7368 ( .ip(n7114), .op(n6258) );
  inv_1 U7369 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[2]), .op(n6255) );
  and2_1 U7370 ( .ip1(n7116), .ip2(n6255), .op(n6253) );
  nor2_1 U7371 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[3]), .ip2(n6258), 
        .op(n6254) );
  inv_1 U7372 ( .ip(n7122), .op(n6250) );
  not_ab_or_c_or_d U7373 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[1]), 
        .ip2(n6250), .ip3(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[0]), .ip4(
        n7123), .op(n6252) );
  nor2_1 U7374 ( .ip1(n6250), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[1]), 
        .op(n6251) );
  nor3_1 U7375 ( .ip1(n6255), .ip2(n6254), .ip3(n7116), .op(n6256) );
  not_ab_or_c_or_d U7376 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[3]), 
        .ip2(n6258), .ip3(n6257), .ip4(n6256), .op(n6259) );
  not_ab_or_c_or_d U7377 ( .ip1(n7105), .ip2(n6261), .ip3(n6260), .ip4(n6259), 
        .op(n6262) );
  not_ab_or_c_or_d U7378 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[5]), 
        .ip2(n7104), .ip3(n6263), .ip4(n6262), .op(n6265) );
  not_ab_or_c_or_d U7379 ( .ip1(n7096), .ip2(n6266), .ip3(n6265), .ip4(n6264), 
        .op(n6267) );
  not_ab_or_c_or_d U7380 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[7]), 
        .ip2(n6269), .ip3(n6268), .ip4(n6267), .op(n6274) );
  inv_1 U7381 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[8]), .op(n6280) );
  and2_1 U7382 ( .ip1(n7072), .ip2(n6280), .op(n6273) );
  inv_1 U7383 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[10]), .op(n6287)
         );
  nand2_1 U7384 ( .ip1(n8550), .ip2(n6287), .op(n6272) );
  mux2_1 U7385 ( .ip1(i_i2c_ic_fs_lcnt[11]), .ip2(i_i2c_ic_lcnt[11]), .s(n6270), .op(n7062) );
  inv_1 U7386 ( .ip(n7062), .op(n6290) );
  nor2_1 U7387 ( .ip1(n6290), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[11]), .op(n6286) );
  inv_1 U7388 ( .ip(n6286), .op(n6271) );
  nand2_1 U7389 ( .ip1(n6272), .ip2(n6271), .op(n6284) );
  or4_1 U7390 ( .ip1(n6279), .ip2(n6274), .ip3(n6273), .ip4(n6284), .op(n6278)
         );
  ab_or_c_or_d U7391 ( .ip1(n7048), .ip2(n6277), .ip3(n6276), .ip4(n6275), 
        .op(n6291) );
  nor2_1 U7392 ( .ip1(n6278), .ip2(n6291), .op(n6294) );
  nor3_1 U7393 ( .ip1(n6280), .ip2(n6279), .ip3(n7072), .op(n6281) );
  nor2_1 U7394 ( .ip1(n7071), .ip2(n6281), .op(n6283) );
  nor2_1 U7395 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[9]), .ip2(n6281), 
        .op(n6282) );
  or2_1 U7396 ( .ip1(n6283), .ip2(n6282), .op(n6285) );
  nor2_1 U7397 ( .ip1(n6285), .ip2(n6284), .op(n6289) );
  nor3_1 U7398 ( .ip1(n6287), .ip2(n8550), .ip3(n6286), .op(n6288) );
  not_ab_or_c_or_d U7399 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[11]), 
        .ip2(n6290), .ip3(n6289), .ip4(n6288), .op(n6292) );
  nor2_1 U7400 ( .ip1(n6292), .ip2(n6291), .op(n6293) );
  or2_1 U7401 ( .ip1(n6294), .ip2(n6293), .op(n6295) );
  nand2_1 U7402 ( .ip1(n8911), .ip2(n6299), .op(n6300) );
  nand2_1 U7403 ( .ip1(n6301), .ip2(n6300), .op(n7771) );
  nand2_1 U7404 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[1]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[2]), .op(n6302) );
  nand2_1 U7405 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[3]), .ip2(n7739), .op(n7743) );
  nand2_1 U7406 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[4]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[5]), .op(n6303) );
  nand2_1 U7407 ( .ip1(n7747), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[6]), .op(n7750) );
  nor2_1 U7408 ( .ip1(n6304), .ip2(n7750), .op(n7753) );
  inv_1 U7409 ( .ip(i_ssi_tx_wr_addr[0]), .op(n10198) );
  nor2_2 U7410 ( .ip1(n10198), .ip2(n10199), .op(n10228) );
  nand2_1 U7411 ( .ip1(i_apb_pwdata_int[10]), .ip2(n10354), .op(n6312) );
  inv_1 U7412 ( .ip(i_ssi_U_dff_tx_mem[74]), .op(n6310) );
  or2_1 U7413 ( .ip1(n10354), .ip2(n6310), .op(n6311) );
  nand2_1 U7414 ( .ip1(n6312), .ip2(n6311), .op(n4502) );
  inv_1 U7415 ( .ip(i_ssi_tx_wr_addr[2]), .op(n10220) );
  nand2_1 U7416 ( .ip1(i_apb_pwdata_int[10]), .ip2(n5608), .op(n6315) );
  inv_1 U7417 ( .ip(i_ssi_U_dff_tx_mem[10]), .op(n6313) );
  or2_1 U7418 ( .ip1(n5608), .ip2(n6313), .op(n6314) );
  nand2_1 U7419 ( .ip1(n6315), .ip2(n6314), .op(n4566) );
  nand2_1 U7420 ( .ip1(i_apb_pwdata_int[13]), .ip2(n10354), .op(n6318) );
  inv_1 U7421 ( .ip(i_ssi_U_dff_tx_mem[77]), .op(n6316) );
  or2_1 U7422 ( .ip1(n10354), .ip2(n6316), .op(n6317) );
  nand2_1 U7423 ( .ip1(n6318), .ip2(n6317), .op(n4499) );
  nand2_1 U7424 ( .ip1(i_apb_pwdata_int[13]), .ip2(n5608), .op(n6321) );
  inv_1 U7425 ( .ip(i_ssi_U_dff_tx_mem[13]), .op(n6319) );
  or2_1 U7426 ( .ip1(n5608), .ip2(n6319), .op(n6320) );
  nand2_1 U7427 ( .ip1(n6321), .ip2(n6320), .op(n4563) );
  inv_1 U7428 ( .ip(i_apb_pwdata_int[4]), .op(n10959) );
  nand2_1 U7429 ( .ip1(i_apb_pwdata_int[4]), .ip2(n10354), .op(n6324) );
  inv_1 U7430 ( .ip(i_ssi_U_dff_tx_mem[68]), .op(n6322) );
  or2_1 U7431 ( .ip1(n10354), .ip2(n6322), .op(n6323) );
  nand2_1 U7432 ( .ip1(n6324), .ip2(n6323), .op(n4508) );
  nand2_1 U7433 ( .ip1(i_apb_pwdata_int[4]), .ip2(n5608), .op(n6327) );
  inv_1 U7434 ( .ip(i_ssi_U_dff_tx_mem[4]), .op(n6325) );
  or2_1 U7435 ( .ip1(n5608), .ip2(n6325), .op(n6326) );
  nand2_1 U7436 ( .ip1(n6327), .ip2(n6326), .op(n4572) );
  nand2_1 U7437 ( .ip1(i_apb_pwdata_int[6]), .ip2(n5608), .op(n6330) );
  inv_1 U7438 ( .ip(i_ssi_U_dff_tx_mem[6]), .op(n6328) );
  or2_1 U7439 ( .ip1(n5608), .ip2(n6328), .op(n6329) );
  nand2_1 U7440 ( .ip1(n6330), .ip2(n6329), .op(n4570) );
  nand2_1 U7441 ( .ip1(i_apb_pwdata_int[3]), .ip2(n5608), .op(n6333) );
  inv_1 U7442 ( .ip(i_ssi_U_dff_tx_mem[3]), .op(n6331) );
  or2_1 U7443 ( .ip1(n5608), .ip2(n6331), .op(n6332) );
  nand2_1 U7444 ( .ip1(n6333), .ip2(n6332), .op(n4573) );
  nand2_1 U7445 ( .ip1(i_apb_pwdata_int[6]), .ip2(n10354), .op(n6336) );
  inv_1 U7446 ( .ip(i_ssi_U_dff_tx_mem[70]), .op(n6334) );
  or2_1 U7447 ( .ip1(n10354), .ip2(n6334), .op(n6335) );
  nand2_1 U7448 ( .ip1(n6336), .ip2(n6335), .op(n4506) );
  nand2_1 U7449 ( .ip1(i_apb_pwdata_int[1]), .ip2(n10354), .op(n6340) );
  inv_1 U7450 ( .ip(i_ssi_U_dff_tx_mem[65]), .op(n6338) );
  or2_1 U7451 ( .ip1(n10354), .ip2(n6338), .op(n6339) );
  nand2_1 U7452 ( .ip1(n6340), .ip2(n6339), .op(n4511) );
  nand2_1 U7453 ( .ip1(i_apb_pwdata_int[1]), .ip2(n5608), .op(n6343) );
  inv_1 U7454 ( .ip(i_ssi_U_dff_tx_mem[1]), .op(n6341) );
  or2_1 U7455 ( .ip1(n5608), .ip2(n6341), .op(n6342) );
  nand2_1 U7456 ( .ip1(n6343), .ip2(n6342), .op(n4575) );
  inv_1 U7457 ( .ip(i_i2c_mst_debug_cstate[1]), .op(n7918) );
  nand2_1 U7458 ( .ip1(n7918), .ip2(i_i2c_mst_debug_cstate[2]), .op(n7683) );
  nor2_1 U7459 ( .ip1(i_i2c_mst_debug_cstate[4]), .ip2(n7683), .op(n6360) );
  and2_1 U7460 ( .ip1(n6360), .ip2(n7685), .op(n7858) );
  inv_1 U7461 ( .ip(i_i2c_U_DW_apb_i2c_mstfsm_delay_stop_en), .op(n6344) );
  nand2_1 U7462 ( .ip1(n7858), .ip2(n6344), .op(n6347) );
  nand2_1 U7463 ( .ip1(i_i2c_mst_debug_cstate[0]), .ip2(
        i_i2c_mst_debug_cstate[3]), .op(n6345) );
  nor2_1 U7464 ( .ip1(n6345), .ip2(n6358), .op(n7856) );
  inv_1 U7465 ( .ip(n7856), .op(n6346) );
  nand2_1 U7466 ( .ip1(n6347), .ip2(n6346), .op(n6348) );
  inv_1 U7467 ( .ip(i_i2c_byte_wait_scl), .op(n7401) );
  and2_1 U7468 ( .ip1(n6348), .ip2(n7401), .op(n11857) );
  or2_1 U7469 ( .ip1(i_i2c_re_start_en), .ip2(i_i2c_start_en), .op(
        i_i2c_U_DW_apb_i2c_toggle_N30) );
  nor2_1 U7470 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_mst_tx_bwen), .ip2(
        i_i2c_mst_rx_bwen), .op(n6349) );
  nor4_1 U7471 ( .ip1(n11857), .ip2(n6349), .ip3(i_i2c_U_DW_apb_i2c_toggle_N30), .ip4(n6352), .op(i_i2c_U_DW_apb_i2c_tx_shift_byte_wait_en) );
  inv_1 U7472 ( .ip(n6352), .op(n9533) );
  inv_1 U7473 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_sda_int_q), .op(n7709) );
  inv_1 U7474 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_scl_int_q), .op(n8065) );
  nor4_1 U7475 ( .ip1(n9533), .ip2(n7709), .ip3(n8065), .ip4(n11833), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_s_det_int) );
  nor2_1 U7476 ( .ip1(i_i2c_mst_debug_cstate[0]), .ip2(
        i_i2c_mst_debug_cstate[3]), .op(n6350) );
  and2_1 U7477 ( .ip1(n6350), .ip2(n7684), .op(n7919) );
  inv_1 U7478 ( .ip(n7919), .op(n7778) );
  and2_1 U7479 ( .ip1(n7917), .ip2(i_i2c_mst_debug_cstate[1]), .op(n7802) );
  nand2_1 U7480 ( .ip1(n7802), .ip2(n7829), .op(n11062) );
  inv_1 U7481 ( .ip(i_i2c_ack_det), .op(n8068) );
  nor2_1 U7482 ( .ip1(n6353), .ip2(n6352), .op(n6354) );
  inv_1 U7483 ( .ip(n5591), .op(n8145) );
  or2_1 U7484 ( .ip1(n8068), .ip2(n9473), .op(n11073) );
  nor2_1 U7485 ( .ip1(n11062), .ip2(n11073), .op(n6382) );
  inv_1 U7486 ( .ip(i_i2c_U_DW_apb_i2c_sync_tx_empty_int_inv), .op(n11861) );
  inv_1 U7487 ( .ip(i_i2c_mst_rxbyte_rdy), .op(n8055) );
  nand2_1 U7488 ( .ip1(i_i2c_ic_abort_sync), .ip2(
        i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_chk_win), .op(n6357) );
  nand2_1 U7489 ( .ip1(n6357), .ip2(i_i2c_U_DW_apb_i2c_mstfsm_byte_waiting_q), 
        .op(n7853) );
  inv_1 U7490 ( .ip(n6358), .op(n7793) );
  nand2_1 U7491 ( .ip1(n7793), .ip2(n7685), .op(n11021) );
  nor2_1 U7492 ( .ip1(n7853), .ip2(n11021), .op(n7865) );
  nand2_1 U7493 ( .ip1(n7865), .ip2(i_i2c_tx_fifo_data_buf[8]), .op(n8126) );
  nor2_1 U7494 ( .ip1(n8055), .ip2(n8126), .op(n6368) );
  inv_1 U7495 ( .ip(n6359), .op(n11068) );
  inv_1 U7496 ( .ip(n11068), .op(n10941) );
  inv_1 U7497 ( .ip(i_i2c_ic_abort_sync), .op(n8105) );
  and2_1 U7498 ( .ip1(n10941), .ip2(n8105), .op(n7791) );
  inv_1 U7499 ( .ip(i_i2c_tx_fifo_data_buf[8]), .op(n11055) );
  inv_1 U7500 ( .ip(i_i2c_mst_debug_cstate[0]), .op(n7830) );
  and2_1 U7501 ( .ip1(n6360), .ip2(n7830), .op(n8109) );
  inv_1 U7502 ( .ip(n8109), .op(n8746) );
  inv_1 U7503 ( .ip(n10942), .op(n11071) );
  nor2_1 U7504 ( .ip1(n11055), .ip2(n11071), .op(n6364) );
  and2_1 U7505 ( .ip1(n6360), .ip2(i_i2c_mst_debug_cstate[3]), .op(n10943) );
  inv_1 U7506 ( .ip(n10943), .op(n11023) );
  inv_1 U7507 ( .ip(i_i2c_U_DW_apb_i2c_mstfsm_old_is_read), .op(n6361) );
  nand3_1 U7508 ( .ip1(n6361), .ip2(i_i2c_tx_fifo_data_buf[8]), .ip3(
        i_i2c_U_DW_apb_i2c_mstfsm_addr_2byte_sent), .op(n7875) );
  inv_1 U7509 ( .ip(n7875), .op(n6362) );
  nand2_1 U7510 ( .ip1(n10919), .ip2(n6362), .op(n7810) );
  inv_1 U7511 ( .ip(n7810), .op(n6363) );
  nor2_1 U7512 ( .ip1(n6364), .ip2(n6363), .op(n10932) );
  inv_1 U7513 ( .ip(n10932), .op(n6365) );
  nor2_1 U7514 ( .ip1(n7791), .ip2(n6365), .op(n6366) );
  nor2_1 U7515 ( .ip1(n6366), .ip2(n11073), .op(n6367) );
  nor2_1 U7516 ( .ip1(n6368), .ip2(n6367), .op(n6369) );
  nor2_1 U7517 ( .ip1(n11861), .ip2(n6369), .op(n6381) );
  nor2_1 U7518 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_slv_arb_lost), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_mst_arb_lost), .op(n8985) );
  nand2_1 U7519 ( .ip1(n8985), .ip2(n11055), .op(n10145) );
  inv_1 U7520 ( .ip(n10145), .op(n6370) );
  nand2_1 U7521 ( .ip1(n6370), .ip2(i_i2c_slv_tx_cmplt), .op(n6371) );
  inv_1 U7522 ( .ip(i_i2c_slv_debug_cstate[3]), .op(n11019) );
  and3_1 U7523 ( .ip1(n11019), .ip2(i_i2c_slv_debug_cstate[1]), .ip3(
        i_i2c_slv_debug_cstate[2]), .op(n7272) );
  and2_1 U7524 ( .ip1(n7272), .ip2(i_i2c_slv_debug_cstate[0]), .op(n11272) );
  or2_1 U7525 ( .ip1(i_i2c_s_det), .ip2(i_i2c_p_det), .op(n11083) );
  inv_1 U7526 ( .ip(n11083), .op(n9577) );
  nand2_1 U7527 ( .ip1(n11272), .ip2(n9577), .op(n11057) );
  nor2_1 U7528 ( .ip1(n6371), .ip2(n11057), .op(n10140) );
  nand2_1 U7529 ( .ip1(n10140), .ip2(i_i2c_slv_ack_det), .op(n9567) );
  nor2_1 U7530 ( .ip1(n11861), .ip2(n9567), .op(n9598) );
  nand2_1 U7531 ( .ip1(i_i2c_scl_s_hld_cmplt), .ip2(i_i2c_scl_s_setup_cmplt), 
        .op(n7868) );
  and2_1 U7532 ( .ip1(n7830), .ip2(i_i2c_mst_debug_cstate[3]), .op(n7874) );
  nand2_1 U7533 ( .ip1(n7793), .ip2(n7874), .op(n7844) );
  nor2_1 U7534 ( .ip1(n7868), .ip2(n7844), .op(n6373) );
  inv_1 U7535 ( .ip(n7895), .op(n11127) );
  nor2_1 U7536 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_N252), .ip2(n11127), .op(n6372) );
  nor2_1 U7537 ( .ip1(n6373), .ip2(n6372), .op(n7889) );
  inv_1 U7538 ( .ip(n7889), .op(n6374) );
  nand3_1 U7539 ( .ip1(n6374), .ip2(i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv), 
        .ip3(i_i2c_scl_s_hld_cmplt), .op(n6379) );
  nor2_1 U7540 ( .ip1(i_i2c_slv_debug_cstate[0]), .ip2(n11083), .op(n6375) );
  nand2_1 U7541 ( .ip1(n7272), .ip2(n6375), .op(n9565) );
  inv_1 U7542 ( .ip(n9565), .op(n6377) );
  inv_1 U7543 ( .ip(i_i2c_U_DW_apb_i2c_sync_tx_empty_sync_r), .op(n8099) );
  nand2_1 U7544 ( .ip1(n8099), .ip2(i_i2c_U_DW_apb_i2c_slvfsm_slv_tx_flush), 
        .op(n6376) );
  and2_1 U7545 ( .ip1(n6376), .ip2(i_i2c_U_DW_apb_i2c_sync_tx_empty_int_inv), 
        .op(n9566) );
  nand2_1 U7546 ( .ip1(n6377), .ip2(n9566), .op(n7969) );
  inv_1 U7547 ( .ip(n7869), .op(n7831) );
  inv_1 U7548 ( .ip(n7868), .op(n7845) );
  nand3_1 U7549 ( .ip1(n7831), .ip2(n7845), .ip3(n7874), .op(n6378) );
  nand3_1 U7550 ( .ip1(n6379), .ip2(n7969), .ip3(n6378), .op(n6380) );
  or4_1 U7551 ( .ip1(n6382), .ip2(n6381), .ip3(n9598), .ip4(n6380), .op(
        i_i2c_U_DW_apb_i2c_tx_shift_N90) );
  inv_1 U7552 ( .ip(i_ssi_U_sclkgen_ssi_cnt[13]), .op(n9784) );
  nor2_1 U7553 ( .ip1(i_ssi_baudr[3]), .ip2(i_ssi_baudr[4]), .op(n6383) );
  nor2_1 U7554 ( .ip1(i_ssi_baudr[8]), .ip2(i_ssi_baudr[7]), .op(n6384) );
  nor2_1 U7555 ( .ip1(i_ssi_baudr[6]), .ip2(i_ssi_baudr[5]), .op(n6396) );
  nand2_1 U7556 ( .ip1(n6384), .ip2(n6396), .op(n6385) );
  nor2_1 U7557 ( .ip1(n6423), .ip2(n6385), .op(n6415) );
  nor2_1 U7558 ( .ip1(i_ssi_baudr[11]), .ip2(i_ssi_baudr[12]), .op(n6386) );
  nor2_1 U7559 ( .ip1(i_ssi_baudr[10]), .ip2(i_ssi_baudr[9]), .op(n6412) );
  nand2_1 U7560 ( .ip1(n6386), .ip2(n6412), .op(n6407) );
  nor2_1 U7561 ( .ip1(n6407), .ip2(i_ssi_baudr[13]), .op(n6387) );
  nand2_1 U7562 ( .ip1(n6415), .ip2(n6387), .op(n7379) );
  xor2_1 U7563 ( .ip1(i_ssi_baudr[14]), .ip2(n7379), .op(n6388) );
  xor2_1 U7564 ( .ip1(n9784), .ip2(n6388), .op(n6447) );
  inv_1 U7565 ( .ip(i_ssi_U_sclkgen_ssi_cnt[14]), .op(n9791) );
  inv_1 U7566 ( .ip(i_ssi_baudr[14]), .op(n6390) );
  inv_1 U7567 ( .ip(i_ssi_baudr[13]), .op(n6389) );
  nand2_1 U7568 ( .ip1(n6390), .ip2(n6389), .op(n6391) );
  nor2_1 U7569 ( .ip1(n6407), .ip2(n6391), .op(n6392) );
  nand2_1 U7570 ( .ip1(n6415), .ip2(n6392), .op(n6393) );
  xor2_1 U7571 ( .ip1(n6415), .ip2(i_ssi_baudr[9]), .op(n6395) );
  xnor2_1 U7572 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[8]), .ip2(n6395), .op(n6404) );
  nand2_1 U7573 ( .ip1(n6397), .ip2(n6396), .op(n6398) );
  xnor2_1 U7574 ( .ip1(i_ssi_baudr[7]), .ip2(n6398), .op(n6399) );
  xnor2_1 U7575 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[6]), .ip2(n6399), .op(n6403) );
  nand2_1 U7576 ( .ip1(n6415), .ip2(n6412), .op(n6400) );
  xnor2_1 U7577 ( .ip1(i_ssi_baudr[11]), .ip2(n6400), .op(n6401) );
  xnor2_1 U7578 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[10]), .ip2(n6401), .op(n6402)
         );
  and3_1 U7579 ( .ip1(n6404), .ip2(n6403), .ip3(n6402), .op(n6411) );
  xor2_1 U7580 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[9]), .ip2(i_ssi_baudr[10]), .op(
        n10996) );
  inv_1 U7581 ( .ip(i_ssi_baudr[9]), .op(n6405) );
  nand2_1 U7582 ( .ip1(n6415), .ip2(n6405), .op(n6406) );
  inv_1 U7583 ( .ip(i_ssi_U_sclkgen_ssi_cnt[12]), .op(n9783) );
  inv_1 U7584 ( .ip(n6407), .op(n6408) );
  nand2_1 U7585 ( .ip1(n6415), .ip2(n6408), .op(n7354) );
  xor2_1 U7586 ( .ip1(i_ssi_baudr[13]), .ip2(n7354), .op(n6409) );
  xnor2_1 U7587 ( .ip1(n9783), .ip2(n6409), .op(n6410) );
  nand3_1 U7588 ( .ip1(n6411), .ip2(n5515), .ip3(n6410), .op(n6445) );
  inv_1 U7589 ( .ip(n6412), .op(n6413) );
  nor2_1 U7590 ( .ip1(n6413), .ip2(i_ssi_baudr[11]), .op(n6414) );
  nand2_1 U7591 ( .ip1(n6415), .ip2(n6414), .op(n7373) );
  xor2_1 U7592 ( .ip1(i_ssi_baudr[12]), .ip2(n7373), .op(n6416) );
  xor2_1 U7593 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[11]), .ip2(n6416), .op(n6443) );
  xor2_1 U7594 ( .ip1(i_ssi_baudr[1]), .ip2(i_ssi_baudr[2]), .op(n6417) );
  xor2_1 U7595 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[1]), .ip2(n6417), .op(n6418) );
  buf_2 U7596 ( .ip(i_ssi_ssi_en_int), .op(n10802) );
  xor2_1 U7597 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[0]), .ip2(i_ssi_baudr[1]), .op(
        n11004) );
  inv_1 U7598 ( .ip(i_ssi_U_sclkgen_ssi_cnt[15]), .op(n7394) );
  inv_1 U7599 ( .ip(n7329), .op(n6428) );
  nor2_1 U7600 ( .ip1(n6428), .ip2(i_ssi_baudr[3]), .op(n6420) );
  xnor2_1 U7601 ( .ip1(n6421), .ip2(n6420), .op(n6426) );
  xnor2_1 U7602 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[2]), .ip2(n6429), .op(n6430) );
  inv_1 U7603 ( .ip(i_ssi_baudr[4]), .op(n6434) );
  nand2_1 U7604 ( .ip1(n5356), .ip2(n6434), .op(n6436) );
  nor2_1 U7605 ( .ip1(i_ssi_baudr[1]), .ip2(n6436), .op(n7340) );
  inv_1 U7606 ( .ip(i_ssi_baudr[5]), .op(n10008) );
  nand2_1 U7607 ( .ip1(n7340), .ip2(n10008), .op(n7366) );
  xor2_1 U7608 ( .ip1(i_ssi_baudr[6]), .ip2(n7366), .op(n6435) );
  xor2_1 U7609 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[5]), .ip2(n6435), .op(n6441) );
  inv_1 U7610 ( .ip(n6436), .op(n9747) );
  inv_1 U7611 ( .ip(i_ssi_baudr[1]), .op(n10973) );
  nand2_1 U7612 ( .ip1(n10973), .ip2(n10008), .op(n6437) );
  or2_1 U7613 ( .ip1(i_ssi_baudr[6]), .ip2(i_ssi_baudr[7]), .op(n9752) );
  nor2_1 U7614 ( .ip1(n6437), .ip2(n9752), .op(n6438) );
  nand2_1 U7615 ( .ip1(n9747), .ip2(n6438), .op(n7361) );
  xor2_1 U7616 ( .ip1(i_ssi_baudr[8]), .ip2(n7361), .op(n6439) );
  xor2_1 U7617 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[7]), .ip2(n6439), .op(n6440) );
  nand4_1 U7618 ( .ip1(n6443), .ip2(n6442), .ip3(n6441), .ip4(n6440), .op(
        n6444) );
  nor4_1 U7619 ( .ip1(n6447), .ip2(n6446), .ip3(n6445), .ip4(n6444), .op(
        i_ssi_U_sclkgen_N74) );
  nand2_1 U7620 ( .ip1(n7919), .ip2(n6448), .op(i_i2c_U_DW_apb_i2c_mstfsm_N487) );
  nor2_1 U7621 ( .ip1(i_i2c_slv_tx_cmplt), .ip2(n10145), .op(n6449) );
  and2_1 U7622 ( .ip1(n11272), .ip2(n6449), .op(n11859) );
  inv_1 U7623 ( .ip(n6453), .op(n6450) );
  nor3_1 U7624 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[14]), .ip2(
        n6450), .ip3(n6504), .op(n6509) );
  inv_1 U7625 ( .ip(n6451), .op(n6452) );
  nor2_1 U7626 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[15]), .ip2(
        n6452), .op(n6508) );
  nor2_1 U7627 ( .ip1(n5996), .ip2(n6453), .op(n6506) );
  nor2_1 U7628 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[13]), .ip2(
        n5988), .op(n6500) );
  nor2_1 U7629 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[11]), .ip2(
        n6498), .op(n6494) );
  inv_1 U7630 ( .ip(n6495), .op(n6492) );
  nor2_1 U7631 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[9]), .ip2(n5532), .op(n6486) );
  inv_1 U7632 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[7]), .op(n7702)
         );
  nand2_1 U7633 ( .ip1(n7702), .ip2(n6480), .op(n6484) );
  nand2_1 U7634 ( .ip1(n5285), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[5]), .op(n6471) );
  nand3_1 U7635 ( .ip1(n6471), .ip2(n6455), .ip3(n5940), .op(n6475) );
  inv_1 U7636 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[5]), .op(n7719)
         );
  nand2_1 U7637 ( .ip1(n6454), .ip2(n7719), .op(n6474) );
  inv_1 U7638 ( .ip(n6455), .op(n6469) );
  nor2_1 U7639 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[3]), .ip2(n5937), .op(n6464) );
  inv_1 U7640 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[1]), .op(n7708)
         );
  nand2_1 U7641 ( .ip1(n6458), .ip2(n7708), .op(n6462) );
  inv_1 U7642 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[0]), .op(n6456)
         );
  nand2_1 U7643 ( .ip1(n6457), .ip2(n6456), .op(n6461) );
  nor2_1 U7644 ( .ip1(n5934), .ip2(n6465), .op(n6460) );
  nor2_1 U7645 ( .ip1(n7708), .ip2(n6458), .op(n6459) );
  not_ab_or_c_or_d U7646 ( .ip1(n6462), .ip2(n6461), .ip3(n6460), .ip4(n6459), 
        .op(n6463) );
  not_ab_or_c_or_d U7647 ( .ip1(n6465), .ip2(n5934), .ip3(n6464), .ip4(n6463), 
        .op(n6468) );
  nor2_1 U7648 ( .ip1(n5927), .ip2(n6466), .op(n6467) );
  not_ab_or_c_or_d U7649 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[4]), 
        .ip2(n6469), .ip3(n6468), .ip4(n6467), .op(n6470) );
  nand2_1 U7650 ( .ip1(n6471), .ip2(n6470), .op(n6473) );
  nand4_1 U7651 ( .ip1(n6475), .ip2(n6474), .ip3(n6473), .ip4(n6472), .op(
        n6479) );
  inv_1 U7652 ( .ip(n6476), .op(n6477) );
  nand2_1 U7653 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[6]), .ip2(
        n6477), .op(n6478) );
  nand2_1 U7654 ( .ip1(n6479), .ip2(n6478), .op(n6483) );
  nor2_1 U7655 ( .ip1(n5972), .ip2(n6487), .op(n6482) );
  nor2_1 U7656 ( .ip1(n7702), .ip2(n6480), .op(n6481) );
  not_ab_or_c_or_d U7657 ( .ip1(n6484), .ip2(n6483), .ip3(n6482), .ip4(n6481), 
        .op(n6485) );
  not_ab_or_c_or_d U7658 ( .ip1(n6487), .ip2(n5972), .ip3(n6486), .ip4(n6485), 
        .op(n6491) );
  inv_1 U7659 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[9]), .op(n6489)
         );
  nor2_1 U7660 ( .ip1(n6489), .ip2(n6488), .op(n6490) );
  not_ab_or_c_or_d U7661 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[10]), 
        .ip2(n6492), .ip3(n6491), .ip4(n6490), .op(n6493) );
  not_ab_or_c_or_d U7662 ( .ip1(n6495), .ip2(n5979), .ip3(n6494), .ip4(n6493), 
        .op(n6497) );
  nor2_1 U7663 ( .ip1(n5987), .ip2(n6501), .op(n6496) );
  not_ab_or_c_or_d U7664 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[11]), 
        .ip2(n6498), .ip3(n6497), .ip4(n6496), .op(n6499) );
  not_ab_or_c_or_d U7665 ( .ip1(n6501), .ip2(n5987), .ip3(n6500), .ip4(n6499), 
        .op(n6505) );
  inv_1 U7666 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[13]), .op(n7694)
         );
  nor2_1 U7667 ( .ip1(n7694), .ip2(n6502), .op(n6503) );
  inv_1 U7668 ( .ip(i_i2c_ic_enable_sync), .op(n11018) );
  inv_1 U7669 ( .ip(i_ahb_U_mux_hsel_prev[3]), .op(n6510) );
  nand2_1 U7670 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hresp[0]), .op(
        n6515) );
  nand2_1 U7671 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hresp[0]), .op(n6514) );
  nor4_1 U7672 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(i_ahb_U_mux_hsel_prev[3]), .ip3(i_ahb_U_mux_hsel_prev[2]), .ip4(i_ahb_U_mux_hsel_prev[1]), .op(n6678)
         );
  nand2_1 U7673 ( .ip1(n6678), .ip2(i_ahb_hresp_none_0_), .op(n6513) );
  inv_1 U7674 ( .ip(i_ahb_U_mux_hsel_prev[1]), .op(n6511) );
  nand2_1 U7675 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hresp[0]), .op(
        n6512) );
  nand4_1 U7676 ( .ip1(n6515), .ip2(n6514), .ip3(n6513), .ip4(n6512), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hresp[0]) );
  nand2_1 U7677 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[31]), .op(
        n6520) );
  nand2_1 U7678 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[31]), .op(n6519) );
  nand2_1 U7679 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[31]), .op(
        n6518) );
  inv_1 U7680 ( .ip(i_ahb_U_mux_hsel_prev[2]), .op(n6516) );
  and2_1 U7681 ( .ip1(n5616), .ip2(n6676), .op(n6521) );
  nand2_1 U7682 ( .ip1(n6521), .ip2(i_ssi_prdata[31]), .op(n6517) );
  nand2_1 U7683 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[27]), .op(n6525) );
  nand2_1 U7684 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[27]), .op(
        n6524) );
  nand2_1 U7685 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[27]), .op(
        n6523) );
  nand2_1 U7686 ( .ip1(n6521), .ip2(i_ssi_prdata[27]), .op(n6522) );
  mux2_1 U7687 ( .ip1(i_i2c_prdata[8]), .ip2(i_ssi_prdata[8]), .s(n5616), .op(
        n6526) );
  nand2_1 U7688 ( .ip1(n6676), .ip2(n6526), .op(n6530) );
  nand2_1 U7689 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[8]), .op(
        n6529) );
  nand2_1 U7690 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[8]), .op(
        n6528) );
  nand2_1 U7691 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[8]), .op(n6527) );
  mux2_1 U7692 ( .ip1(i_i2c_prdata[21]), .ip2(i_ssi_prdata[21]), .s(n5616), 
        .op(n6531) );
  nand2_1 U7693 ( .ip1(n6676), .ip2(n6531), .op(n6535) );
  nand2_1 U7694 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[21]), .op(
        n6534) );
  nand2_1 U7695 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[21]), .op(n6533) );
  nand2_1 U7696 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[21]), .op(
        n6532) );
  mux2_1 U7697 ( .ip1(i_i2c_prdata[17]), .ip2(i_ssi_prdata[17]), .s(n5616), 
        .op(n6536) );
  nand2_1 U7698 ( .ip1(n6676), .ip2(n6536), .op(n6540) );
  nand2_1 U7699 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[17]), .op(
        n6539) );
  nand2_1 U7700 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[17]), .op(
        n6538) );
  nand2_1 U7701 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[17]), .op(n6537) );
  mux2_1 U7702 ( .ip1(i_i2c_prdata[29]), .ip2(i_ssi_prdata[29]), .s(n5616), 
        .op(n6541) );
  nand2_1 U7703 ( .ip1(n6676), .ip2(n6541), .op(n6545) );
  nand2_1 U7704 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[29]), .op(
        n6544) );
  nand2_1 U7705 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[29]), .op(
        n6543) );
  nand2_1 U7706 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[29]), .op(n6542) );
  mux2_1 U7707 ( .ip1(i_i2c_prdata[0]), .ip2(i_ssi_prdata[0]), .s(n5616), .op(
        n6546) );
  nand2_1 U7708 ( .ip1(n6676), .ip2(n6546), .op(n6550) );
  nand2_1 U7709 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[0]), .op(
        n6549) );
  nand2_1 U7710 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[0]), .op(
        n6548) );
  nand2_1 U7711 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[0]), .op(n6547) );
  mux2_1 U7712 ( .ip1(i_i2c_prdata[18]), .ip2(i_ssi_prdata[18]), .s(n5616), 
        .op(n6551) );
  nand2_1 U7713 ( .ip1(n6676), .ip2(n6551), .op(n6555) );
  nand2_1 U7714 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[18]), .op(
        n6554) );
  nand2_1 U7715 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[18]), .op(n6553) );
  nand2_1 U7716 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[18]), .op(
        n6552) );
  mux2_1 U7717 ( .ip1(i_i2c_prdata[24]), .ip2(i_ssi_prdata[24]), .s(n5616), 
        .op(n6556) );
  nand2_1 U7718 ( .ip1(n6676), .ip2(n6556), .op(n6560) );
  nand2_1 U7719 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[24]), .op(
        n6559) );
  nand2_1 U7720 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[24]), .op(n6558) );
  nand2_1 U7721 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[24]), .op(
        n6557) );
  mux2_1 U7722 ( .ip1(i_i2c_prdata[2]), .ip2(i_ssi_prdata[2]), .s(n5616), .op(
        n6561) );
  nand2_1 U7723 ( .ip1(n6676), .ip2(n6561), .op(n6565) );
  nand2_1 U7724 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[2]), .op(
        n6564) );
  nand2_1 U7725 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[2]), .op(
        n6563) );
  nand2_1 U7726 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[2]), .op(n6562) );
  mux2_1 U7727 ( .ip1(i_i2c_prdata[12]), .ip2(i_ssi_prdata[12]), .s(n5616), 
        .op(n6566) );
  nand2_1 U7728 ( .ip1(n6676), .ip2(n6566), .op(n6570) );
  nand2_1 U7729 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[12]), .op(
        n6569) );
  nand2_1 U7730 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[12]), .op(n6568) );
  nand2_1 U7731 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[12]), .op(
        n6567) );
  mux2_1 U7732 ( .ip1(i_i2c_prdata[28]), .ip2(i_ssi_prdata[28]), .s(n5617), 
        .op(n6571) );
  nand2_1 U7733 ( .ip1(n6676), .ip2(n6571), .op(n6575) );
  nand2_1 U7734 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[28]), .op(
        n6574) );
  nand2_1 U7735 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[28]), .op(
        n6573) );
  nand2_1 U7736 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[28]), .op(n6572) );
  mux2_1 U7737 ( .ip1(i_i2c_prdata[22]), .ip2(i_ssi_prdata[22]), .s(n5617), 
        .op(n6576) );
  nand2_1 U7738 ( .ip1(n6676), .ip2(n6576), .op(n6580) );
  nand2_1 U7739 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[22]), .op(
        n6579) );
  nand2_1 U7740 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[22]), .op(
        n6578) );
  nand2_1 U7741 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[22]), .op(n6577) );
  mux2_1 U7742 ( .ip1(i_i2c_prdata[4]), .ip2(i_ssi_prdata[4]), .s(n5616), .op(
        n6581) );
  nand2_1 U7743 ( .ip1(n6676), .ip2(n6581), .op(n6585) );
  nand2_1 U7744 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[4]), .op(
        n6584) );
  nand2_1 U7745 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[4]), .op(
        n6583) );
  nand2_1 U7746 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[4]), .op(n6582) );
  mux2_1 U7747 ( .ip1(i_i2c_prdata[19]), .ip2(i_ssi_prdata[19]), .s(n5617), 
        .op(n6586) );
  nand2_1 U7748 ( .ip1(n6676), .ip2(n6586), .op(n6590) );
  nand2_1 U7749 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[19]), .op(
        n6589) );
  nand2_1 U7750 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[19]), .op(n6588) );
  nand2_1 U7751 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[19]), .op(
        n6587) );
  mux2_1 U7752 ( .ip1(i_i2c_prdata[5]), .ip2(i_ssi_prdata[5]), .s(n5617), .op(
        n6591) );
  nand2_1 U7753 ( .ip1(n6676), .ip2(n6591), .op(n6595) );
  nand2_1 U7754 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[5]), .op(
        n6594) );
  nand2_1 U7755 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[5]), .op(n6593) );
  nand2_1 U7756 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[5]), .op(
        n6592) );
  mux2_1 U7757 ( .ip1(i_i2c_prdata[6]), .ip2(i_ssi_prdata[6]), .s(n5617), .op(
        n6596) );
  nand2_1 U7758 ( .ip1(n6676), .ip2(n6596), .op(n6600) );
  nand2_1 U7759 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[6]), .op(
        n6599) );
  nand2_1 U7760 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[6]), .op(
        n6598) );
  nand2_1 U7761 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[6]), .op(n6597) );
  mux2_1 U7762 ( .ip1(i_i2c_prdata[11]), .ip2(i_ssi_prdata[11]), .s(n5617), 
        .op(n6601) );
  nand2_1 U7763 ( .ip1(n6676), .ip2(n6601), .op(n6605) );
  nand2_1 U7764 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[11]), .op(
        n6604) );
  nand2_1 U7765 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[11]), .op(
        n6603) );
  nand2_1 U7766 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[11]), .op(n6602) );
  mux2_1 U7767 ( .ip1(i_i2c_prdata[3]), .ip2(i_ssi_prdata[3]), .s(n5617), .op(
        n6606) );
  nand2_1 U7768 ( .ip1(n6676), .ip2(n6606), .op(n6610) );
  nand2_1 U7769 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[3]), .op(
        n6609) );
  nand2_1 U7770 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[3]), .op(n6608) );
  nand2_1 U7771 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[3]), .op(
        n6607) );
  mux2_1 U7772 ( .ip1(i_i2c_prdata[7]), .ip2(i_ssi_prdata[7]), .s(n5617), .op(
        n6611) );
  nand2_1 U7773 ( .ip1(n6676), .ip2(n6611), .op(n6615) );
  nand2_1 U7774 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[7]), .op(
        n6614) );
  nand2_1 U7775 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[7]), .op(n6613) );
  nand2_1 U7776 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[7]), .op(
        n6612) );
  mux2_1 U7777 ( .ip1(i_i2c_prdata[26]), .ip2(i_ssi_prdata[26]), .s(n5617), 
        .op(n6616) );
  nand2_1 U7778 ( .ip1(n6676), .ip2(n6616), .op(n6620) );
  nand2_1 U7779 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[26]), .op(
        n6619) );
  nand2_1 U7780 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[26]), .op(
        n6618) );
  nand2_1 U7781 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[26]), .op(n6617) );
  mux2_1 U7782 ( .ip1(i_i2c_prdata[25]), .ip2(i_ssi_prdata[25]), .s(n5617), 
        .op(n6621) );
  nand2_1 U7783 ( .ip1(n6676), .ip2(n6621), .op(n6625) );
  nand2_1 U7784 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[25]), .op(
        n6624) );
  nand2_1 U7785 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[25]), .op(n6623) );
  nand2_1 U7786 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[25]), .op(
        n6622) );
  mux2_1 U7787 ( .ip1(i_i2c_prdata[16]), .ip2(i_ssi_prdata[16]), .s(n5617), 
        .op(n6626) );
  nand2_1 U7788 ( .ip1(n6676), .ip2(n6626), .op(n6630) );
  nand2_1 U7789 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[16]), .op(
        n6629) );
  nand2_1 U7790 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[16]), .op(n6628) );
  nand2_1 U7791 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[16]), .op(
        n6627) );
  mux2_1 U7792 ( .ip1(i_i2c_prdata[23]), .ip2(i_ssi_prdata[23]), .s(n5617), 
        .op(n6631) );
  nand2_1 U7793 ( .ip1(n6676), .ip2(n6631), .op(n6635) );
  nand2_1 U7794 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[23]), .op(
        n6634) );
  nand2_1 U7795 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[23]), .op(
        n6633) );
  nand2_1 U7796 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[23]), .op(n6632) );
  mux2_1 U7797 ( .ip1(i_i2c_prdata[14]), .ip2(i_ssi_prdata[14]), .s(n5617), 
        .op(n6636) );
  nand2_1 U7798 ( .ip1(n6676), .ip2(n6636), .op(n6640) );
  nand2_1 U7799 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[14]), .op(
        n6639) );
  nand2_1 U7800 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[14]), .op(n6638) );
  nand2_1 U7801 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[14]), .op(
        n6637) );
  mux2_1 U7802 ( .ip1(i_i2c_prdata[20]), .ip2(i_ssi_prdata[20]), .s(n5617), 
        .op(n6641) );
  nand2_1 U7803 ( .ip1(n6676), .ip2(n6641), .op(n6645) );
  nand2_1 U7804 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[20]), .op(
        n6644) );
  nand2_1 U7805 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[20]), .op(n6643) );
  nand2_1 U7806 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[20]), .op(
        n6642) );
  mux2_1 U7807 ( .ip1(i_i2c_prdata[10]), .ip2(i_ssi_prdata[10]), .s(n5617), 
        .op(n6646) );
  nand2_1 U7808 ( .ip1(n6676), .ip2(n6646), .op(n6650) );
  nand2_1 U7809 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[10]), .op(
        n6649) );
  nand2_1 U7810 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[10]), .op(n6648) );
  nand2_1 U7811 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[10]), .op(
        n6647) );
  mux2_1 U7812 ( .ip1(i_i2c_prdata[1]), .ip2(i_ssi_prdata[1]), .s(n5617), .op(
        n6651) );
  nand2_1 U7813 ( .ip1(n6676), .ip2(n6651), .op(n6655) );
  nand2_1 U7814 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[1]), .op(
        n6654) );
  nand2_1 U7815 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[1]), .op(
        n6653) );
  nand2_1 U7816 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[1]), .op(n6652) );
  mux2_1 U7817 ( .ip1(i_i2c_prdata[30]), .ip2(i_ssi_prdata[30]), .s(n5617), 
        .op(n6656) );
  nand2_1 U7818 ( .ip1(n6676), .ip2(n6656), .op(n6660) );
  nand2_1 U7819 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[30]), .op(
        n6659) );
  nand2_1 U7820 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[30]), .op(n6658) );
  nand2_1 U7821 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[30]), .op(
        n6657) );
  mux2_1 U7822 ( .ip1(i_i2c_prdata[15]), .ip2(i_ssi_prdata[15]), .s(n5617), 
        .op(n6661) );
  nand2_1 U7823 ( .ip1(n6676), .ip2(n6661), .op(n6665) );
  nand2_1 U7824 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[15]), .op(
        n6664) );
  nand2_1 U7825 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[15]), .op(
        n6663) );
  nand2_1 U7826 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[15]), .op(n6662) );
  mux2_1 U7827 ( .ip1(i_i2c_prdata[9]), .ip2(i_ssi_prdata[9]), .s(n5617), .op(
        n6666) );
  nand2_1 U7828 ( .ip1(n6676), .ip2(n6666), .op(n6670) );
  nand2_1 U7829 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[9]), .op(
        n6669) );
  nand2_1 U7830 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[9]), .op(n6668) );
  nand2_1 U7831 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[9]), .op(
        n6667) );
  mux2_1 U7832 ( .ip1(i_i2c_prdata[13]), .ip2(i_ssi_prdata[13]), .s(n5617), 
        .op(n6671) );
  nand2_1 U7833 ( .ip1(n6676), .ip2(n6671), .op(n6675) );
  nand2_1 U7834 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hrdata[13]), .op(
        n6674) );
  nand2_1 U7835 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hrdata[13]), .op(
        n6673) );
  nand2_1 U7836 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(
        ex_i_ahb_AHB_Slave_PID_hrdata[13]), .op(n6672) );
  nand2_1 U7837 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hready_resp), .op(
        n6682) );
  nand2_1 U7838 ( .ip1(n6676), .ip2(i_apb_hready_resp), .op(n6681) );
  nand2_1 U7839 ( .ip1(n6678), .ip2(n6677), .op(n6680) );
  nand2_1 U7840 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hready_resp), .op(
        n6679) );
  nand2_1 U7841 ( .ip1(i_ssi_reg_addr[1]), .ip2(i_ssi_reg_addr[2]), .op(n11463) );
  inv_1 U7842 ( .ip(i_ssi_reg_addr[3]), .op(n6684) );
  nand3_1 U7843 ( .ip1(n6685), .ip2(n6684), .ip3(i_ssi_reg_addr[4]), .op(
        n10752) );
  nor2_1 U7844 ( .ip1(n11463), .ip2(n10752), .op(n11661) );
  inv_1 U7845 ( .ip(n11661), .op(n11644) );
  inv_1 U7846 ( .ip(n6687), .op(n11663) );
  nor2_1 U7847 ( .ip1(n11644), .ip2(n11663), .op(n10081) );
  inv_1 U7848 ( .ip(i_ssi_reg_addr[0]), .op(n6807) );
  nand2_1 U7849 ( .ip1(n10081), .ip2(n6807), .op(n11665) );
  nand2_1 U7850 ( .ip1(n6687), .ip2(n11632), .op(n6688) );
  inv_1 U7851 ( .ip(i_ssi_rx_rd_addr[2]), .op(n6690) );
  nor3_1 U7852 ( .ip1(i_ssi_rx_rd_addr[1]), .ip2(i_ssi_rx_rd_addr[0]), .ip3(
        n6690), .op(n11614) );
  nand2_1 U7853 ( .ip1(n11614), .ip2(i_ssi_U_dff_rx_mem[58]), .op(n6701) );
  nand2_1 U7854 ( .ip1(i_ssi_rx_rd_addr[1]), .ip2(i_ssi_rx_rd_addr[0]), .op(
        n6936) );
  nor2_1 U7855 ( .ip1(i_ssi_rx_rd_addr[2]), .ip2(n6936), .op(n11618) );
  inv_1 U7856 ( .ip(i_ssi_rx_rd_addr[1]), .op(n6692) );
  nand3_1 U7857 ( .ip1(i_ssi_rx_rd_addr[2]), .ip2(i_ssi_rx_rd_addr[0]), .ip3(
        n6692), .op(n11616) );
  inv_1 U7858 ( .ip(i_ssi_U_dff_rx_mem[42]), .op(n6689) );
  nor2_1 U7859 ( .ip1(n11616), .ip2(n6689), .op(n6698) );
  nand2_1 U7860 ( .ip1(i_ssi_rx_rd_addr[1]), .ip2(i_ssi_rx_rd_addr[2]), .op(
        n10130) );
  nor2_1 U7861 ( .ip1(i_ssi_rx_rd_addr[0]), .ip2(n10130), .op(n11617) );
  nand2_1 U7862 ( .ip1(n11617), .ip2(i_ssi_U_dff_rx_mem[26]), .op(n6696) );
  nor2_1 U7863 ( .ip1(n6936), .ip2(n6690), .op(n11620) );
  nand2_1 U7864 ( .ip1(n11620), .ip2(i_ssi_U_dff_rx_mem[10]), .op(n6695) );
  inv_1 U7865 ( .ip(i_ssi_rx_rd_addr[0]), .op(n10127) );
  nand2_1 U7866 ( .ip1(n10127), .ip2(n6690), .op(n6691) );
  nor2_1 U7867 ( .ip1(i_ssi_rx_rd_addr[1]), .ip2(n6691), .op(n11627) );
  nand2_1 U7868 ( .ip1(n11627), .ip2(i_ssi_U_dff_rx_mem[122]), .op(n6694) );
  nor2_1 U7869 ( .ip1(n6692), .ip2(n6691), .op(n11628) );
  nand2_1 U7870 ( .ip1(n11628), .ip2(i_ssi_U_dff_rx_mem[90]), .op(n6693) );
  nand4_1 U7871 ( .ip1(n6696), .ip2(n6695), .ip3(n6694), .ip4(n6693), .op(
        n6697) );
  not_ab_or_c_or_d U7872 ( .ip1(i_ssi_U_dff_rx_mem[74]), .ip2(n11618), .ip3(
        n6698), .ip4(n6697), .op(n6700) );
  nor3_1 U7873 ( .ip1(i_ssi_rx_rd_addr[2]), .ip2(i_ssi_rx_rd_addr[1]), .ip3(
        n10127), .op(n11619) );
  nand2_1 U7874 ( .ip1(n11619), .ip2(i_ssi_U_dff_rx_mem[106]), .op(n6699) );
  nand3_1 U7875 ( .ip1(n6701), .ip2(n6700), .ip3(n6699), .op(n6702) );
  nand2_1 U7876 ( .ip1(n6937), .ip2(n6702), .op(n6713) );
  nand2_1 U7877 ( .ip1(n11663), .ip2(i_ssi_prdata[10]), .op(n6712) );
  nor2_1 U7878 ( .ip1(n6807), .ip2(n11644), .op(n6703) );
  nor2_1 U7879 ( .ip1(n6703), .ip2(n11663), .op(n11651) );
  nor2_1 U7880 ( .ip1(i_ssi_reg_addr[4]), .ip2(i_ssi_reg_addr[5]), .op(n6805)
         );
  nor2_1 U7881 ( .ip1(i_ssi_reg_addr[0]), .ip2(i_ssi_reg_addr[3]), .op(n6704)
         );
  and2_1 U7882 ( .ip1(n6805), .ip2(n6704), .op(n11469) );
  nor2_1 U7883 ( .ip1(i_ssi_reg_addr[1]), .ip2(i_ssi_reg_addr[2]), .op(n11481)
         );
  nand2_1 U7884 ( .ip1(n11469), .ip2(n11481), .op(n11470) );
  inv_1 U7885 ( .ip(n11470), .op(n11592) );
  nand2_1 U7886 ( .ip1(n11592), .ip2(i_ssi_ctrlr0[10]), .op(n6709) );
  inv_1 U7887 ( .ip(n11481), .op(n11485) );
  nor2_1 U7888 ( .ip1(i_ssi_reg_addr[3]), .ip2(n6807), .op(n6705) );
  nand2_1 U7889 ( .ip1(n6705), .ip2(n6805), .op(n10136) );
  nor2_1 U7890 ( .ip1(n11485), .ip2(n10136), .op(n11636) );
  nand2_1 U7891 ( .ip1(n11636), .ip2(i_ssi_U_regfile_ctrlr1_int[10]), .op(
        n6708) );
  inv_1 U7892 ( .ip(i_ssi_reg_addr[1]), .op(n6706) );
  and2_1 U7893 ( .ip1(n6706), .ip2(i_ssi_reg_addr[2]), .op(n11468) );
  inv_1 U7894 ( .ip(n11468), .op(n11603) );
  nor2_1 U7895 ( .ip1(n10136), .ip2(n11603), .op(n11635) );
  nand2_1 U7896 ( .ip1(n11635), .ip2(i_ssi_baudr[10]), .op(n6707) );
  nand3_1 U7897 ( .ip1(n6709), .ip2(n6708), .ip3(n6707), .op(n6710) );
  nand2_1 U7898 ( .ip1(n11651), .ip2(n6710), .op(n6711) );
  nand4_1 U7899 ( .ip1(n11665), .ip2(n6713), .ip3(n6712), .ip4(n6711), .op(
        n4227) );
  nand2_1 U7900 ( .ip1(n11663), .ip2(i_ssi_prdata[11]), .op(n6731) );
  nand2_1 U7901 ( .ip1(n11592), .ip2(i_ssi_ctrlr0[11]), .op(n6716) );
  nand2_1 U7902 ( .ip1(n11636), .ip2(n5391), .op(n6715) );
  nand2_1 U7903 ( .ip1(n11635), .ip2(i_ssi_baudr[11]), .op(n6714) );
  nand3_1 U7904 ( .ip1(n6716), .ip2(n6715), .ip3(n6714), .op(n6717) );
  nand2_1 U7905 ( .ip1(n11651), .ip2(n6717), .op(n6730) );
  nand2_1 U7906 ( .ip1(n11617), .ip2(i_ssi_U_dff_rx_mem[27]), .op(n6727) );
  inv_1 U7907 ( .ip(i_ssi_U_dff_rx_mem[43]), .op(n6718) );
  nor2_1 U7908 ( .ip1(n11616), .ip2(n6718), .op(n6724) );
  nand2_1 U7909 ( .ip1(n11619), .ip2(i_ssi_U_dff_rx_mem[107]), .op(n6722) );
  nand2_1 U7910 ( .ip1(n11614), .ip2(i_ssi_U_dff_rx_mem[59]), .op(n6721) );
  nand2_1 U7911 ( .ip1(n11618), .ip2(i_ssi_U_dff_rx_mem[75]), .op(n6720) );
  nand2_1 U7912 ( .ip1(n11620), .ip2(i_ssi_U_dff_rx_mem[11]), .op(n6719) );
  nand4_1 U7913 ( .ip1(n6722), .ip2(n6721), .ip3(n6720), .ip4(n6719), .op(
        n6723) );
  not_ab_or_c_or_d U7914 ( .ip1(i_ssi_U_dff_rx_mem[91]), .ip2(n11628), .ip3(
        n6724), .ip4(n6723), .op(n6726) );
  nand2_1 U7915 ( .ip1(n11627), .ip2(i_ssi_U_dff_rx_mem[123]), .op(n6725) );
  nand3_1 U7916 ( .ip1(n6727), .ip2(n6726), .ip3(n6725), .op(n6728) );
  nand2_1 U7917 ( .ip1(n6937), .ip2(n6728), .op(n6729) );
  nand4_1 U7918 ( .ip1(n11665), .ip2(n6731), .ip3(n6730), .ip4(n6729), .op(
        n4226) );
  nand2_1 U7919 ( .ip1(n11663), .ip2(i_ssi_prdata[15]), .op(n6749) );
  nand2_1 U7920 ( .ip1(n11592), .ip2(i_ssi_cfs[3]), .op(n6734) );
  nand2_1 U7921 ( .ip1(n11636), .ip2(n5434), .op(n6733) );
  nand2_1 U7922 ( .ip1(n11635), .ip2(i_ssi_baudr[15]), .op(n6732) );
  nand3_1 U7923 ( .ip1(n6734), .ip2(n6733), .ip3(n6732), .op(n6735) );
  nand2_1 U7924 ( .ip1(n11651), .ip2(n6735), .op(n6748) );
  nand2_1 U7925 ( .ip1(n11617), .ip2(i_ssi_U_dff_rx_mem[31]), .op(n6745) );
  inv_1 U7926 ( .ip(i_ssi_U_dff_rx_mem[47]), .op(n6736) );
  nor2_1 U7927 ( .ip1(n11616), .ip2(n6736), .op(n6742) );
  nand2_1 U7928 ( .ip1(n11628), .ip2(i_ssi_U_dff_rx_mem[95]), .op(n6740) );
  nand2_1 U7929 ( .ip1(n11627), .ip2(i_ssi_U_dff_rx_mem[127]), .op(n6739) );
  nand2_1 U7930 ( .ip1(n11619), .ip2(i_ssi_U_dff_rx_mem[111]), .op(n6738) );
  nand2_1 U7931 ( .ip1(n11614), .ip2(i_ssi_U_dff_rx_mem[63]), .op(n6737) );
  nand4_1 U7932 ( .ip1(n6740), .ip2(n6739), .ip3(n6738), .ip4(n6737), .op(
        n6741) );
  not_ab_or_c_or_d U7933 ( .ip1(i_ssi_U_dff_rx_mem[15]), .ip2(n11620), .ip3(
        n6742), .ip4(n6741), .op(n6744) );
  nand2_1 U7934 ( .ip1(n11618), .ip2(i_ssi_U_dff_rx_mem[79]), .op(n6743) );
  nand3_1 U7935 ( .ip1(n6745), .ip2(n6744), .ip3(n6743), .op(n6746) );
  nand2_1 U7936 ( .ip1(n6937), .ip2(n6746), .op(n6747) );
  nand4_1 U7937 ( .ip1(n11665), .ip2(n6749), .ip3(n6748), .ip4(n6747), .op(
        n4222) );
  nand2_1 U7938 ( .ip1(n11663), .ip2(i_ssi_prdata[7]), .op(n6766) );
  nand2_1 U7939 ( .ip1(n11635), .ip2(i_ssi_baudr[7]), .op(n6751) );
  nand2_1 U7940 ( .ip1(n11636), .ip2(i_ssi_U_regfile_ctrlr1_int[7]), .op(n6750) );
  nand2_1 U7941 ( .ip1(n6751), .ip2(n6750), .op(n6752) );
  nand2_1 U7942 ( .ip1(n11651), .ip2(n6752), .op(n6765) );
  nand2_1 U7943 ( .ip1(n11628), .ip2(i_ssi_U_dff_rx_mem[87]), .op(n6762) );
  inv_1 U7944 ( .ip(i_ssi_U_dff_rx_mem[39]), .op(n6753) );
  nor2_1 U7945 ( .ip1(n11616), .ip2(n6753), .op(n6759) );
  nand2_1 U7946 ( .ip1(n11617), .ip2(i_ssi_U_dff_rx_mem[23]), .op(n6757) );
  nand2_1 U7947 ( .ip1(n11620), .ip2(i_ssi_U_dff_rx_mem[7]), .op(n6756) );
  nand2_1 U7948 ( .ip1(n11614), .ip2(i_ssi_U_dff_rx_mem[55]), .op(n6755) );
  nand2_1 U7949 ( .ip1(n11618), .ip2(i_ssi_U_dff_rx_mem[71]), .op(n6754) );
  nand4_1 U7950 ( .ip1(n6757), .ip2(n6756), .ip3(n6755), .ip4(n6754), .op(
        n6758) );
  not_ab_or_c_or_d U7951 ( .ip1(i_ssi_U_dff_rx_mem[119]), .ip2(n11627), .ip3(
        n6759), .ip4(n6758), .op(n6761) );
  nand2_1 U7952 ( .ip1(n11619), .ip2(i_ssi_U_dff_rx_mem[103]), .op(n6760) );
  nand3_1 U7953 ( .ip1(n6762), .ip2(n6761), .ip3(n6760), .op(n6763) );
  nand2_1 U7954 ( .ip1(n6937), .ip2(n6763), .op(n6764) );
  nand4_1 U7955 ( .ip1(n11665), .ip2(n6766), .ip3(n6765), .ip4(n6764), .op(
        n4230) );
  nand2_1 U7956 ( .ip1(n11663), .ip2(i_ssi_prdata[14]), .op(n6784) );
  nand2_1 U7957 ( .ip1(n11592), .ip2(i_ssi_cfs[2]), .op(n6769) );
  nand2_1 U7958 ( .ip1(n11636), .ip2(i_ssi_U_regfile_ctrlr1_int[14]), .op(
        n6768) );
  nand2_1 U7959 ( .ip1(n11635), .ip2(i_ssi_baudr[14]), .op(n6767) );
  nand3_1 U7960 ( .ip1(n6769), .ip2(n6768), .ip3(n6767), .op(n6770) );
  nand2_1 U7961 ( .ip1(n11651), .ip2(n6770), .op(n6783) );
  nand2_1 U7962 ( .ip1(n11614), .ip2(i_ssi_U_dff_rx_mem[62]), .op(n6780) );
  inv_1 U7963 ( .ip(i_ssi_U_dff_rx_mem[46]), .op(n6771) );
  nor2_1 U7964 ( .ip1(n11616), .ip2(n6771), .op(n6777) );
  nand2_1 U7965 ( .ip1(n11628), .ip2(i_ssi_U_dff_rx_mem[94]), .op(n6775) );
  nand2_1 U7966 ( .ip1(n11617), .ip2(i_ssi_U_dff_rx_mem[30]), .op(n6774) );
  nand2_1 U7967 ( .ip1(n11619), .ip2(i_ssi_U_dff_rx_mem[110]), .op(n6773) );
  nand2_1 U7968 ( .ip1(n11620), .ip2(i_ssi_U_dff_rx_mem[14]), .op(n6772) );
  nand4_1 U7969 ( .ip1(n6775), .ip2(n6774), .ip3(n6773), .ip4(n6772), .op(
        n6776) );
  not_ab_or_c_or_d U7970 ( .ip1(i_ssi_U_dff_rx_mem[78]), .ip2(n11618), .ip3(
        n6777), .ip4(n6776), .op(n6779) );
  nand2_1 U7971 ( .ip1(n11627), .ip2(i_ssi_U_dff_rx_mem[126]), .op(n6778) );
  nand3_1 U7972 ( .ip1(n6780), .ip2(n6779), .ip3(n6778), .op(n6781) );
  nand2_1 U7973 ( .ip1(n6937), .ip2(n6781), .op(n6782) );
  nand4_1 U7974 ( .ip1(n11665), .ip2(n6784), .ip3(n6783), .ip4(n6782), .op(
        n4223) );
  nand2_1 U7975 ( .ip1(n11663), .ip2(i_ssi_prdata[6]), .op(n6803) );
  nand2_1 U7976 ( .ip1(n6805), .ip2(i_ssi_reg_addr[3]), .op(n11609) );
  nor2_1 U7977 ( .ip1(i_ssi_reg_addr[0]), .ip2(n11609), .op(n11482) );
  inv_1 U7978 ( .ip(i_ssi_reg_addr[2]), .op(n6785) );
  and2_1 U7979 ( .ip1(n6785), .ip2(i_ssi_reg_addr[1]), .op(n6816) );
  and2_1 U7980 ( .ip1(n11482), .ip2(n6816), .op(n11647) );
  nand2_1 U7981 ( .ip1(n11647), .ip2(i_ssi_U_regfile_sr_6_), .op(n6788) );
  nand2_1 U7982 ( .ip1(n11635), .ip2(i_ssi_baudr[6]), .op(n6787) );
  nand2_1 U7983 ( .ip1(n11636), .ip2(i_ssi_U_regfile_ctrlr1_int[6]), .op(n6786) );
  nand3_1 U7984 ( .ip1(n6788), .ip2(n6787), .ip3(n6786), .op(n6789) );
  nand2_1 U7985 ( .ip1(n11651), .ip2(n6789), .op(n6802) );
  nand2_1 U7986 ( .ip1(n11618), .ip2(i_ssi_U_dff_rx_mem[70]), .op(n6799) );
  inv_1 U7987 ( .ip(i_ssi_U_dff_rx_mem[38]), .op(n6790) );
  nor2_1 U7988 ( .ip1(n11616), .ip2(n6790), .op(n6796) );
  nand2_1 U7989 ( .ip1(n11627), .ip2(i_ssi_U_dff_rx_mem[118]), .op(n6794) );
  nand2_1 U7990 ( .ip1(n11619), .ip2(i_ssi_U_dff_rx_mem[102]), .op(n6793) );
  nand2_1 U7991 ( .ip1(n11620), .ip2(i_ssi_U_dff_rx_mem[6]), .op(n6792) );
  nand2_1 U7992 ( .ip1(n11617), .ip2(i_ssi_U_dff_rx_mem[22]), .op(n6791) );
  nand4_1 U7993 ( .ip1(n6794), .ip2(n6793), .ip3(n6792), .ip4(n6791), .op(
        n6795) );
  not_ab_or_c_or_d U7994 ( .ip1(i_ssi_U_dff_rx_mem[54]), .ip2(n11614), .ip3(
        n6796), .ip4(n6795), .op(n6798) );
  nand2_1 U7995 ( .ip1(n11628), .ip2(i_ssi_U_dff_rx_mem[86]), .op(n6797) );
  nand3_1 U7996 ( .ip1(n6799), .ip2(n6798), .ip3(n6797), .op(n6800) );
  nand2_1 U7997 ( .ip1(n6937), .ip2(n6800), .op(n6801) );
  nand4_1 U7998 ( .ip1(n11665), .ip2(n6803), .ip3(n6802), .ip4(n6801), .op(
        n4231) );
  and2_1 U7999 ( .ip1(i_ssi_reg_addr[3]), .ip2(i_ssi_reg_addr[0]), .op(n6804)
         );
  nand2_1 U8000 ( .ip1(n6805), .ip2(n6804), .op(n11484) );
  inv_1 U8001 ( .ip(n6816), .op(n9810) );
  nor2_1 U8002 ( .ip1(n11484), .ip2(n9810), .op(n11640) );
  inv_1 U8003 ( .ip(n11640), .op(n10005) );
  nor2_1 U8004 ( .ip1(n10005), .ip2(n10139), .op(n10846) );
  inv_1 U8005 ( .ip(n10846), .op(n6806) );
  nor2_1 U8006 ( .ip1(i_apb_pwdata_int[5]), .ip2(n6806), .op(n9702) );
  xor2_1 U8007 ( .ip1(i_ssi_U_regfile_multi_mst_edge), .ip2(
        i_ssi_fsm_multi_mst), .op(n10015) );
  nor2_1 U8008 ( .ip1(i_ssi_risr[5]), .ip2(n10015), .op(n6812) );
  or2_1 U8009 ( .ip1(i_ssi_imr[5]), .ip2(n10846), .op(n9700) );
  nand2_1 U8010 ( .ip1(n6816), .ip2(n6807), .op(n6808) );
  nor2_1 U8011 ( .ip1(n10752), .ip2(n6808), .op(n11467) );
  inv_1 U8012 ( .ip(n11467), .op(n10760) );
  nor2_1 U8013 ( .ip1(n11485), .ip2(n10752), .op(n11457) );
  nand2_1 U8014 ( .ip1(n11457), .ip2(i_ssi_reg_addr[0]), .op(n6809) );
  and2_1 U8015 ( .ip1(n10760), .ip2(n6809), .op(n11462) );
  or2_1 U8016 ( .ip1(n11462), .ip2(n11663), .op(n9991) );
  and3_1 U8017 ( .ip1(n9991), .ip2(i_ssi_risr[5]), .ip3(i_ssi_mst_contention), 
        .op(n6810) );
  nor2_1 U8018 ( .ip1(n9700), .ip2(n6810), .op(n6811) );
  nor4_1 U8019 ( .ip1(n9702), .ip2(n6812), .ip3(n5291), .ip4(n6811), .op(n4239) );
  and2_1 U8020 ( .ip1(n11854), .ip2(n5588), .op(n10758) );
  nand2_1 U8021 ( .ip1(i_ssi_U_fifo_U_tx_fifo_empty_n), .ip2(i_ssi_tx_full), 
        .op(n6813) );
  nand2_1 U8022 ( .ip1(n10758), .ip2(n6813), .op(n9921) );
  or2_1 U8023 ( .ip1(n5588), .ip2(n11854), .op(n9926) );
  nand2_1 U8024 ( .ip1(n9921), .ip2(n9926), .op(n6814) );
  xnor2_1 U8025 ( .ip1(i_ssi_U_fifo_unconnected_tx_wrd_count[0]), .ip2(n6814), 
        .op(n6815) );
  inv_1 U8026 ( .ip(n6815), .op(n6819) );
  nand2_1 U8027 ( .ip1(n11469), .ip2(n6816), .op(n11475) );
  nor2_1 U8028 ( .ip1(n11475), .ip2(n10139), .op(n9699) );
  inv_1 U8029 ( .ip(i_apb_pwdata_int[0]), .op(n6817) );
  nand2_1 U8030 ( .ip1(n9699), .ip2(n6817), .op(n6818) );
  and2_1 U8031 ( .ip1(n6818), .ip2(n10802), .op(n10759) );
  and2_1 U8032 ( .ip1(n6819), .ip2(n10759), .op(n11853) );
  inv_1 U8033 ( .ip(i_apb_U_DW_apb_ahbsif_pipeline_c), .op(n10094) );
  or2_1 U8034 ( .ip1(i_apb_U_DW_apb_ahbsif_state[1]), .ip2(
        i_apb_U_DW_apb_ahbsif_state[0]), .op(n6849) );
  inv_1 U8035 ( .ip(n6849), .op(n10105) );
  nand2_1 U8036 ( .ip1(n10105), .ip2(i_apb_U_DW_apb_ahbsif_state[2]), .op(
        n6859) );
  nor2_1 U8037 ( .ip1(n10094), .ip2(n6859), .op(n6829) );
  and2_1 U8038 ( .ip1(i_apb_U_DW_apb_ahbsif_state[0]), .ip2(
        i_apb_U_DW_apb_ahbsif_state[1]), .op(n7416) );
  inv_1 U8039 ( .ip(i_apb_U_DW_apb_ahbsif_state[2]), .op(n10098) );
  nand2_1 U8040 ( .ip1(n7416), .ip2(n10098), .op(n7428) );
  inv_1 U8041 ( .ip(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[14]), .op(n6821) );
  inv_1 U8042 ( .ip(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[15]), .op(n6820) );
  nand3_1 U8043 ( .ip1(n6821), .ip2(n6820), .ip3(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[16]), .op(n6827) );
  nor4_1 U8044 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[29]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[28]), .ip3(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[25]), .ip4(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[24]), .op(n6824) );
  nor4_1 U8045 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[21]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[20]), .ip3(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[19]), .ip4(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[18]), .op(n6823) );
  nor4_1 U8046 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[17]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[23]), .ip3(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[26]), .ip4(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[22]), .op(n6822) );
  nor3_1 U8047 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[31]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[27]), .ip3(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[30]), .op(n6826) );
  nand2_1 U8048 ( .ip1(n6825), .ip2(n6826), .op(n11158) );
  inv_1 U8049 ( .ip(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[13]), .op(n9661) );
  and3_1 U8050 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_hready), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_htrans[1]), .ip3(n9661), .op(n6828) );
  inv_1 U8051 ( .ip(n7413), .op(n7405) );
  nor2_1 U8052 ( .ip1(n7428), .ip2(n7405), .op(n7418) );
  nor2_1 U8053 ( .ip1(n6829), .ip2(n7418), .op(n6837) );
  inv_1 U8054 ( .ip(i_apb_pclk_en), .op(n10100) );
  inv_1 U8055 ( .ip(i_apb_U_DW_apb_ahbsif_state[0]), .op(n10099) );
  nand3_1 U8056 ( .ip1(n10099), .ip2(i_apb_U_DW_apb_ahbsif_state[1]), .ip3(
        i_apb_U_DW_apb_ahbsif_state[2]), .op(n7173) );
  nand2_1 U8057 ( .ip1(n7428), .ip2(n7173), .op(n10083) );
  nand2_1 U8058 ( .ip1(n10083), .ip2(n10094), .op(n6841) );
  ab_or_c_or_d U8059 ( .ip1(n6849), .ip2(n6841), .ip3(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite), .ip4(n7413), .op(n6833) );
  nor2_1 U8060 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_hwrite_c), .ip2(n10094), 
        .op(n6830) );
  nand2_1 U8061 ( .ip1(n10083), .ip2(n6830), .op(n6843) );
  inv_1 U8062 ( .ip(i_apb_U_DW_apb_ahbsif_state[1]), .op(n10101) );
  nand2_1 U8063 ( .ip1(n10101), .ip2(i_apb_U_DW_apb_ahbsif_state[2]), .op(
        n6831) );
  and2_1 U8064 ( .ip1(n6843), .ip2(n6831), .op(n6832) );
  nand2_1 U8065 ( .ip1(n6833), .ip2(n6832), .op(
        i_apb_U_DW_apb_ahbsif_nextstate[2]) );
  inv_1 U8066 ( .ip(i_apb_U_DW_apb_ahbsif_nextstate[2]), .op(n10087) );
  and2_1 U8067 ( .ip1(i_apb_U_DW_apb_ahbsif_pipeline_c), .ip2(
        i_apb_U_DW_apb_ahbsif_piped_hwrite_c), .op(n6834) );
  nand2_1 U8068 ( .ip1(n10083), .ip2(n6834), .op(n6844) );
  nand2_1 U8069 ( .ip1(n10101), .ip2(i_apb_U_DW_apb_ahbsif_state[0]), .op(
        n7408) );
  nand2_1 U8070 ( .ip1(n6844), .ip2(n7408), .op(n6835) );
  nand2_1 U8071 ( .ip1(i_apb_pclk_en), .ip2(n6835), .op(n6836) );
  nand3_1 U8072 ( .ip1(n10099), .ip2(n10098), .ip3(
        i_apb_U_DW_apb_ahbsif_state[1]), .op(n9609) );
  nand2_1 U8073 ( .ip1(n6836), .ip2(n9609), .op(
        i_apb_U_DW_apb_ahbsif_nextstate[1]) );
  or2_1 U8074 ( .ip1(n10087), .ip2(i_apb_U_DW_apb_ahbsif_nextstate[1]), .op(
        n9607) );
  or2_1 U8075 ( .ip1(n10100), .ip2(n9607), .op(n9611) );
  nor2_1 U8076 ( .ip1(n6837), .ip2(n9611), .op(n6855) );
  nand2_1 U8077 ( .ip1(i_apb_U_DW_apb_ahbsif_nextstate[1]), .ip2(n10087), .op(
        n6853) );
  inv_1 U8078 ( .ip(n7408), .op(n9684) );
  nor2_1 U8079 ( .ip1(n9684), .ip2(i_apb_pclk_en), .op(n6840) );
  inv_1 U8080 ( .ip(n9609), .op(n6838) );
  nand2_1 U8081 ( .ip1(i_apb_pclk_en), .ip2(n6859), .op(n6856) );
  nor2_1 U8082 ( .ip1(n6838), .ip2(n6856), .op(n6839) );
  nor2_1 U8083 ( .ip1(n6840), .ip2(n6839), .op(n6848) );
  or2_1 U8084 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite), .ip2(i_apb_pclk_en), 
        .op(n6851) );
  nor2_1 U8085 ( .ip1(n6841), .ip2(n7413), .op(n6842) );
  nand2_1 U8086 ( .ip1(n6851), .ip2(n6842), .op(n6846) );
  mux2_1 U8087 ( .ip1(n6844), .ip2(n6843), .s(i_apb_pclk_en), .op(n6845) );
  nand2_1 U8088 ( .ip1(n6846), .ip2(n6845), .op(n6847) );
  or2_1 U8089 ( .ip1(i_apb_U_DW_apb_ahbsif_state[2]), .ip2(n6849), .op(n10085)
         );
  nor2_1 U8090 ( .ip1(n10085), .ip2(n7413), .op(n6850) );
  nand2_1 U8091 ( .ip1(n6851), .ip2(n6850), .op(n6852) );
  nand2_1 U8092 ( .ip1(n10091), .ip2(i_apb_pclk_en), .op(n6857) );
  nor2_1 U8093 ( .ip1(i_apb_U_DW_apb_ahbsif_use_saved_c), .ip2(n11117), .op(
        n6854) );
  or2_1 U8094 ( .ip1(n6855), .ip2(n6854), .op(n6892) );
  nand2_1 U8095 ( .ip1(n6892), .ip2(i_apb_U_DW_apb_ahbsif_piped_haddr_c[4]), 
        .op(n6867) );
  nor3_1 U8096 ( .ip1(n7418), .ip2(n6856), .ip3(n9607), .op(n7266) );
  nand2_1 U8097 ( .ip1(n7239), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[4]), 
        .op(n6866) );
  inv_1 U8098 ( .ip(n9611), .op(n6861) );
  inv_1 U8099 ( .ip(n6857), .op(n6858) );
  nand2_1 U8100 ( .ip1(n5249), .ip2(i_ssi_reg_addr[2]), .op(n6865) );
  nand2_1 U8101 ( .ip1(n6858), .ip2(i_apb_U_DW_apb_ahbsif_use_saved_c), .op(
        n6863) );
  inv_1 U8102 ( .ip(n6859), .op(n6860) );
  nand3_1 U8103 ( .ip1(n6861), .ip2(n6860), .ip3(n10094), .op(n6862) );
  nand2_1 U8104 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[4]), 
        .op(n6864) );
  nand4_1 U8105 ( .ip1(n6867), .ip2(n6866), .ip3(n6865), .ip4(n6864), .op(
        n4724) );
  nand2_1 U8106 ( .ip1(n6892), .ip2(i_apb_U_DW_apb_ahbsif_piped_haddr_c[7]), 
        .op(n6871) );
  nand2_1 U8107 ( .ip1(n7239), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[7]), 
        .op(n6870) );
  nand2_1 U8108 ( .ip1(n5249), .ip2(i_ssi_reg_addr[5]), .op(n6869) );
  nand2_1 U8109 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[7]), 
        .op(n6868) );
  nand4_1 U8110 ( .ip1(n6871), .ip2(n6870), .ip3(n6869), .ip4(n6868), .op(
        n4721) );
  nand2_1 U8111 ( .ip1(n6892), .ip2(i_apb_U_DW_apb_ahbsif_piped_haddr_c[16]), 
        .op(n6875) );
  nand2_1 U8112 ( .ip1(n7239), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[16]), 
        .op(n6874) );
  nand2_1 U8113 ( .ip1(n5249), .ip2(i_apb_paddr[16]), .op(n6873) );
  nand2_1 U8114 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[16]), 
        .op(n6872) );
  nand4_1 U8115 ( .ip1(n6875), .ip2(n6874), .ip3(n6873), .ip4(n6872), .op(
        n4716) );
  nand2_1 U8116 ( .ip1(n6892), .ip2(i_apb_U_DW_apb_ahbsif_piped_haddr_c[5]), 
        .op(n6879) );
  nand2_1 U8117 ( .ip1(n7239), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[5]), 
        .op(n6878) );
  nand2_1 U8118 ( .ip1(n5249), .ip2(i_ssi_reg_addr[3]), .op(n6877) );
  nand2_1 U8119 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[5]), 
        .op(n6876) );
  nand4_1 U8120 ( .ip1(n6879), .ip2(n6878), .ip3(n6877), .ip4(n6876), .op(
        n4723) );
  nand2_1 U8121 ( .ip1(n6892), .ip2(i_apb_U_DW_apb_ahbsif_piped_haddr_c[6]), 
        .op(n6883) );
  nand2_1 U8122 ( .ip1(n7239), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[6]), 
        .op(n6882) );
  nand2_1 U8123 ( .ip1(n5249), .ip2(i_ssi_reg_addr[4]), .op(n6881) );
  nand2_1 U8124 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[6]), 
        .op(n6880) );
  nand4_1 U8125 ( .ip1(n6883), .ip2(n6882), .ip3(n6881), .ip4(n6880), .op(
        n4722) );
  nand2_1 U8126 ( .ip1(n6892), .ip2(i_apb_U_DW_apb_ahbsif_piped_haddr_c[3]), 
        .op(n6887) );
  nand2_1 U8127 ( .ip1(n7239), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[3]), 
        .op(n6886) );
  nand2_1 U8128 ( .ip1(n5249), .ip2(i_ssi_reg_addr[1]), .op(n6885) );
  nand2_1 U8129 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[3]), 
        .op(n6884) );
  nand4_1 U8130 ( .ip1(n6887), .ip2(n6886), .ip3(n6885), .ip4(n6884), .op(
        n4725) );
  nand2_1 U8131 ( .ip1(n6892), .ip2(i_apb_U_DW_apb_ahbsif_piped_haddr_c[12]), 
        .op(n6891) );
  nand2_1 U8132 ( .ip1(n7239), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[12]), 
        .op(n6890) );
  nand2_1 U8133 ( .ip1(n5249), .ip2(i_apb_paddr[12]), .op(n6889) );
  nand2_1 U8134 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[12]), 
        .op(n6888) );
  nand4_1 U8135 ( .ip1(n6891), .ip2(n6890), .ip3(n6889), .ip4(n6888), .op(
        n4720) );
  nand2_1 U8136 ( .ip1(n6892), .ip2(i_apb_U_DW_apb_ahbsif_piped_haddr_c[2]), 
        .op(n6896) );
  nand2_1 U8137 ( .ip1(n7239), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[2]), 
        .op(n6895) );
  nand2_1 U8138 ( .ip1(n5249), .ip2(i_ssi_reg_addr[0]), .op(n6894) );
  nand2_1 U8139 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[2]), 
        .op(n6893) );
  nand4_1 U8140 ( .ip1(n6896), .ip2(n6895), .ip3(n6894), .ip4(n6893), .op(
        n4726) );
  inv_1 U8141 ( .ip(i_ssi_U_fifo_unconnected_rx_wrd_count[2]), .op(n6903) );
  nand2_1 U8142 ( .ip1(i_ssi_U_fifo_U_rx_fifo_empty_n), .ip2(n6937), .op(
        n10128) );
  inv_1 U8143 ( .ip(i_ssi_U_fifo_rx_push_edge), .op(n6897) );
  nand2_1 U8144 ( .ip1(i_ssi_U_fifo_U_rx_fifo_empty_n), .ip2(i_ssi_rx_full), 
        .op(n6898) );
  and2_1 U8145 ( .ip1(n11837), .ip2(n6898), .op(n6899) );
  nand2_1 U8146 ( .ip1(n10128), .ip2(n6899), .op(n6909) );
  nand2_1 U8147 ( .ip1(i_ssi_U_fifo_unconnected_rx_wrd_count[0]), .ip2(n6909), 
        .op(n6917) );
  inv_1 U8148 ( .ip(n10128), .op(n10749) );
  nand2_1 U8149 ( .ip1(n10749), .ip2(n10713), .op(n6915) );
  inv_1 U8150 ( .ip(n6915), .op(n6900) );
  mux2_1 U8151 ( .ip1(n6900), .ip2(i_ssi_U_fifo_unconnected_rx_wrd_count[0]), 
        .s(i_ssi_U_fifo_unconnected_rx_wrd_count[1]), .op(n6901) );
  nand2_1 U8152 ( .ip1(n6917), .ip2(n6901), .op(n6902) );
  xnor2_1 U8153 ( .ip1(n6903), .ip2(n6902), .op(n6904) );
  inv_1 U8154 ( .ip(n6904), .op(n6905) );
  and2_1 U8155 ( .ip1(n6905), .ip2(n10759), .op(n11850) );
  nand3_1 U8156 ( .ip1(i_ssi_U_fifo_unconnected_rx_wrd_count[2]), .ip2(
        i_ssi_U_fifo_unconnected_rx_wrd_count[1]), .ip3(
        i_ssi_U_fifo_unconnected_rx_wrd_count[0]), .op(n6906) );
  nor3_1 U8157 ( .ip1(n10713), .ip2(n6906), .ip3(n6937), .op(n6907) );
  nor2_1 U8158 ( .ip1(i_ssi_rx_full), .ip2(n6907), .op(n6908) );
  inv_1 U8159 ( .ip(n10759), .op(n10748) );
  not_ab_or_c_or_d U8160 ( .ip1(n6937), .ip2(n10713), .ip3(n6908), .ip4(n10748), .op(n11871) );
  inv_1 U8161 ( .ip(i_ssi_rxftlr[2]), .op(n10848) );
  nand2_1 U8162 ( .ip1(n6915), .ip2(n6909), .op(n6911) );
  inv_1 U8163 ( .ip(n6911), .op(n6910) );
  nand2_1 U8164 ( .ip1(n6910), .ip2(i_ssi_U_fifo_unconnected_rx_wrd_count[0]), 
        .op(n6913) );
  inv_1 U8165 ( .ip(i_ssi_U_fifo_unconnected_rx_wrd_count[0]), .op(n6914) );
  nand2_1 U8166 ( .ip1(n6911), .ip2(n6914), .op(n6912) );
  and2_1 U8167 ( .ip1(n6913), .ip2(n6912), .op(n10123) );
  nor3_1 U8168 ( .ip1(n10123), .ip2(i_ssi_rxftlr[0]), .ip3(i_ssi_rxftlr[1]), 
        .op(n6921) );
  inv_1 U8169 ( .ip(i_ssi_U_fifo_unconnected_rx_wrd_count[1]), .op(n6919) );
  nand2_1 U8170 ( .ip1(n6915), .ip2(n6914), .op(n6916) );
  nand2_1 U8171 ( .ip1(n6917), .ip2(n6916), .op(n6918) );
  xnor2_1 U8172 ( .ip1(n6919), .ip2(n6918), .op(n6920) );
  inv_1 U8173 ( .ip(n6920), .op(n10124) );
  nor2_1 U8174 ( .ip1(n6921), .ip2(n10124), .op(n6924) );
  nand2_1 U8175 ( .ip1(i_ssi_rxftlr[0]), .ip2(i_ssi_rxftlr[1]), .op(n10847) );
  and3_1 U8176 ( .ip1(n10759), .ip2(n10848), .ip3(n10847), .op(n6922) );
  nor2_1 U8177 ( .ip1(n6922), .ip2(n11850), .op(n6923) );
  not_ab_or_c_or_d U8178 ( .ip1(i_ssi_rxftlr[1]), .ip2(n10123), .ip3(n6924), 
        .ip4(n6923), .op(n6925) );
  ab_or_c_or_d U8179 ( .ip1(n11850), .ip2(n10848), .ip3(n6925), .ip4(n11871), 
        .op(n11830) );
  xor2_1 U8180 ( .ip1(i_ssi_cfs[3]), .ip2(i_ssi_U_mstfsm_ctrl_cnt[3]), .op(
        n6927) );
  xor2_1 U8181 ( .ip1(i_ssi_cfs[2]), .ip2(i_ssi_U_mstfsm_ctrl_cnt[2]), .op(
        n6926) );
  nor2_1 U8182 ( .ip1(n6927), .ip2(n6926), .op(n6931) );
  xor2_1 U8183 ( .ip1(i_ssi_cfs[0]), .ip2(i_ssi_U_mstfsm_ctrl_cnt[0]), .op(
        n6929) );
  nor2_1 U8184 ( .ip1(n6929), .ip2(n6928), .op(n6930) );
  nand2_1 U8185 ( .ip1(n6931), .ip2(n6930), .op(n6933) );
  inv_1 U8186 ( .ip(i_ssi_U_mstfsm_c_done_ir), .op(n6932) );
  nand2_1 U8187 ( .ip1(n6933), .ip2(n6932), .op(n6934) );
  and2_1 U8188 ( .ip1(n6934), .ip2(n9972), .op(n11831) );
  inv_1 U8189 ( .ip(i_ssi_U_fifo_U_rx_fifo_empty_n), .op(n6935) );
  nor2_1 U8190 ( .ip1(n6936), .ip2(n6935), .op(n6938) );
  nand2_1 U8191 ( .ip1(n6938), .ip2(n6937), .op(n10131) );
  nand2_1 U8192 ( .ip1(n10749), .ip2(i_ssi_U_fifo_U_rx_fifo_rd_addr_at_max), 
        .op(n6939) );
  nand2_1 U8193 ( .ip1(n6939), .ip2(n10759), .op(n10133) );
  nor2_1 U8194 ( .ip1(n5614), .ip2(n10133), .op(i_ssi_U_fifo_U_rx_fifo_N46) );
  inv_1 U8195 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[15]), .op(
        n7158) );
  nand2_1 U8196 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[13]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[14]), .op(n7157) );
  nand2_1 U8197 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[10]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[11]), .op(n7156) );
  nand2_1 U8198 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[7]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[8]), .op(n7155) );
  nand2_1 U8199 ( .ip1(n8754), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[15]), .op(n6946) );
  nor2_1 U8200 ( .ip1(n8754), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[15]), .op(n6947) );
  nand2_1 U8201 ( .ip1(n8773), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[14]), .op(n6944) );
  or2_1 U8202 ( .ip1(n6947), .ip2(n6944), .op(n6945) );
  nand2_1 U8203 ( .ip1(n6946), .ip2(n6945), .op(n6954) );
  nor2_1 U8204 ( .ip1(n8773), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[14]), .op(n6948) );
  nor2_1 U8205 ( .ip1(n6948), .ip2(n6947), .op(n6957) );
  nand2_1 U8206 ( .ip1(n8778), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[13]), .op(n6951) );
  nor2_1 U8207 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[13]), .ip2(
        n8778), .op(n6956) );
  nand2_1 U8208 ( .ip1(n8620), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[12]), .op(n6949) );
  or2_1 U8209 ( .ip1(n6956), .ip2(n6949), .op(n6950) );
  nand2_1 U8210 ( .ip1(n6951), .ip2(n6950), .op(n6952) );
  and2_1 U8211 ( .ip1(n6957), .ip2(n6952), .op(n6953) );
  nor2_1 U8212 ( .ip1(n6954), .ip2(n6953), .op(n6972) );
  nor2_1 U8213 ( .ip1(n8620), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[12]), .op(n6955) );
  nor2_1 U8214 ( .ip1(n6956), .ip2(n6955), .op(n6958) );
  nand2_1 U8215 ( .ip1(n6958), .ip2(n6957), .op(n6977) );
  nand2_1 U8216 ( .ip1(n5273), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[11]), .op(n6961) );
  nor2_1 U8217 ( .ip1(n5273), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[11]), .op(n6962) );
  nand2_1 U8218 ( .ip1(n8761), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[10]), .op(n6959) );
  or2_1 U8219 ( .ip1(n6962), .ip2(n6959), .op(n6960) );
  nand2_1 U8220 ( .ip1(n6961), .ip2(n6960), .op(n6969) );
  nand2_1 U8221 ( .ip1(n5265), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[9]), .op(n6966) );
  nor2_1 U8222 ( .ip1(n5265), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[9]), .op(n6973) );
  nand2_1 U8223 ( .ip1(n5264), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[8]), .op(n6964) );
  or2_1 U8224 ( .ip1(n6973), .ip2(n6964), .op(n6965) );
  nand2_1 U8225 ( .ip1(n6966), .ip2(n6965), .op(n6967) );
  and2_1 U8226 ( .ip1(n6975), .ip2(n6967), .op(n6968) );
  nor2_1 U8227 ( .ip1(n6969), .ip2(n6968), .op(n6970) );
  or2_1 U8228 ( .ip1(n6977), .ip2(n6970), .op(n6971) );
  nand2_1 U8229 ( .ip1(n6972), .ip2(n6971), .op(n7017) );
  nor2_1 U8230 ( .ip1(n5264), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[8]), .op(n6974) );
  nor2_1 U8231 ( .ip1(n6974), .ip2(n6973), .op(n6976) );
  nand2_1 U8232 ( .ip1(n6976), .ip2(n6975), .op(n6978) );
  nor2_1 U8233 ( .ip1(n6978), .ip2(n6977), .op(n7015) );
  nand2_1 U8234 ( .ip1(n5597), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[7]), .op(n6981) );
  nor2_1 U8235 ( .ip1(n5597), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[7]), .op(n6982) );
  nand2_1 U8236 ( .ip1(n5598), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[6]), .op(n6979) );
  or2_1 U8237 ( .ip1(n6982), .ip2(n6979), .op(n6980) );
  nand2_1 U8238 ( .ip1(n6981), .ip2(n6980), .op(n6989) );
  nor2_1 U8239 ( .ip1(n5598), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[6]), .op(n6983) );
  nor2_1 U8240 ( .ip1(n6983), .ip2(n6982), .op(n7008) );
  nand2_1 U8241 ( .ip1(n8800), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[5]), .op(n6986) );
  nor2_1 U8242 ( .ip1(n8800), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[5]), .op(n7006) );
  nand2_1 U8243 ( .ip1(n8822), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[4]), .op(n6984) );
  or2_1 U8244 ( .ip1(n7006), .ip2(n6984), .op(n6985) );
  nand2_1 U8245 ( .ip1(n6986), .ip2(n6985), .op(n6987) );
  and2_1 U8246 ( .ip1(n7008), .ip2(n6987), .op(n6988) );
  nor2_1 U8247 ( .ip1(n6989), .ip2(n6988), .op(n7013) );
  nand2_1 U8248 ( .ip1(n5274), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[3]), .op(n6993) );
  nor2_1 U8249 ( .ip1(n5274), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[3]), .op(n6999) );
  nand2_1 U8250 ( .ip1(n8807), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[2]), .op(n6991) );
  or2_1 U8251 ( .ip1(n6999), .ip2(n6991), .op(n6992) );
  nand2_1 U8252 ( .ip1(n6993), .ip2(n6992), .op(n7004) );
  nand2_1 U8253 ( .ip1(n8811), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[1]), .op(n6998) );
  nor2_1 U8254 ( .ip1(n6994), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[0]), .op(n6996) );
  nor2_1 U8255 ( .ip1(n8811), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[1]), .op(n6995) );
  or2_1 U8256 ( .ip1(n6996), .ip2(n6995), .op(n6997) );
  nand2_1 U8257 ( .ip1(n6998), .ip2(n6997), .op(n7002) );
  nor2_1 U8258 ( .ip1(n8807), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[2]), .op(n7000) );
  nor2_1 U8259 ( .ip1(n7000), .ip2(n6999), .op(n7001) );
  and2_1 U8260 ( .ip1(n7002), .ip2(n7001), .op(n7003) );
  nor2_1 U8261 ( .ip1(n7004), .ip2(n7003), .op(n7011) );
  nor2_1 U8262 ( .ip1(n8822), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[4]), .op(n7007) );
  nor2_1 U8263 ( .ip1(n7007), .ip2(n7006), .op(n7009) );
  nand2_1 U8264 ( .ip1(n7009), .ip2(n7008), .op(n7010) );
  or2_1 U8265 ( .ip1(n7011), .ip2(n7010), .op(n7012) );
  nand2_1 U8266 ( .ip1(n7013), .ip2(n7012), .op(n7014) );
  and2_1 U8267 ( .ip1(n7015), .ip2(n7014), .op(n7016) );
  nor2_1 U8268 ( .ip1(n7017), .ip2(n7016), .op(n7020) );
  inv_1 U8269 ( .ip(n7018), .op(n7019) );
  nand2_1 U8270 ( .ip1(n7020), .ip2(n7019), .op(n7150) );
  nor2_1 U8271 ( .ip1(n8550), .ip2(n7062), .op(n7022) );
  nand2_1 U8272 ( .ip1(n7063), .ip2(n7022), .op(n7045) );
  nor2_1 U8273 ( .ip1(n7048), .ip2(n7044), .op(n7032) );
  inv_1 U8274 ( .ip(n7036), .op(n7023) );
  nand2_1 U8275 ( .ip1(n7032), .ip2(n7023), .op(n7024) );
  nor2_1 U8276 ( .ip1(n7045), .ip2(n7024), .op(n7029) );
  nor2_1 U8277 ( .ip1(n7096), .ip2(n7093), .op(n7027) );
  nor2_4 U8278 ( .ip1(n7090), .ip2(n7028), .op(n7073) );
  nand2_1 U8279 ( .ip1(n7029), .ip2(n7073), .op(n7030) );
  xnor2_1 U8280 ( .ip1(n7031), .ip2(n7030), .op(n8530) );
  nand2_1 U8281 ( .ip1(n5277), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[15]), .op(n7039) );
  nor2_1 U8282 ( .ip1(n5277), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[15]), .op(n7040) );
  inv_1 U8283 ( .ip(n7032), .op(n7033) );
  nor2_1 U8284 ( .ip1(n7045), .ip2(n7033), .op(n7034) );
  nand2_1 U8285 ( .ip1(n7034), .ip2(n7073), .op(n7035) );
  xnor2_1 U8286 ( .ip1(n7036), .ip2(n7035), .op(n8392) );
  nand2_1 U8287 ( .ip1(n5276), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[14]), .op(n7037) );
  or2_1 U8288 ( .ip1(n7040), .ip2(n7037), .op(n7038) );
  nand2_1 U8289 ( .ip1(n7039), .ip2(n7038), .op(n7054) );
  nor2_1 U8290 ( .ip1(n5276), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[14]), .op(n7041) );
  nor2_1 U8291 ( .ip1(n7041), .ip2(n7040), .op(n7057) );
  nor2_1 U8292 ( .ip1(n7045), .ip2(n7048), .op(n7042) );
  nand2_1 U8293 ( .ip1(n7042), .ip2(n7073), .op(n7043) );
  nand2_1 U8294 ( .ip1(n5268), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[13]), .op(n7051) );
  nor2_1 U8295 ( .ip1(n5268), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[13]), .op(n7055) );
  inv_1 U8296 ( .ip(n7045), .op(n7046) );
  nand2_1 U8297 ( .ip1(n7073), .ip2(n7046), .op(n7047) );
  xnor2_1 U8298 ( .ip1(n7048), .ip2(n7047), .op(n8537) );
  nand2_1 U8299 ( .ip1(n5275), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[12]), .op(n7049) );
  or2_1 U8300 ( .ip1(n7055), .ip2(n7049), .op(n7050) );
  nand2_1 U8301 ( .ip1(n7051), .ip2(n7050), .op(n7052) );
  and2_1 U8302 ( .ip1(n7057), .ip2(n7052), .op(n7053) );
  nor2_1 U8303 ( .ip1(n7054), .ip2(n7053), .op(n7082) );
  nor2_1 U8304 ( .ip1(n5275), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[12]), .op(n7056) );
  nor2_1 U8305 ( .ip1(n7056), .ip2(n7055), .op(n7058) );
  nand2_1 U8306 ( .ip1(n7058), .ip2(n7057), .op(n7087) );
  inv_1 U8307 ( .ip(n7063), .op(n7059) );
  nor2_1 U8308 ( .ip1(n7059), .ip2(n8550), .op(n7060) );
  nand2_1 U8309 ( .ip1(n7073), .ip2(n7060), .op(n7061) );
  nand2_1 U8310 ( .ip1(n5269), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[11]), .op(n7066) );
  nor2_1 U8311 ( .ip1(n5269), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[11]), .op(n7067) );
  nand2_1 U8312 ( .ip1(n7073), .ip2(n7063), .op(n8549) );
  nand2_1 U8313 ( .ip1(n8408), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[10]), .op(n7064) );
  or2_1 U8314 ( .ip1(n7067), .ip2(n7064), .op(n7065) );
  nand2_1 U8315 ( .ip1(n7066), .ip2(n7065), .op(n7079) );
  nor2_1 U8316 ( .ip1(n8408), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[10]), .op(n7068) );
  nor2_1 U8317 ( .ip1(n7068), .ip2(n7067), .op(n7085) );
  inv_1 U8318 ( .ip(n7072), .op(n7069) );
  nand2_1 U8319 ( .ip1(n8858), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[9]), .op(n7076) );
  nor2_1 U8320 ( .ip1(n8858), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[9]), .op(n7083) );
  nand2_1 U8321 ( .ip1(n5259), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[8]), .op(n7074) );
  or2_1 U8322 ( .ip1(n7083), .ip2(n7074), .op(n7075) );
  nand2_1 U8323 ( .ip1(n7076), .ip2(n7075), .op(n7077) );
  and2_1 U8324 ( .ip1(n7085), .ip2(n7077), .op(n7078) );
  nor2_1 U8325 ( .ip1(n7079), .ip2(n7078), .op(n7080) );
  or2_1 U8326 ( .ip1(n7087), .ip2(n7080), .op(n7081) );
  nand2_1 U8327 ( .ip1(n7082), .ip2(n7081), .op(n7145) );
  nor2_1 U8328 ( .ip1(n5259), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[8]), .op(n7084) );
  nor2_1 U8329 ( .ip1(n7084), .ip2(n7083), .op(n7086) );
  nand2_1 U8330 ( .ip1(n7086), .ip2(n7085), .op(n7088) );
  nor2_1 U8331 ( .ip1(n7088), .ip2(n7087), .op(n7143) );
  inv_1 U8332 ( .ip(n7094), .op(n7089) );
  nor2_1 U8333 ( .ip1(n7089), .ip2(n7096), .op(n7091) );
  inv_1 U8334 ( .ip(n7090), .op(n7106) );
  nand2_1 U8335 ( .ip1(n7091), .ip2(n7106), .op(n7092) );
  nand2_1 U8336 ( .ip1(n5266), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[7]), .op(n7099) );
  nor2_1 U8337 ( .ip1(n5266), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[7]), .op(n7100) );
  nand2_1 U8338 ( .ip1(n7106), .ip2(n7094), .op(n7095) );
  xnor2_1 U8339 ( .ip1(n7096), .ip2(n7095), .op(n8429) );
  nand2_1 U8340 ( .ip1(n5278), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[6]), .op(n7097) );
  or2_1 U8341 ( .ip1(n7100), .ip2(n7097), .op(n7098) );
  nand2_1 U8342 ( .ip1(n7099), .ip2(n7098), .op(n7112) );
  nor2_1 U8343 ( .ip1(n5278), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[6]), .op(n7101) );
  nor2_1 U8344 ( .ip1(n7101), .ip2(n7100), .op(n7136) );
  inv_1 U8345 ( .ip(n7105), .op(n7102) );
  nand2_1 U8346 ( .ip1(n7106), .ip2(n7102), .op(n7103) );
  xnor2_2 U8347 ( .ip1(n7104), .ip2(n7103), .op(n8879) );
  nand2_1 U8348 ( .ip1(n8879), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[5]), .op(n7109) );
  nor2_1 U8349 ( .ip1(n8879), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[5]), .op(n7134) );
  xor2_1 U8350 ( .ip1(n7106), .ip2(n7105), .op(n8435) );
  nand2_1 U8351 ( .ip1(n8457), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[4]), .op(n7107) );
  or2_1 U8352 ( .ip1(n7134), .ip2(n7107), .op(n7108) );
  nand2_1 U8353 ( .ip1(n7109), .ip2(n7108), .op(n7110) );
  and2_1 U8354 ( .ip1(n7136), .ip2(n7110), .op(n7111) );
  nor2_1 U8355 ( .ip1(n7112), .ip2(n7111), .op(n7141) );
  inv_1 U8356 ( .ip(n7113), .op(n7117) );
  nand2_1 U8357 ( .ip1(n8442), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[3]), .op(n7120) );
  nor2_1 U8358 ( .ip1(n8442), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[3]), .op(n7128) );
  xnor2_1 U8359 ( .ip1(n7117), .ip2(n7116), .op(n8443) );
  nand2_1 U8360 ( .ip1(n5280), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[2]), .op(n7118) );
  or2_1 U8361 ( .ip1(n7128), .ip2(n7118), .op(n7119) );
  nand2_1 U8362 ( .ip1(n7120), .ip2(n7119), .op(n7133) );
  nand2_1 U8363 ( .ip1(n5245), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[1]), .op(n7127) );
  nor2_1 U8364 ( .ip1(n7121), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[0]), .op(n7125) );
  nor2_1 U8365 ( .ip1(n5245), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[1]), .op(n7124) );
  or2_1 U8366 ( .ip1(n7125), .ip2(n7124), .op(n7126) );
  nand2_1 U8367 ( .ip1(n7127), .ip2(n7126), .op(n7131) );
  nor2_1 U8368 ( .ip1(n5280), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[2]), .op(n7129) );
  nor2_1 U8369 ( .ip1(n7129), .ip2(n7128), .op(n7130) );
  and2_1 U8370 ( .ip1(n7131), .ip2(n7130), .op(n7132) );
  nor2_1 U8371 ( .ip1(n7133), .ip2(n7132), .op(n7139) );
  nor2_1 U8372 ( .ip1(n8457), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[4]), .op(n7135) );
  nor2_1 U8373 ( .ip1(n7135), .ip2(n7134), .op(n7137) );
  nand2_1 U8374 ( .ip1(n7137), .ip2(n7136), .op(n7138) );
  or2_1 U8375 ( .ip1(n7139), .ip2(n7138), .op(n7140) );
  nand2_1 U8376 ( .ip1(n7141), .ip2(n7140), .op(n7142) );
  and2_1 U8377 ( .ip1(n7143), .ip2(n7142), .op(n7144) );
  nor2_1 U8378 ( .ip1(n7145), .ip2(n7144), .op(n7148) );
  inv_1 U8379 ( .ip(n8911), .op(n11052) );
  nand2_1 U8380 ( .ip1(n11052), .ip2(n7146), .op(n7147) );
  nand2_1 U8381 ( .ip1(n7148), .ip2(n7147), .op(n7149) );
  nand2_1 U8382 ( .ip1(n7150), .ip2(n7149), .op(n8385) );
  inv_1 U8383 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[0]), .op(n8345) );
  nand2_1 U8384 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[1]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[2]), .op(n7151) );
  nor2_1 U8385 ( .ip1(n8345), .ip2(n7151), .op(n8350) );
  nand2_1 U8386 ( .ip1(n5594), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[6]), .op(n8364) );
  nor2_1 U8387 ( .ip1(n7155), .ip2(n8364), .op(n8368) );
  nand2_1 U8388 ( .ip1(n8368), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[9]), .op(n8372) );
  nor2_1 U8389 ( .ip1(n7156), .ip2(n8372), .op(n8376) );
  nand2_1 U8390 ( .ip1(n8376), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[12]), .op(n8380) );
  nor2_1 U8391 ( .ip1(n7157), .ip2(n8380), .op(n8382) );
  xnor2_1 U8392 ( .ip1(n7158), .ip2(n8382), .op(n7159) );
  nand2_1 U8393 ( .ip1(n9890), .ip2(n7165), .op(n7163) );
  nor2_1 U8394 ( .ip1(n11836), .ip2(n7161), .op(n7162) );
  nand2_1 U8395 ( .ip1(n7163), .ip2(n7162), .op(n7168) );
  or2_1 U8396 ( .ip1(n7165), .ip2(n7164), .op(n7166) );
  nor2_1 U8397 ( .ip1(n7166), .ip2(n9890), .op(n7167) );
  nor2_1 U8398 ( .ip1(n7168), .ip2(n7167), .op(n4190) );
  nand2_1 U8399 ( .ip1(n5249), .ip2(i_apb_paddr[29]), .op(n7171) );
  nand2_1 U8400 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[29]), 
        .op(n7170) );
  nand2_1 U8401 ( .ip1(n7239), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[29]), 
        .op(n7169) );
  nand3_1 U8402 ( .ip1(n7171), .ip2(n7170), .ip3(n7169), .op(n4703) );
  nand2_1 U8403 ( .ip1(n10098), .ip2(i_apb_U_DW_apb_ahbsif_pipeline_c), .op(
        n10096) );
  nor2_1 U8404 ( .ip1(n10096), .ip2(n10105), .op(n9681) );
  nor2_1 U8405 ( .ip1(n9681), .ip2(n10095), .op(n7172) );
  nor2_1 U8406 ( .ip1(n7406), .ip2(n7172), .op(n7176) );
  nand2_1 U8407 ( .ip1(n7406), .ip2(n7173), .op(n7174) );
  nand2_1 U8408 ( .ip1(n7174), .ip2(n10083), .op(n7175) );
  and2_1 U8409 ( .ip1(n7175), .ip2(n10085), .op(n7177) );
  nand2_1 U8410 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[29]), 
        .op(n7182) );
  inv_1 U8411 ( .ip(n7406), .op(n7178) );
  nand2_1 U8412 ( .ip1(n7178), .ip2(n10095), .op(n7179) );
  nand2_1 U8413 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[29]), 
        .op(n7181) );
  nand2_1 U8414 ( .ip1(n7182), .ip2(n7181), .op(n4729) );
  nand2_1 U8415 ( .ip1(n5249), .ip2(i_apb_paddr[31]), .op(n7185) );
  nand2_1 U8416 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[31]), 
        .op(n7184) );
  nand2_1 U8417 ( .ip1(n7239), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[31]), 
        .op(n7183) );
  nand3_1 U8418 ( .ip1(n7185), .ip2(n7184), .ip3(n7183), .op(n4701) );
  nand2_1 U8419 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[31]), 
        .op(n7187) );
  nand2_1 U8420 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[31]), 
        .op(n7186) );
  nand2_1 U8421 ( .ip1(n7187), .ip2(n7186), .op(n4727) );
  nand2_1 U8422 ( .ip1(n5249), .ip2(i_apb_paddr[24]), .op(n7190) );
  nand2_1 U8423 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[24]), 
        .op(n7189) );
  nand2_1 U8424 ( .ip1(n7239), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[24]), 
        .op(n7188) );
  nand3_1 U8425 ( .ip1(n7190), .ip2(n7189), .ip3(n7188), .op(n4708) );
  nand2_1 U8426 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[24]), 
        .op(n7192) );
  nand2_1 U8427 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[24]), 
        .op(n7191) );
  nand2_1 U8428 ( .ip1(n7192), .ip2(n7191), .op(n4734) );
  nand2_1 U8429 ( .ip1(n5249), .ip2(i_apb_paddr[27]), .op(n7195) );
  nand2_1 U8430 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[27]), 
        .op(n7194) );
  nand2_1 U8431 ( .ip1(n7239), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[27]), 
        .op(n7193) );
  nand3_1 U8432 ( .ip1(n7195), .ip2(n7194), .ip3(n7193), .op(n4705) );
  nand2_1 U8433 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[27]), 
        .op(n7197) );
  nand2_1 U8434 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[27]), 
        .op(n7196) );
  nand2_1 U8435 ( .ip1(n7197), .ip2(n7196), .op(n4731) );
  nand2_1 U8436 ( .ip1(n5249), .ip2(i_apb_paddr[28]), .op(n7200) );
  nand2_1 U8437 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[28]), 
        .op(n7199) );
  nand2_1 U8438 ( .ip1(n7239), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[28]), 
        .op(n7198) );
  nand3_1 U8439 ( .ip1(n7200), .ip2(n7199), .ip3(n7198), .op(n4704) );
  nand2_1 U8440 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[28]), 
        .op(n7203) );
  nand2_1 U8441 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[28]), 
        .op(n7202) );
  nand2_1 U8442 ( .ip1(n7203), .ip2(n7202), .op(n4730) );
  nand2_1 U8443 ( .ip1(n5249), .ip2(i_apb_paddr[30]), .op(n7206) );
  nand2_1 U8444 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[30]), 
        .op(n7205) );
  nand2_1 U8445 ( .ip1(n7266), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[30]), 
        .op(n7204) );
  nand3_1 U8446 ( .ip1(n7206), .ip2(n7205), .ip3(n7204), .op(n4702) );
  nand2_1 U8447 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[30]), 
        .op(n7208) );
  nand2_1 U8448 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[30]), 
        .op(n7207) );
  nand2_1 U8449 ( .ip1(n7208), .ip2(n7207), .op(n4728) );
  nand2_1 U8450 ( .ip1(n5249), .ip2(i_apb_paddr[13]), .op(n7211) );
  nand2_1 U8451 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[13]), 
        .op(n7210) );
  nand2_1 U8452 ( .ip1(n7266), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[13]), 
        .op(n7209) );
  nand3_1 U8453 ( .ip1(n7211), .ip2(n7210), .ip3(n7209), .op(n4719) );
  nand2_1 U8454 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[13]), 
        .op(n7213) );
  nand2_1 U8455 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[13]), 
        .op(n7212) );
  nand2_1 U8456 ( .ip1(n7213), .ip2(n7212), .op(n4745) );
  nand2_1 U8457 ( .ip1(n5249), .ip2(i_apb_paddr[14]), .op(n7216) );
  nand2_1 U8458 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[14]), 
        .op(n7215) );
  nand2_1 U8459 ( .ip1(n7239), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[14]), 
        .op(n7214) );
  nand3_1 U8460 ( .ip1(n7216), .ip2(n7215), .ip3(n7214), .op(n4718) );
  nand2_1 U8461 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[14]), 
        .op(n7218) );
  nand2_1 U8462 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[14]), 
        .op(n7217) );
  nand2_1 U8463 ( .ip1(n7218), .ip2(n7217), .op(n4744) );
  nand2_1 U8464 ( .ip1(n5249), .ip2(i_apb_paddr[15]), .op(n7221) );
  nand2_1 U8465 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[15]), 
        .op(n7220) );
  nand2_1 U8466 ( .ip1(n7239), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[15]), 
        .op(n7219) );
  nand3_1 U8467 ( .ip1(n7221), .ip2(n7220), .ip3(n7219), .op(n4717) );
  nand2_1 U8468 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[15]), 
        .op(n7223) );
  nand2_1 U8469 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[15]), 
        .op(n7222) );
  nand2_1 U8470 ( .ip1(n7223), .ip2(n7222), .op(n4743) );
  nand2_1 U8471 ( .ip1(n5249), .ip2(i_apb_paddr[17]), .op(n7226) );
  nand2_1 U8472 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[17]), 
        .op(n7225) );
  nand2_1 U8473 ( .ip1(n7239), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[17]), 
        .op(n7224) );
  nand3_1 U8474 ( .ip1(n7226), .ip2(n7225), .ip3(n7224), .op(n4715) );
  nand2_1 U8475 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[17]), 
        .op(n7228) );
  nand2_1 U8476 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[17]), 
        .op(n7227) );
  nand2_1 U8477 ( .ip1(n7228), .ip2(n7227), .op(n4741) );
  nand2_1 U8478 ( .ip1(n5249), .ip2(i_apb_paddr[18]), .op(n7231) );
  nand2_1 U8479 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[18]), 
        .op(n7230) );
  nand2_1 U8480 ( .ip1(n7266), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[18]), 
        .op(n7229) );
  nand3_1 U8481 ( .ip1(n7231), .ip2(n7230), .ip3(n7229), .op(n4714) );
  nand2_1 U8482 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[18]), 
        .op(n7233) );
  nand2_1 U8483 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[18]), 
        .op(n7232) );
  nand2_1 U8484 ( .ip1(n7233), .ip2(n7232), .op(n4740) );
  nand2_1 U8485 ( .ip1(n5249), .ip2(i_apb_paddr[20]), .op(n7236) );
  nand2_1 U8486 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[20]), 
        .op(n7235) );
  nand2_1 U8487 ( .ip1(n7239), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[20]), 
        .op(n7234) );
  nand3_1 U8488 ( .ip1(n7236), .ip2(n7235), .ip3(n7234), .op(n4712) );
  nand2_1 U8489 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[20]), 
        .op(n7238) );
  nand2_1 U8490 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[20]), 
        .op(n7237) );
  nand2_1 U8491 ( .ip1(n7238), .ip2(n7237), .op(n4738) );
  nand2_1 U8492 ( .ip1(n5249), .ip2(i_apb_paddr[21]), .op(n7242) );
  nand2_1 U8493 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[21]), 
        .op(n7241) );
  nand2_1 U8494 ( .ip1(n7239), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[21]), 
        .op(n7240) );
  nand3_1 U8495 ( .ip1(n7242), .ip2(n7241), .ip3(n7240), .op(n4711) );
  nand2_1 U8496 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[21]), 
        .op(n7244) );
  nand2_1 U8497 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[21]), 
        .op(n7243) );
  nand2_1 U8498 ( .ip1(n7244), .ip2(n7243), .op(n4737) );
  nand2_1 U8499 ( .ip1(n5249), .ip2(i_apb_paddr[19]), .op(n7247) );
  nand2_1 U8500 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[19]), 
        .op(n7246) );
  nand2_1 U8501 ( .ip1(n7266), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[19]), 
        .op(n7245) );
  nand3_1 U8502 ( .ip1(n7247), .ip2(n7246), .ip3(n7245), .op(n4713) );
  nand2_1 U8503 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[19]), 
        .op(n7249) );
  nand2_1 U8504 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[19]), 
        .op(n7248) );
  nand2_1 U8505 ( .ip1(n7249), .ip2(n7248), .op(n4739) );
  nand2_1 U8506 ( .ip1(n5249), .ip2(i_apb_paddr[22]), .op(n7252) );
  nand2_1 U8507 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[22]), 
        .op(n7251) );
  nand2_1 U8508 ( .ip1(n7266), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[22]), 
        .op(n7250) );
  nand3_1 U8509 ( .ip1(n7252), .ip2(n7251), .ip3(n7250), .op(n4710) );
  nand2_1 U8510 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[22]), 
        .op(n7254) );
  nand2_1 U8511 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[22]), 
        .op(n7253) );
  nand2_1 U8512 ( .ip1(n7254), .ip2(n7253), .op(n4736) );
  nand2_1 U8513 ( .ip1(n5249), .ip2(i_apb_paddr[23]), .op(n7257) );
  nand2_1 U8514 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[23]), 
        .op(n7256) );
  nand2_1 U8515 ( .ip1(n7266), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[23]), 
        .op(n7255) );
  nand3_1 U8516 ( .ip1(n7257), .ip2(n7256), .ip3(n7255), .op(n4709) );
  nand2_1 U8517 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[23]), 
        .op(n7259) );
  nand2_1 U8518 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[23]), 
        .op(n7258) );
  nand2_1 U8519 ( .ip1(n7259), .ip2(n7258), .op(n4735) );
  nand2_1 U8520 ( .ip1(n5249), .ip2(i_apb_paddr[25]), .op(n7262) );
  nand2_1 U8521 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[25]), 
        .op(n7261) );
  nand2_1 U8522 ( .ip1(n7266), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[25]), 
        .op(n7260) );
  nand3_1 U8523 ( .ip1(n7262), .ip2(n7261), .ip3(n7260), .op(n4707) );
  nand2_1 U8524 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[25]), 
        .op(n7264) );
  nand2_1 U8525 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[25]), 
        .op(n7263) );
  nand2_1 U8526 ( .ip1(n7264), .ip2(n7263), .op(n4733) );
  nand2_1 U8527 ( .ip1(n5249), .ip2(i_apb_paddr[26]), .op(n7269) );
  nand2_1 U8528 ( .ip1(n7265), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[26]), 
        .op(n7268) );
  nand2_1 U8529 ( .ip1(n7266), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[26]), 
        .op(n7267) );
  nand3_1 U8530 ( .ip1(n7269), .ip2(n7268), .ip3(n7267), .op(n4706) );
  nand2_1 U8531 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[26]), 
        .op(n7271) );
  nand2_1 U8532 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[26]), 
        .op(n7270) );
  nand2_1 U8533 ( .ip1(n7271), .ip2(n7270), .op(n4732) );
  xor2_1 U8534 ( .ip1(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_flg_sync), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_flg_sync_q), .op(
        i_i2c_tx_abrt_flg_edg) );
  or2_1 U8535 ( .ip1(i_i2c_mst_activity_sync), .ip2(i_i2c_slv_activity_sync), 
        .op(i_i2c_activity) );
  inv_1 U8536 ( .ip(n11272), .op(n11280) );
  nor2_1 U8537 ( .ip1(i_i2c_slv_debug_cstate[0]), .ip2(
        i_i2c_slv_debug_cstate[2]), .op(n7302) );
  inv_1 U8538 ( .ip(i_i2c_slv_debug_cstate[1]), .op(n7959) );
  and2_1 U8539 ( .ip1(n7302), .ip2(n7959), .op(n11242) );
  nor2_1 U8540 ( .ip1(n11242), .ip2(n7272), .op(n11279) );
  or2_1 U8541 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[0]), .ip2(
        n11280), .op(n7298) );
  inv_1 U8542 ( .ip(i_i2c_ic_sda_setup[7]), .op(n7293) );
  inv_1 U8543 ( .ip(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[6]), .op(
        n11283) );
  inv_1 U8544 ( .ip(i_i2c_ic_sda_setup[5]), .op(n7288) );
  nor2_1 U8545 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[5]), .ip2(
        n7288), .op(n7290) );
  inv_1 U8546 ( .ip(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[4]), .op(n9329) );
  nor2_1 U8547 ( .ip1(i_i2c_ic_sda_setup[4]), .ip2(n9329), .op(n7287) );
  inv_1 U8548 ( .ip(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[2]), .op(
        n11259) );
  inv_1 U8549 ( .ip(i_i2c_ic_sda_setup[3]), .op(n7280) );
  nor2_1 U8550 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[3]), .ip2(
        n7280), .op(n7278) );
  inv_1 U8551 ( .ip(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[1]), .op(
        n11253) );
  nand2_1 U8552 ( .ip1(i_i2c_ic_sda_setup[1]), .ip2(n11253), .op(n7276) );
  inv_1 U8553 ( .ip(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[0]), .op(
        n11251) );
  nand2_1 U8554 ( .ip1(i_i2c_ic_sda_setup[0]), .ip2(n11251), .op(n7275) );
  nor2_1 U8555 ( .ip1(i_i2c_ic_sda_setup[2]), .ip2(n11259), .op(n7274) );
  nor2_1 U8556 ( .ip1(i_i2c_ic_sda_setup[1]), .ip2(n11253), .op(n7273) );
  not_ab_or_c_or_d U8557 ( .ip1(n7276), .ip2(n7275), .ip3(n7274), .ip4(n7273), 
        .op(n7277) );
  not_ab_or_c_or_d U8558 ( .ip1(i_i2c_ic_sda_setup[2]), .ip2(n11259), .ip3(
        n7278), .ip4(n7277), .op(n7279) );
  or2_1 U8559 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[3]), .ip2(
        n7279), .op(n7282) );
  or2_1 U8560 ( .ip1(n7280), .ip2(n7279), .op(n7281) );
  nand2_1 U8561 ( .ip1(n7282), .ip2(n7281), .op(n7283) );
  or2_1 U8562 ( .ip1(i_i2c_ic_sda_setup[4]), .ip2(n7283), .op(n7285) );
  or2_1 U8563 ( .ip1(n9329), .ip2(n7283), .op(n7284) );
  nand2_1 U8564 ( .ip1(n7285), .ip2(n7284), .op(n7286) );
  not_ab_or_c_or_d U8565 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[5]), .ip2(n7288), .ip3(n7287), .ip4(n7286), .op(n7289) );
  not_ab_or_c_or_d U8566 ( .ip1(i_i2c_ic_sda_setup[6]), .ip2(n11283), .ip3(
        n7290), .ip4(n7289), .op(n7292) );
  nor2_1 U8567 ( .ip1(i_i2c_ic_sda_setup[6]), .ip2(n11283), .op(n7291) );
  ab_or_c_or_d U8568 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[7]), 
        .ip2(n7293), .ip3(n7292), .ip4(n7291), .op(n7296) );
  inv_1 U8569 ( .ip(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[7]), .op(n7294) );
  nand2_1 U8570 ( .ip1(i_i2c_ic_sda_setup[7]), .ip2(n7294), .op(n7295) );
  nand2_1 U8571 ( .ip1(n7296), .ip2(n7295), .op(n11254) );
  or2_1 U8572 ( .ip1(n11254), .ip2(n11280), .op(n7297) );
  nand2_1 U8573 ( .ip1(n7298), .ip2(n7297), .op(n7299) );
  nor2_1 U8574 ( .ip1(n11279), .ip2(n7299), .op(n11252) );
  or2_1 U8575 ( .ip1(n11280), .ip2(n11252), .op(n7301) );
  or2_1 U8576 ( .ip1(n11251), .ip2(n11252), .op(n7300) );
  nand2_1 U8577 ( .ip1(n7301), .ip2(n7300), .op(n5211) );
  or2_1 U8578 ( .ip1(i_i2c_slv_debug_cstate[3]), .ip2(
        i_i2c_slv_debug_cstate[1]), .op(n9592) );
  inv_1 U8579 ( .ip(n9592), .op(n9584) );
  nand2_1 U8580 ( .ip1(n9584), .ip2(n7302), .op(i_i2c_U_DW_apb_i2c_slvfsm_N284) );
  nand2_1 U8581 ( .ip1(n7302), .ip2(n11019), .op(n9585) );
  inv_1 U8582 ( .ip(i_i2c_U_DW_apb_i2c_slvfsm_N284), .op(n7303) );
  or2_1 U8583 ( .ip1(n9585), .ip2(n7303), .op(n7305) );
  inv_1 U8584 ( .ip(i_i2c_slv_rx_2addr), .op(n11078) );
  or2_1 U8585 ( .ip1(n11078), .ip2(n7303), .op(n7304) );
  nand2_1 U8586 ( .ip1(n7305), .ip2(n7304), .op(n5224) );
  nand2_1 U8587 ( .ip1(i_i2c_ic_clr_rx_over_en), .ip2(n11839), .op(n7306) );
  nand2_1 U8588 ( .ip1(i_i2c_ic_clr_intr_en), .ip2(n11839), .op(n7312) );
  nand3_1 U8589 ( .ip1(n7306), .ip2(n7312), .ip3(i_i2c_ic_raw_intr_stat[1]), 
        .op(n7307) );
  inv_1 U8590 ( .ip(i_i2c_ic_en), .op(n11449) );
  or2_1 U8591 ( .ip1(n7307), .ip2(n11449), .op(n7311) );
  inv_1 U8592 ( .ip(i_i2c_U_DW_apb_i2c_fifo_rx_pop_dly), .op(n7308) );
  nand3_1 U8593 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_rx_error_ir), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_rx_push_sync_dly), .ip3(n7308), .op(n7309) );
  or2_1 U8594 ( .ip1(n7309), .ip2(n11449), .op(n7310) );
  nand2_1 U8595 ( .ip1(n7311), .ip2(n7310), .op(n4645) );
  inv_1 U8596 ( .ip(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_empty_n), .op(n5240) );
  nand2_1 U8597 ( .ip1(i_i2c_ic_clr_rx_under_en), .ip2(n11839), .op(n7313) );
  nand3_1 U8598 ( .ip1(n7313), .ip2(n7312), .ip3(i_i2c_ic_raw_intr_stat[0]), 
        .op(n7314) );
  or2_1 U8599 ( .ip1(n7314), .ip2(n11449), .op(n7317) );
  nand3_1 U8600 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_rx_error_ir), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_rx_pop_dly), .ip3(n5240), .op(n7315) );
  or2_1 U8601 ( .ip1(n7315), .ip2(n11449), .op(n7316) );
  nand2_1 U8602 ( .ip1(n7317), .ip2(n7316), .op(n4646) );
  nor2_1 U8603 ( .ip1(n9989), .ip2(n10982), .op(n7318) );
  nand2_1 U8604 ( .ip1(n7319), .ip2(n7318), .op(n7320) );
  inv_1 U8605 ( .ip(n7320), .op(n5226) );
  inv_1 U8606 ( .ip(i_ssi_fsm_multi_mst), .op(n7322) );
  nand2_1 U8607 ( .ip1(n11851), .ip2(n9988), .op(n7321) );
  xnor2_1 U8608 ( .ip1(n7322), .ip2(n7321), .op(n7323) );
  inv_1 U8609 ( .ip(n7323), .op(n4241) );
  inv_1 U8610 ( .ip(i_ssi_U_sclkgen_ssi_cnt[7]), .op(n7326) );
  nand2_1 U8611 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[6]), .ip2(
        i_ssi_U_sclkgen_ssi_cnt[5]), .op(n7325) );
  nand2_1 U8612 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[3]), .ip2(
        i_ssi_U_sclkgen_ssi_cnt[0]), .op(n7324) );
  nand2_1 U8613 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[1]), .ip2(
        i_ssi_U_sclkgen_ssi_cnt[2]), .op(n9763) );
  nor2_1 U8614 ( .ip1(n7324), .ip2(n9763), .op(n9765) );
  nand2_1 U8615 ( .ip1(n9765), .ip2(i_ssi_U_sclkgen_ssi_cnt[4]), .op(n9768) );
  nor2_1 U8616 ( .ip1(n7325), .ip2(n9768), .op(n9770) );
  xnor2_1 U8617 ( .ip1(n7326), .ip2(n9770), .op(n7382) );
  xor2_1 U8618 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[9]), .ip2(i_ssi_baudr[9]), .op(
        n7327) );
  inv_1 U8619 ( .ip(i_ssi_baudr[8]), .op(n10029) );
  xnor2_1 U8620 ( .ip1(n7327), .ip2(n5394), .op(n7328) );
  inv_1 U8621 ( .ip(n7328), .op(n7348) );
  xor2_1 U8622 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[3]), .ip2(n7329), .op(n7335) );
  inv_1 U8623 ( .ip(n7335), .op(n7331) );
  xor2_1 U8624 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[4]), .ip2(i_ssi_baudr[4]), .op(
        n7351) );
  inv_1 U8625 ( .ip(n7351), .op(n7330) );
  nand2_1 U8626 ( .ip1(n7331), .ip2(n7330), .op(n7332) );
  nand2_1 U8627 ( .ip1(n7332), .ip2(n6433), .op(n7333) );
  mux2_1 U8628 ( .ip1(n6433), .ip2(n7333), .s(i_ssi_U_sclkgen_ssi_cnt[2]), 
        .op(n7334) );
  nand2_1 U8629 ( .ip1(n7334), .ip2(i_ssi_U_sclkgen_ssi_cnt[1]), .op(n7347) );
  nor2_1 U8630 ( .ip1(n6432), .ip2(n7351), .op(n7336) );
  mux2_1 U8631 ( .ip1(n6432), .ip2(n7336), .s(n7335), .op(n7337) );
  inv_1 U8632 ( .ip(n7337), .op(n7345) );
  xor2_1 U8633 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[8]), .ip2(i_ssi_baudr[8]), .op(
        n7338) );
  xor2_1 U8634 ( .ip1(n7338), .ip2(n7361), .op(n7339) );
  xnor2_1 U8635 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[5]), .ip2(i_ssi_baudr[5]), .op(
        n7341) );
  xnor2_1 U8636 ( .ip1(n7341), .ip2(n7340), .op(n7342) );
  inv_1 U8637 ( .ip(n7342), .op(n7343) );
  nand2_1 U8638 ( .ip1(n7339), .ip2(n7343), .op(n7344) );
  nor2_1 U8639 ( .ip1(n7345), .ip2(n7344), .op(n7346) );
  inv_1 U8640 ( .ip(i_ssi_U_sclkgen_ssi_cnt[1]), .op(n9754) );
  xor2_1 U8641 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[2]), .ip2(i_ssi_baudr[2]), .op(
        n7349) );
  ab_or_c_or_d U8642 ( .ip1(n7351), .ip2(n9763), .ip3(n9764), .ip4(n7350), 
        .op(n7352) );
  xnor2_1 U8643 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[14]), .ip2(i_ssi_baudr[14]), 
        .op(n7353) );
  xnor2_1 U8644 ( .ip1(n7353), .ip2(n7379), .op(n7356) );
  xor2_1 U8645 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[13]), .ip2(i_ssi_baudr[13]), 
        .op(n7355) );
  xor2_1 U8646 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[7]), .ip2(i_ssi_baudr[7]), .op(
        n7358) );
  nor2_1 U8647 ( .ip1(i_ssi_baudr[6]), .ip2(n7366), .op(n7357) );
  xnor2_1 U8648 ( .ip1(n7358), .ip2(n7357), .op(n7377) );
  xor2_1 U8649 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[11]), .ip2(i_ssi_baudr[11]), 
        .op(n7364) );
  nor2_1 U8650 ( .ip1(i_ssi_baudr[9]), .ip2(i_ssi_baudr[8]), .op(n7360) );
  inv_1 U8651 ( .ip(i_ssi_baudr[10]), .op(n7359) );
  nand2_1 U8652 ( .ip1(n7360), .ip2(n7359), .op(n7362) );
  or2_1 U8653 ( .ip1(n7362), .ip2(n7361), .op(n7363) );
  xnor2_1 U8654 ( .ip1(n7364), .ip2(n7363), .op(n7365) );
  inv_1 U8655 ( .ip(n7365), .op(n7369) );
  xor2_1 U8656 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[6]), .ip2(i_ssi_baudr[6]), .op(
        n7367) );
  xor2_1 U8657 ( .ip1(n7367), .ip2(n7366), .op(n7368) );
  and2_1 U8658 ( .ip1(n7369), .ip2(n7368), .op(n7376) );
  xor2_1 U8659 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[10]), .ip2(i_ssi_baudr[10]), 
        .op(n7372) );
  xnor2_1 U8660 ( .ip1(n7372), .ip2(n7371), .op(n7375) );
  xnor2_1 U8661 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[15]), .ip2(i_ssi_baudr[15]), 
        .op(n7381) );
  nor2_1 U8662 ( .ip1(i_ssi_baudr[14]), .ip2(n7379), .op(n7380) );
  xnor2_1 U8663 ( .ip1(n7381), .ip2(n7380), .op(n9794) );
  or2_1 U8664 ( .ip1(n7397), .ip2(n5291), .op(n7386) );
  inv_1 U8665 ( .ip(n5435), .op(n9755) );
  inv_1 U8666 ( .ip(n9755), .op(n9760) );
  nand2_1 U8667 ( .ip1(n7382), .ip2(n9760), .op(n7383) );
  inv_1 U8668 ( .ip(n7383), .op(i_ssi_U_sclkgen_N47) );
  inv_1 U8669 ( .ip(i_ssi_U_sclkgen_ssi_cnt[10]), .op(n7385) );
  nand2_1 U8670 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[9]), .ip2(
        i_ssi_U_sclkgen_ssi_cnt[8]), .op(n7384) );
  nand2_1 U8671 ( .ip1(n9770), .ip2(i_ssi_U_sclkgen_ssi_cnt[7]), .op(n9774) );
  nor2_1 U8672 ( .ip1(n7384), .ip2(n9774), .op(n9776) );
  xnor2_1 U8673 ( .ip1(n7385), .ip2(n9776), .op(n7387) );
  nand2_1 U8674 ( .ip1(n7387), .ip2(n5284), .op(n7388) );
  inv_1 U8675 ( .ip(n7388), .op(i_ssi_U_sclkgen_N50) );
  xnor2_1 U8676 ( .ip1(n6422), .ip2(n9765), .op(n7389) );
  nand2_1 U8677 ( .ip1(n7389), .ip2(n5284), .op(n7390) );
  inv_1 U8678 ( .ip(n7390), .op(i_ssi_U_sclkgen_N44) );
  nand2_1 U8679 ( .ip1(n5435), .ip2(n9764), .op(n7391) );
  nand2_1 U8680 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[12]), .ip2(
        i_ssi_U_sclkgen_ssi_cnt[11]), .op(n7392) );
  nand2_1 U8681 ( .ip1(n9776), .ip2(i_ssi_U_sclkgen_ssi_cnt[10]), .op(n9780)
         );
  nor2_1 U8682 ( .ip1(n7392), .ip2(n9780), .op(n9787) );
  and2_1 U8683 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[13]), .ip2(
        i_ssi_U_sclkgen_ssi_cnt[14]), .op(n7393) );
  and2_1 U8684 ( .ip1(n9787), .ip2(n7393), .op(n9789) );
  xor2_1 U8685 ( .ip1(n7394), .ip2(n9789), .op(n7395) );
  or2_1 U8686 ( .ip1(n7395), .ip2(n5291), .op(n7396) );
  nor2_1 U8687 ( .ip1(n5477), .ip2(n7396), .op(i_ssi_U_sclkgen_N55) );
  or2_1 U8688 ( .ip1(n7917), .ip2(n10926), .op(n11022) );
  or2_1 U8689 ( .ip1(n10919), .ip2(n10941), .op(n8968) );
  nor2_1 U8690 ( .ip1(n11022), .ip2(n8968), .op(n7400) );
  nand2_1 U8691 ( .ip1(n10943), .ip2(i_i2c_mst_debug_cstate[0]), .op(n10917)
         );
  inv_1 U8692 ( .ip(n10917), .op(n10938) );
  and2_1 U8693 ( .ip1(i_i2c_tx_fifo_data_buf[8]), .ip2(
        i_i2c_U_DW_apb_i2c_sync_ic_rstrt_en_sync_inv), .op(n7851) );
  inv_1 U8694 ( .ip(n7851), .op(n7399) );
  nand2_1 U8695 ( .ip1(n10938), .ip2(n7399), .op(n11064) );
  nand2_1 U8696 ( .ip1(n7400), .ip2(n11064), .op(n7402) );
  nand2_1 U8697 ( .ip1(n7402), .ip2(n7401), .op(n9488) );
  xor2_1 U8698 ( .ip1(n7829), .ip2(i_i2c_ack_det), .op(n7803) );
  nand2_1 U8699 ( .ip1(n7802), .ip2(n7803), .op(n7905) );
  inv_1 U8700 ( .ip(n7905), .op(n7403) );
  nor2_1 U8701 ( .ip1(n7403), .ip2(n9473), .op(n7404) );
  nor2_1 U8702 ( .ip1(n9488), .ip2(n7404), .op(n11834) );
  nor2_1 U8703 ( .ip1(n8065), .ip2(n6352), .op(n11835) );
  inv_1 U8704 ( .ip(i_i2c_ic_hs), .op(n11840) );
  inv_1 U8705 ( .ip(i_ssi_ssi_rst_n), .op(n11841) );
  inv_1 U8706 ( .ip(i_i2c_ic_rst_n), .op(n11843) );
  inv_1 U8707 ( .ip(i_i2c_ic_rst_n), .op(n11842) );
  inv_1 U8708 ( .ip(PRESETn_presetn), .op(n11845) );
  nand2_1 U8709 ( .ip1(n7405), .ip2(n10098), .op(n7415) );
  mux2_1 U8710 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_hwrite_c), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwrite), .s(n9690), .op(n4846) );
  nor2_1 U8711 ( .ip1(n10099), .ip2(n7406), .op(n7410) );
  inv_1 U8712 ( .ip(n7410), .op(n7407) );
  nand2_1 U8713 ( .ip1(n7407), .ip2(i_apb_U_DW_apb_ahbsif_state[1]), .op(n7409) );
  nand2_1 U8714 ( .ip1(n7409), .ip2(n7408), .op(n7423) );
  nor2_1 U8715 ( .ip1(n7413), .ip2(n7410), .op(n7411) );
  not_ab_or_c_or_d U8716 ( .ip1(i_apb_U_DW_apb_ahbsif_state[0]), .ip2(n7413), 
        .ip3(n10101), .ip4(n7411), .op(n7412) );
  not_ab_or_c_or_d U8717 ( .ip1(n9684), .ip2(n7413), .ip3(
        i_apb_U_DW_apb_ahbsif_state[2]), .ip4(n7412), .op(n7414) );
  or2_1 U8718 ( .ip1(i_apb_pclk_en), .ip2(n7414), .op(n7421) );
  nor2_1 U8719 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_hwrite_c), .ip2(n7428), .op(
        n7417) );
  nor2_1 U8720 ( .ip1(n7416), .ip2(n7415), .op(n10103) );
  nor4_1 U8721 ( .ip1(n10105), .ip2(n7418), .ip3(n7417), .ip4(n10103), .op(
        n7419) );
  nand2_1 U8722 ( .ip1(i_apb_pclk_en), .ip2(n7419), .op(n7420) );
  nand2_1 U8723 ( .ip1(n7421), .ip2(n7420), .op(n7422) );
  mux2_1 U8724 ( .ip1(n7423), .ip2(i_apb_U_DW_apb_ahbsif_pipeline_c), .s(n7422), .op(n4847) );
  nand2_1 U8725 ( .ip1(n10091), .ip2(n9684), .op(n7424) );
  nand2_1 U8726 ( .ip1(n7424), .ip2(i_apb_U_DW_apb_ahbsif_use_saved_c), .op(
        n7427) );
  inv_1 U8727 ( .ip(n10095), .op(n10093) );
  inv_1 U8728 ( .ip(n10083), .op(n10092) );
  nand2_1 U8729 ( .ip1(n10092), .ip2(n10085), .op(n7425) );
  nand2_1 U8730 ( .ip1(n10093), .ip2(n7425), .op(n7426) );
  nand2_1 U8731 ( .ip1(n7427), .ip2(n7426), .op(n4819) );
  or2_1 U8732 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[16]), .ip2(n9690), 
        .op(n4835) );
  nand2_1 U8733 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[16]), 
        .op(n7431) );
  nand2_1 U8734 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[16]), 
        .op(n7430) );
  nor3_1 U8735 ( .ip1(n7428), .ip2(n10094), .ip3(n10095), .op(n9692) );
  nand2_1 U8736 ( .ip1(n9692), .ip2(i_apb_U_DW_apb_ahbsif_piped_haddr_c[16]), 
        .op(n7429) );
  nand3_1 U8737 ( .ip1(n7431), .ip2(n7430), .ip3(n7429), .op(n4742) );
  xor2_1 U8738 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_tx_pop_flg_sync), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_pop_flg_sync_q), .op(i_i2c_tx_pop_sync) );
  inv_1 U8739 ( .ip(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_empty_n), .op(n11862) );
  inv_1 U8740 ( .ip(i_i2c_tx_fifo_rst_n), .op(n11026) );
  inv_1 U8741 ( .ip(i_i2c_tx_pop_sync), .op(n11216) );
  nor2_1 U8742 ( .ip1(n11216), .ip2(n11862), .op(n11215) );
  inv_1 U8743 ( .ip(i_i2c_tx_push), .op(n9626) );
  not_ab_or_c_or_d U8744 ( .ip1(i_i2c_tx_full), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_empty_n), .ip3(n11215), .ip4(n9626), 
        .op(n7434) );
  inv_1 U8745 ( .ip(n11215), .op(n11227) );
  nor2_1 U8746 ( .ip1(i_i2c_tx_push), .ip2(n11227), .op(n7964) );
  nor2_1 U8747 ( .ip1(n7434), .ip2(n7964), .op(n7432) );
  xor2_1 U8748 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[0]), .ip2(n7432), 
        .op(n7433) );
  nor2_1 U8749 ( .ip1(n11026), .ip2(n7433), .op(n11867) );
  inv_1 U8750 ( .ip(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[0]), .op(n7436) );
  nor2_1 U8751 ( .ip1(n7434), .ip2(n7436), .op(n7966) );
  nor2_1 U8752 ( .ip1(n7964), .ip2(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[1]), 
        .op(n7435) );
  not_ab_or_c_or_d U8753 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[1]), 
        .ip2(n7436), .ip3(n7966), .ip4(n7435), .op(n7437) );
  xnor2_1 U8754 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[2]), .ip2(n7437), 
        .op(n11031) );
  nor2_1 U8755 ( .ip1(n11026), .ip2(n11031), .op(n11866) );
  inv_1 U8756 ( .ip(i_i2c_ic_clk_in_a), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_U_SYNC_N2) );
  inv_1 U8757 ( .ip(i_i2c_ic_data_in_a), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_U_SYNC_N2) );
  inv_1 U8758 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[4]), .op(
        n7507) );
  inv_1 U8759 ( .ip(i_i2c_ic_fs_spklen[5]), .op(n7549) );
  nor2_1 U8760 ( .ip1(n7549), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[5]), .op(n7450) );
  and2_1 U8761 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[3]), 
        .ip2(n7438), .op(n7448) );
  inv_1 U8762 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[3]), .op(
        n7506) );
  nor2_1 U8763 ( .ip1(n7440), .ip2(n7501), .op(n7446) );
  inv_1 U8764 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[0]), .op(
        n7495) );
  nand2_1 U8765 ( .ip1(n7495), .ip2(i_i2c_ic_fs_spklen[0]), .op(n7444) );
  inv_1 U8766 ( .ip(n7439), .op(n7442) );
  and2_1 U8767 ( .ip1(n7501), .ip2(n7440), .op(n7441) );
  not_ab_or_c_or_d U8768 ( .ip1(n7444), .ip2(n7443), .ip3(n7442), .ip4(n7441), 
        .op(n7445) );
  not_ab_or_c_or_d U8769 ( .ip1(i_i2c_ic_fs_spklen[3]), .ip2(n7506), .ip3(
        n7446), .ip4(n7445), .op(n7447) );
  not_ab_or_c_or_d U8770 ( .ip1(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[4]), .ip2(n9095), .ip3(
        n7448), .ip4(n7447), .op(n7449) );
  ab_or_c_or_d U8771 ( .ip1(i_i2c_ic_fs_spklen[4]), .ip2(n7507), .ip3(n7450), 
        .ip4(n7449), .op(n7453) );
  and2_1 U8772 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[5]), 
        .ip2(n7549), .op(n7451) );
  not_ab_or_c_or_d U8773 ( .ip1(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[6]), .ip2(n9093), .ip3(
        n7451), .ip4(n7454), .op(n7452) );
  nand2_1 U8774 ( .ip1(n7453), .ip2(n7452), .op(n7459) );
  inv_1 U8775 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[6]), .op(
        n7513) );
  nand2_1 U8776 ( .ip1(n7513), .ip2(i_i2c_ic_fs_spklen[6]), .op(n7455) );
  nor2_1 U8777 ( .ip1(n7455), .ip2(n7454), .op(n7456) );
  nor2_1 U8778 ( .ip1(n7457), .ip2(n7456), .op(n7458) );
  nand2_1 U8779 ( .ip1(n7459), .ip2(n7458), .op(n7461) );
  nand2_1 U8780 ( .ip1(n7461), .ip2(n7460), .op(n7492) );
  nand2_1 U8781 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[3]), 
        .ip2(n7462), .op(n7464) );
  nand2_1 U8782 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[4]), 
        .ip2(n9094), .op(n7463) );
  nand2_1 U8783 ( .ip1(n7464), .ip2(n7463), .op(n7474) );
  nor2_1 U8784 ( .ip1(n7470), .ip2(n7501), .op(n7472) );
  nor2_1 U8785 ( .ip1(n7465), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[0]), .op(n7467) );
  nor2_1 U8786 ( .ip1(n7467), .ip2(n7466), .op(n7468) );
  not_ab_or_c_or_d U8787 ( .ip1(n7501), .ip2(n7470), .ip3(n7469), .ip4(n7468), 
        .op(n7471) );
  not_ab_or_c_or_d U8788 ( .ip1(i_i2c_ic_hs_spklen[3]), .ip2(n7506), .ip3(
        n7472), .ip4(n7471), .op(n7473) );
  or2_1 U8789 ( .ip1(n7474), .ip2(n7473), .op(n7478) );
  nor2_1 U8790 ( .ip1(n7479), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[5]), .op(n7476) );
  nor2_1 U8791 ( .ip1(n9094), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[4]), .op(n7475) );
  nor2_1 U8792 ( .ip1(n7476), .ip2(n7475), .op(n7477) );
  nand2_1 U8793 ( .ip1(n7478), .ip2(n7477), .op(n7483) );
  nand2_1 U8794 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[6]), 
        .ip2(n9092), .op(n7481) );
  nand2_1 U8795 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[5]), 
        .ip2(n7479), .op(n7480) );
  nand2_1 U8796 ( .ip1(n7483), .ip2(n7482), .op(n7487) );
  nor2_1 U8797 ( .ip1(n9092), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[6]), .op(n7485) );
  nor2_1 U8798 ( .ip1(n7485), .ip2(n7484), .op(n7486) );
  nand2_1 U8799 ( .ip1(n7487), .ip2(n7486), .op(n7490) );
  inv_1 U8800 ( .ip(n7488), .op(n7489) );
  nand2_1 U8801 ( .ip1(n7490), .ip2(n7489), .op(n7491) );
  nand2_1 U8802 ( .ip1(n7492), .ip2(n7491), .op(n9529) );
  xnor2_1 U8803 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_U_scl_sync_data_d_int_0_), 
        .ip2(i_i2c_U_DW_apb_i2c_rx_filter_scl_clk_int), .op(n7493) );
  nand2_1 U8804 ( .ip1(n9529), .ip2(n7493), .op(n7517) );
  nor2_1 U8805 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[0]), 
        .ip2(n7517), .op(n11865) );
  nor2_1 U8806 ( .ip1(n7495), .ip2(n7517), .op(n7494) );
  mux2_1 U8807 ( .ip1(n7494), .ip2(n11865), .s(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[1]), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_N83) );
  nand2_1 U8808 ( .ip1(n11865), .ip2(n7501), .op(n7500) );
  inv_1 U8809 ( .ip(n7517), .op(n7498) );
  nor2_1 U8810 ( .ip1(n7501), .ip2(n7495), .op(n7496) );
  mux2_1 U8811 ( .ip1(n7501), .ip2(n7496), .s(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[1]), .op(n7497) );
  nand2_1 U8812 ( .ip1(n7498), .ip2(n7497), .op(n7499) );
  nand2_1 U8813 ( .ip1(n7500), .ip2(n7499), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_N84) );
  nand2_1 U8814 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[1]), 
        .ip2(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[0]), .op(n7503) );
  inv_1 U8815 ( .ip(n7503), .op(n7502) );
  nand2_1 U8816 ( .ip1(n7502), .ip2(n7501), .op(n7505) );
  nor3_1 U8817 ( .ip1(n7504), .ip2(n7506), .ip3(n7503), .op(n7509) );
  not_ab_or_c_or_d U8818 ( .ip1(n7506), .ip2(n7505), .ip3(n7509), .ip4(n7517), 
        .op(i_i2c_U_DW_apb_i2c_rx_filter_N85) );
  xor2_1 U8819 ( .ip1(n7507), .ip2(n7509), .op(n7508) );
  nor2_1 U8820 ( .ip1(n7508), .ip2(n7517), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_N86) );
  nand2_1 U8821 ( .ip1(n7509), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[4]), .op(n7511) );
  xor2_1 U8822 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[5]), 
        .ip2(n7511), .op(n7510) );
  nor2_1 U8823 ( .ip1(n7510), .ip2(n7517), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_N87) );
  inv_1 U8824 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[5]), .op(
        n7512) );
  nor2_1 U8825 ( .ip1(n7512), .ip2(n7511), .op(n7515) );
  xor2_1 U8826 ( .ip1(n7513), .ip2(n7515), .op(n7514) );
  nor2_1 U8827 ( .ip1(n7514), .ip2(n7517), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_N88) );
  and2_1 U8828 ( .ip1(n7515), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[6]), .op(n7516) );
  nor2_1 U8829 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_scl_spklen_cnt[7]), 
        .ip2(n7516), .op(n7518) );
  nor2_1 U8830 ( .ip1(n7518), .ip2(n7517), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_N89) );
  inv_1 U8831 ( .ip(n7519), .op(n7522) );
  nand3_1 U8832 ( .ip1(n7522), .ip2(n7521), .ip3(n7520), .op(n7527) );
  nand2_1 U8833 ( .ip1(n7524), .ip2(n7523), .op(n7525) );
  nand3_1 U8834 ( .ip1(n7527), .ip2(n7526), .ip3(n7525), .op(n7529) );
  nand2_1 U8835 ( .ip1(n7529), .ip2(n7528), .op(n7535) );
  nand2_1 U8836 ( .ip1(n7531), .ip2(n7530), .op(n7532) );
  nand2_1 U8837 ( .ip1(n7533), .ip2(n7532), .op(n7534) );
  nand2_1 U8838 ( .ip1(n7535), .ip2(n7534), .op(n7536) );
  and2_1 U8839 ( .ip1(n7536), .ip2(i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r), .op(
        n7564) );
  inv_1 U8840 ( .ip(n7537), .op(n7539) );
  nand4_1 U8841 ( .ip1(n7540), .ip2(n7539), .ip3(n7538), .ip4(n7542), .op(
        n7548) );
  inv_1 U8842 ( .ip(n7541), .op(n7544) );
  nor2_1 U8843 ( .ip1(n7544), .ip2(n7542), .op(n7546) );
  nor2_1 U8844 ( .ip1(n7544), .ip2(n7543), .op(n7545) );
  or2_1 U8845 ( .ip1(n7546), .ip2(n7545), .op(n7547) );
  nand2_1 U8846 ( .ip1(n7548), .ip2(n7547), .op(n7552) );
  nand2_1 U8847 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[5]), 
        .ip2(n7549), .op(n7550) );
  nand3_1 U8848 ( .ip1(n7552), .ip2(n7551), .ip3(n7550), .op(n7554) );
  inv_1 U8849 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[5]), .op(
        n7580) );
  nand2_1 U8850 ( .ip1(n7580), .ip2(i_i2c_ic_fs_spklen[5]), .op(n7553) );
  nand2_1 U8851 ( .ip1(n7554), .ip2(n7553), .op(n7558) );
  inv_1 U8852 ( .ip(n7555), .op(n7557) );
  not_ab_or_c_or_d U8853 ( .ip1(n7559), .ip2(n7558), .ip3(n7557), .ip4(n7556), 
        .op(n7560) );
  nor3_1 U8854 ( .ip1(n7562), .ip2(n7561), .ip3(n7560), .op(n7563) );
  nor2_1 U8855 ( .ip1(n7564), .ip2(n7563), .op(n7588) );
  inv_1 U8856 ( .ip(n7588), .op(n7566) );
  inv_1 U8857 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_U_sda_sync_data_d_int_0_), 
        .op(n7590) );
  nor2_1 U8858 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[0]), 
        .ip2(n7585), .op(i_i2c_U_DW_apb_i2c_rx_filter_N123) );
  and2_1 U8859 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[1]), 
        .ip2(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[0]), .op(n7569) );
  not_ab_or_c_or_d U8860 ( .ip1(n7568), .ip2(n7567), .ip3(n7569), .ip4(n7585), 
        .op(i_i2c_U_DW_apb_i2c_rx_filter_N124) );
  inv_1 U8861 ( .ip(n7569), .op(n7570) );
  and2_1 U8862 ( .ip1(n7569), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[2]), .op(n7572) );
  not_ab_or_c_or_d U8863 ( .ip1(n7571), .ip2(n7570), .ip3(n7572), .ip4(n7585), 
        .op(i_i2c_U_DW_apb_i2c_rx_filter_N125) );
  inv_1 U8864 ( .ip(n7572), .op(n7573) );
  and2_1 U8865 ( .ip1(n7572), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[3]), .op(n7575) );
  not_ab_or_c_or_d U8866 ( .ip1(n7574), .ip2(n7573), .ip3(n7575), .ip4(n7585), 
        .op(i_i2c_U_DW_apb_i2c_rx_filter_N126) );
  inv_1 U8867 ( .ip(n7575), .op(n7576) );
  and2_1 U8868 ( .ip1(n7575), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[4]), .op(n7578) );
  not_ab_or_c_or_d U8869 ( .ip1(n7577), .ip2(n7576), .ip3(n7578), .ip4(n7585), 
        .op(i_i2c_U_DW_apb_i2c_rx_filter_N127) );
  inv_1 U8870 ( .ip(n7578), .op(n7579) );
  and2_1 U8871 ( .ip1(n7578), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[5]), .op(n7581) );
  not_ab_or_c_or_d U8872 ( .ip1(n7580), .ip2(n7579), .ip3(n7581), .ip4(n7585), 
        .op(i_i2c_U_DW_apb_i2c_rx_filter_N128) );
  inv_1 U8873 ( .ip(n7581), .op(n7582) );
  and2_1 U8874 ( .ip1(n7581), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[6]), .op(n7584) );
  not_ab_or_c_or_d U8875 ( .ip1(n7583), .ip2(n7582), .ip3(n7584), .ip4(n7585), 
        .op(i_i2c_U_DW_apb_i2c_rx_filter_N129) );
  nor2_1 U8876 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_spklen_cnt[7]), 
        .ip2(n7584), .op(n7586) );
  nor2_1 U8877 ( .ip1(n7586), .ip2(n7585), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_N130) );
  nand2_1 U8878 ( .ip1(n7588), .ip2(n7587), .op(n7589) );
  mux2_1 U8879 ( .ip1(n7590), .ip2(i_i2c_U_DW_apb_i2c_rx_filter_sda_data_int), 
        .s(n7589), .op(n5129) );
  inv_1 U8880 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[5]), .op(
        n7648) );
  nand2_1 U8881 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[2]), 
        .ip2(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[1]), .op(n7643)
         );
  or2_1 U8882 ( .ip1(n7591), .ip2(n7601), .op(n7639) );
  nand2_1 U8883 ( .ip1(n7639), .ip2(n7640), .op(n7593) );
  inv_1 U8884 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[7]), .op(
        n7592) );
  nand2_1 U8885 ( .ip1(n7593), .ip2(n7592), .op(n7597) );
  inv_1 U8886 ( .ip(n7601), .op(n7594) );
  nand2_1 U8887 ( .ip1(i_i2c_ic_sda_rx_hold_sync[6]), .ip2(n7599), .op(n7600)
         );
  nand2_1 U8888 ( .ip1(n7594), .ip2(n7600), .op(n7595) );
  inv_1 U8889 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[6]), .op(
        n7664) );
  nand2_1 U8890 ( .ip1(n7595), .ip2(n7664), .op(n7596) );
  nand2_1 U8891 ( .ip1(n7597), .ip2(n7596), .op(n7678) );
  nand2_1 U8892 ( .ip1(i_i2c_ic_sda_rx_hold_sync[5]), .ip2(n7613), .op(n7598)
         );
  nand2_1 U8893 ( .ip1(n7599), .ip2(n7598), .op(n7605) );
  nor2_1 U8894 ( .ip1(n7648), .ip2(n7605), .op(n7604) );
  nand2_1 U8895 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[6]), 
        .ip2(n7600), .op(n7602) );
  nor2_1 U8896 ( .ip1(n7602), .ip2(n7601), .op(n7603) );
  nor2_1 U8897 ( .ip1(n7604), .ip2(n7603), .op(n7675) );
  nand2_1 U8898 ( .ip1(n7605), .ip2(n7648), .op(n7608) );
  nand2_1 U8899 ( .ip1(n7611), .ip2(i_i2c_ic_sda_rx_hold_sync[4]), .op(n7614)
         );
  nand2_1 U8900 ( .ip1(n7614), .ip2(n7613), .op(n7606) );
  inv_1 U8901 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[4]), .op(
        n7660) );
  nand2_1 U8902 ( .ip1(n7606), .ip2(n7660), .op(n7607) );
  and2_1 U8903 ( .ip1(n7608), .ip2(n7607), .op(n7634) );
  inv_1 U8904 ( .ip(i_i2c_ic_sda_rx_hold_sync[2]), .op(n7625) );
  nor2_1 U8905 ( .ip1(i_i2c_ic_sda_rx_hold_sync[1]), .ip2(
        i_i2c_ic_sda_rx_hold_sync[0]), .op(n7624) );
  nand2_1 U8906 ( .ip1(n7625), .ip2(n7624), .op(n7609) );
  nand2_1 U8907 ( .ip1(i_i2c_ic_sda_rx_hold_sync[3]), .ip2(n7609), .op(n7610)
         );
  nand2_1 U8908 ( .ip1(n7611), .ip2(n7610), .op(n7629) );
  inv_1 U8909 ( .ip(n7629), .op(n7612) );
  nand2_1 U8910 ( .ip1(n7612), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[3]), .op(n7616) );
  nand3_1 U8911 ( .ip1(n7614), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[4]), .ip3(n7613), .op(
        n7615) );
  nand2_1 U8912 ( .ip1(n7616), .ip2(n7615), .op(n7669) );
  nand2_1 U8913 ( .ip1(n7634), .ip2(n7669), .op(n7617) );
  nand2_1 U8914 ( .ip1(n7675), .ip2(n7617), .op(n7637) );
  nand2_1 U8915 ( .ip1(i_i2c_ic_sda_rx_hold_sync[0]), .ip2(
        i_i2c_ic_sda_rx_hold_sync[1]), .op(n7619) );
  inv_1 U8916 ( .ip(n7624), .op(n7618) );
  and2_1 U8917 ( .ip1(n7619), .ip2(n7618), .op(n7626) );
  inv_1 U8918 ( .ip(n7626), .op(n7621) );
  inv_1 U8919 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[1]), .op(
        n7620) );
  nand2_1 U8920 ( .ip1(n7621), .ip2(n7620), .op(n7623) );
  or2_1 U8921 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[0]), 
        .ip2(i_i2c_ic_sda_rx_hold_sync[0]), .op(n7622) );
  and2_1 U8922 ( .ip1(n7623), .ip2(n7622), .op(n7670) );
  xor2_1 U8923 ( .ip1(n7625), .ip2(n7624), .op(n7630) );
  nand2_1 U8924 ( .ip1(n7626), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[1]), .op(n7627) );
  nand2_1 U8925 ( .ip1(n7628), .ip2(n7627), .op(n7671) );
  nor2_1 U8926 ( .ip1(n7670), .ip2(n7671), .op(n7635) );
  inv_1 U8927 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[3]), .op(
        n7657) );
  nand2_1 U8928 ( .ip1(n7629), .ip2(n7657), .op(n7632) );
  or2_1 U8929 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[2]), 
        .ip2(n7630), .op(n7631) );
  and2_1 U8930 ( .ip1(n7632), .ip2(n7631), .op(n7633) );
  nand2_1 U8931 ( .ip1(n7634), .ip2(n7633), .op(n7679) );
  nor2_1 U8932 ( .ip1(n7635), .ip2(n7679), .op(n7636) );
  nor2_1 U8933 ( .ip1(n7637), .ip2(n7636), .op(n7638) );
  nor2_1 U8934 ( .ip1(n7678), .ip2(n7638), .op(n7642) );
  nand3_1 U8935 ( .ip1(n7639), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[7]), .ip3(n7640), .op(
        n7676) );
  nand2_1 U8936 ( .ip1(n7676), .ip2(n7640), .op(n7641) );
  nor2_1 U8937 ( .ip1(n7642), .ip2(n7641), .op(n7652) );
  nand2_1 U8938 ( .ip1(n7652), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[0]), .op(n7654) );
  nor2_1 U8939 ( .ip1(n7643), .ip2(n7654), .op(n7656) );
  and2_1 U8940 ( .ip1(n7656), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[3]), .op(n7659) );
  nand2_1 U8941 ( .ip1(n7659), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[4]), .op(n7647) );
  nand2_1 U8942 ( .ip1(n7645), .ip2(n6352), .op(n7667) );
  nand3_1 U8943 ( .ip1(n7659), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[5]), .ip3(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[4]), .op(n7663) );
  inv_1 U8944 ( .ip(n7663), .op(n7646) );
  not_ab_or_c_or_d U8945 ( .ip1(n7648), .ip2(n7647), .ip3(n7667), .ip4(n7646), 
        .op(n5091) );
  inv_1 U8946 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[2]), .op(
        n7651) );
  inv_1 U8947 ( .ip(n7654), .op(n7649) );
  nand2_1 U8948 ( .ip1(n7649), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[1]), .op(n7650) );
  not_ab_or_c_or_d U8949 ( .ip1(n7651), .ip2(n7650), .ip3(n7656), .ip4(n7667), 
        .op(n5094) );
  xnor2_1 U8950 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[0]), 
        .ip2(n7652), .op(n7653) );
  nor2_1 U8951 ( .ip1(n7667), .ip2(n7653), .op(n5096) );
  xor2_1 U8952 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[1]), 
        .ip2(n7654), .op(n7655) );
  nor2_1 U8953 ( .ip1(n7667), .ip2(n7655), .op(n5095) );
  xor2_1 U8954 ( .ip1(n7657), .ip2(n7656), .op(n7658) );
  xor2_1 U8955 ( .ip1(n7660), .ip2(n7659), .op(n7661) );
  xor2_1 U8956 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[6]), 
        .ip2(n7663), .op(n7662) );
  nor2_1 U8957 ( .ip1(n7667), .ip2(n7662), .op(n5090) );
  nor2_1 U8958 ( .ip1(n7664), .ip2(n7663), .op(n7665) );
  nor2_1 U8959 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[7]), 
        .ip2(n7665), .op(n7666) );
  nor2_1 U8960 ( .ip1(n7667), .ip2(n7666), .op(n5089) );
  inv_1 U8961 ( .ip(n7668), .op(n7682) );
  inv_1 U8962 ( .ip(n7669), .op(n7674) );
  inv_1 U8963 ( .ip(n7670), .op(n7672) );
  not_ab_or_c_or_d U8964 ( .ip1(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_sda_rx_hold_cnt[0]), .ip2(
        i_i2c_ic_sda_rx_hold_sync[0]), .ip3(n7672), .ip4(n7671), .op(n7673) );
  nand4_1 U8965 ( .ip1(n7676), .ip2(n7675), .ip3(n7674), .ip4(n7673), .op(
        n7677) );
  nor3_1 U8966 ( .ip1(n7679), .ip2(n7678), .ip3(n7677), .op(n7680) );
  nor2_1 U8967 ( .ip1(n9533), .ip2(n7680), .op(n7681) );
  mux2_1 U8968 ( .ip1(n7682), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_sda_post_hold_done), .s(n7681), .op(n5097) );
  inv_1 U8969 ( .ip(i_i2c_ic_master), .op(
        i_i2c_U_DW_apb_i2c_sync_U_ic_master_1_sync_N2) );
  inv_1 U8970 ( .ip(i_i2c_ic_10bit_mst), .op(
        i_i2c_U_DW_apb_i2c_sync_U_ic_10bit_mst_1_sync_N2) );
  nor2_1 U8971 ( .ip1(n7684), .ip2(n7683), .op(n7686) );
  and2_1 U8972 ( .ip1(n7686), .ip2(n7685), .op(n7730) );
  inv_1 U8973 ( .ip(n7730), .op(n8745) );
  nand3_1 U8974 ( .ip1(n8745), .ip2(i_i2c_U_DW_apb_i2c_mstfsm_addr_2byte_sent), 
        .ip3(i_i2c_U_DW_apb_i2c_mstfsm_N487), .op(n7687) );
  nand2_1 U8975 ( .ip1(n7687), .ip2(n10917), .op(n5199) );
  nand2_1 U8976 ( .ip1(n7689), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[14]), .op(n7690) );
  xnor2_1 U8977 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[15]), .ip2(
        n7690), .op(n7691) );
  inv_1 U8978 ( .ip(n7691), .op(n7692) );
  nor2_1 U8979 ( .ip1(n7729), .ip2(n7692), .op(i_i2c_U_DW_apb_i2c_clk_gen_N77)
         );
  nand2_1 U8980 ( .ip1(n7688), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[12]), .op(n7693) );
  not_ab_or_c_or_d U8981 ( .ip1(n7694), .ip2(n7693), .ip3(n7689), .ip4(n7729), 
        .op(i_i2c_U_DW_apb_i2c_clk_gen_N75) );
  nand2_1 U8982 ( .ip1(n7695), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[9]), .op(n7697) );
  not_ab_or_c_or_d U8983 ( .ip1(n5979), .ip2(n7697), .ip3(n7696), .ip4(n7729), 
        .op(i_i2c_U_DW_apb_i2c_clk_gen_N72) );
  or2_1 U8984 ( .ip1(n7716), .ip2(n7698), .op(n7721) );
  nand2_1 U8985 ( .ip1(n7699), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[6]), .op(n7701) );
  nor2_1 U8986 ( .ip1(n7700), .ip2(n7716), .op(n7723) );
  not_ab_or_c_or_d U8987 ( .ip1(n7702), .ip2(n7701), .ip3(n7723), .ip4(n7729), 
        .op(i_i2c_U_DW_apb_i2c_clk_gen_N69) );
  inv_1 U8988 ( .ip(n7716), .op(n7703) );
  nand2_1 U8989 ( .ip1(n7703), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[3]), .op(n7705) );
  nand2_1 U8990 ( .ip1(n7703), .ip2(n6006), .op(n7718) );
  inv_1 U8991 ( .ip(n7718), .op(n7704) );
  not_ab_or_c_or_d U8992 ( .ip1(n5940), .ip2(n7705), .ip3(n7704), .ip4(n7729), 
        .op(i_i2c_U_DW_apb_i2c_clk_gen_N66) );
  inv_1 U8993 ( .ip(n7712), .op(n7706) );
  nand2_1 U8994 ( .ip1(n7706), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[0]), .op(n7707) );
  not_ab_or_c_or_d U8995 ( .ip1(n7708), .ip2(n7707), .ip3(n7714), .ip4(n7729), 
        .op(i_i2c_U_DW_apb_i2c_clk_gen_N63) );
  and2_1 U8996 ( .ip1(n6352), .ip2(n7709), .op(n7710) );
  and2_1 U8997 ( .ip1(n11833), .ip2(n7710), .op(n11864) );
  nor2_1 U8998 ( .ip1(i_i2c_p_det), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_count_en), 
        .op(n7711) );
  nor2_1 U8999 ( .ip1(i_i2c_s_det), .ip2(n7711), .op(n4118) );
  xor2_1 U9000 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[0]), .ip2(n7712), .op(n7713) );
  nor2_1 U9001 ( .ip1(n7729), .ip2(n7713), .op(i_i2c_U_DW_apb_i2c_clk_gen_N62)
         );
  xor2_1 U9002 ( .ip1(n5934), .ip2(n7714), .op(n7715) );
  nor2_1 U9003 ( .ip1(n7729), .ip2(n7715), .op(i_i2c_U_DW_apb_i2c_clk_gen_N64)
         );
  nor2_1 U9004 ( .ip1(n7729), .ip2(n7717), .op(i_i2c_U_DW_apb_i2c_clk_gen_N65)
         );
  nor2_1 U9005 ( .ip1(n7729), .ip2(n7720), .op(i_i2c_U_DW_apb_i2c_clk_gen_N67)
         );
  nor2_1 U9006 ( .ip1(n7729), .ip2(n7722), .op(i_i2c_U_DW_apb_i2c_clk_gen_N68)
         );
  xor2_1 U9007 ( .ip1(n5972), .ip2(n7723), .op(n7724) );
  nor2_1 U9008 ( .ip1(n7729), .ip2(n7724), .op(i_i2c_U_DW_apb_i2c_clk_gen_N70)
         );
  xor2_1 U9009 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_bus_idle_cntr[9]), .ip2(n7725), .op(n7726) );
  xor2_1 U9010 ( .ip1(n5987), .ip2(n7688), .op(n7727) );
  xor2_1 U9011 ( .ip1(n5996), .ip2(n7689), .op(n7728) );
  inv_1 U9012 ( .ip(i_i2c_U_DW_apb_i2c_mstfsm_N382), .op(n7775) );
  nand2_1 U9013 ( .ip1(n7775), .ip2(i_i2c_scl_s_hld_cmplt), .op(n7871) );
  nand2_1 U9014 ( .ip1(n7730), .ip2(n7871), .op(n7900) );
  nand2_1 U9015 ( .ip1(i_i2c_scl_lcnt_cmplt), .ip2(i_i2c_scl_p_setup_cmplt), 
        .op(n9333) );
  inv_1 U9016 ( .ip(n9333), .op(n7731) );
  nand2_1 U9017 ( .ip1(n7856), .ip2(n7731), .op(n7732) );
  nand2_1 U9018 ( .ip1(n7900), .ip2(n7732), .op(n5225) );
  inv_1 U9019 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[0]), .op(n7733) );
  xor2_1 U9020 ( .ip1(n7733), .ip2(n7771), .op(n7734) );
  xor2_1 U9021 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[1]), .ip2(n7736), 
        .op(n7735) );
  inv_1 U9022 ( .ip(n7736), .op(n7737) );
  nand2_1 U9023 ( .ip1(n7737), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[1]), .op(n7738) );
  not_ab_or_c_or_d U9024 ( .ip1(n6255), .ip2(n7738), .ip3(n7739), .ip4(n7774), 
        .op(n5125) );
  inv_1 U9025 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[3]), .op(n7740) );
  xor2_1 U9026 ( .ip1(n7740), .ip2(n7739), .op(n7741) );
  xor2_1 U9027 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[4]), .ip2(n7743), 
        .op(n7742) );
  nor2_1 U9028 ( .ip1(n7774), .ip2(n7742), .op(n5123) );
  inv_1 U9029 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[5]), .op(n7746) );
  inv_1 U9030 ( .ip(n7743), .op(n7744) );
  nand2_1 U9031 ( .ip1(n7744), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[4]), .op(n7745) );
  not_ab_or_c_or_d U9032 ( .ip1(n7746), .ip2(n7745), .ip3(n7747), .ip4(n7774), 
        .op(n5122) );
  xor2_1 U9033 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[7]), .ip2(n7750), 
        .op(n7749) );
  nor2_1 U9034 ( .ip1(n7774), .ip2(n7749), .op(n5120) );
  inv_1 U9035 ( .ip(n7750), .op(n7751) );
  nand2_1 U9036 ( .ip1(n7751), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[7]), .op(n7752) );
  not_ab_or_c_or_d U9037 ( .ip1(n6280), .ip2(n7752), .ip3(n7753), .ip4(n7774), 
        .op(n5119) );
  inv_1 U9038 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[9]), .op(n7754) );
  nor2_1 U9039 ( .ip1(n7774), .ip2(n7755), .op(n5118) );
  xor2_1 U9040 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[10]), .ip2(n7758), .op(n7756) );
  nor2_1 U9041 ( .ip1(n7774), .ip2(n7756), .op(n5117) );
  inv_1 U9042 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[11]), .op(n7762)
         );
  nand2_1 U9043 ( .ip1(n7759), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[10]), .op(n7761) );
  inv_1 U9044 ( .ip(n7757), .op(n7760) );
  inv_1 U9045 ( .ip(n7758), .op(n7759) );
  not_ab_or_c_or_d U9046 ( .ip1(n7762), .ip2(n7761), .ip3(n7763), .ip4(n7774), 
        .op(n5116) );
  nand2_1 U9047 ( .ip1(n7763), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[12]), .op(n7766) );
  xor2_1 U9048 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[13]), .ip2(n7766), .op(n7764) );
  nor2_1 U9049 ( .ip1(n7774), .ip2(n7764), .op(n5114) );
  inv_1 U9050 ( .ip(n7766), .op(n7765) );
  nand2_1 U9051 ( .ip1(n7765), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[13]), .op(n7768) );
  nand2_1 U9052 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[13]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_min_hld_cntr[14]), .op(n7767) );
  nor2_1 U9053 ( .ip1(n7767), .ip2(n7766), .op(n7769) );
  not_ab_or_c_or_d U9054 ( .ip1(n6248), .ip2(n7768), .ip3(n7769), .ip4(n7774), 
        .op(n5113) );
  nor2_1 U9055 ( .ip1(n7774), .ip2(n7770), .op(n5128) );
  inv_1 U9056 ( .ip(n7771), .op(n7772) );
  nor2_1 U9057 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_N382), .ip2(n7772), .op(n7773)
         );
  nor2_1 U9058 ( .ip1(n7774), .ip2(n7773), .op(n5112) );
  inv_1 U9059 ( .ip(n5225), .op(n8991) );
  nand2_1 U9060 ( .ip1(n8991), .ip2(i_i2c_start_en), .op(n7921) );
  inv_1 U9061 ( .ip(i_i2c_scl_s_hld_cmplt), .op(n8337) );
  nor2_1 U9062 ( .ip1(n7775), .ip2(n8337), .op(n7916) );
  nand2_1 U9063 ( .ip1(n7776), .ip2(i_i2c_mst_rx_ack_vld), .op(n7777) );
  nand2_1 U9064 ( .ip1(n9473), .ip2(n7777), .op(n7809) );
  inv_1 U9065 ( .ip(n7809), .op(n7782) );
  inv_1 U9066 ( .ip(n7829), .op(n7786) );
  inv_1 U9067 ( .ip(n7808), .op(n7780) );
  nor2_1 U9068 ( .ip1(n7786), .ip2(n7780), .op(n7781) );
  nand2_1 U9069 ( .ip1(n7782), .ip2(n7781), .op(n11035) );
  inv_1 U9070 ( .ip(n11035), .op(n8119) );
  nand2_1 U9071 ( .ip1(n8119), .ip2(n11055), .op(n7784) );
  nand2_1 U9072 ( .ip1(n7856), .ip2(n9333), .op(n7783) );
  nand2_1 U9073 ( .ip1(n7784), .ip2(n7783), .op(n7790) );
  xor2_1 U9074 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_old_is_read), .ip2(
        i_i2c_tx_fifo_data_buf[8]), .op(n7823) );
  nand2_1 U9075 ( .ip1(n7823), .ip2(i_i2c_U_DW_apb_i2c_mstfsm_addr_2byte_sent), 
        .op(n7887) );
  inv_1 U9076 ( .ip(i_i2c_U_DW_apb_i2c_mstfsm_addr_1byte_sent), .op(n7785) );
  nand2_1 U9077 ( .ip1(n7887), .ip2(n7785), .op(n7847) );
  inv_1 U9078 ( .ip(n7847), .op(n7788) );
  nand2_1 U9079 ( .ip1(n7808), .ip2(n7786), .op(n7787) );
  nor2_1 U9080 ( .ip1(n7787), .ip2(n7809), .op(n7816) );
  inv_1 U9081 ( .ip(i_i2c_U_DW_apb_i2c_sync_ic_10bit_mst_sync_inv), .op(n7825)
         );
  and2_1 U9082 ( .ip1(n7816), .ip2(n7825), .op(n7888) );
  inv_1 U9083 ( .ip(n7888), .op(n7846) );
  nor2_1 U9084 ( .ip1(n7788), .ip2(n7846), .op(n7789) );
  nor2_1 U9085 ( .ip1(n7790), .ip2(n7789), .op(n7884) );
  inv_1 U9086 ( .ip(n8332), .op(n10902) );
  nand3_1 U9087 ( .ip1(n7791), .ip2(i_i2c_ack_det), .ip3(
        i_i2c_U_DW_apb_i2c_sync_tx_empty_int_inv), .op(n7801) );
  inv_1 U9088 ( .ip(i_i2c_U_DW_apb_i2c_sync_ic_rstrt_en_sync_inv), .op(n7852)
         );
  nand3_1 U9089 ( .ip1(n11055), .ip2(
        i_i2c_U_DW_apb_i2c_sync_ic_10bit_mst_sync_inv), .ip3(n7852), .op(n7799) );
  inv_1 U9090 ( .ip(n7874), .op(n7795) );
  nor2_1 U9091 ( .ip1(n7868), .ip2(n7869), .op(n7792) );
  not_ab_or_c_or_d U9092 ( .ip1(n7868), .ip2(n7873), .ip3(n7793), .ip4(n7792), 
        .op(n7794) );
  nor2_1 U9093 ( .ip1(n7795), .ip2(n7794), .op(n7798) );
  or2_1 U9094 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(n11021), .op(n7922) );
  nand2_1 U9095 ( .ip1(n7895), .ip2(i_i2c_scl_s_hld_cmplt), .op(n7796) );
  nand2_1 U9096 ( .ip1(n7922), .ip2(n7796), .op(n7797) );
  not_ab_or_c_or_d U9097 ( .ip1(n7865), .ip2(n7799), .ip3(n7798), .ip4(n7797), 
        .op(n7800) );
  nand2_1 U9098 ( .ip1(n7801), .ip2(n7800), .op(n7807) );
  inv_1 U9099 ( .ip(n7802), .op(n7828) );
  inv_1 U9100 ( .ip(n7803), .op(n7804) );
  nor2_1 U9101 ( .ip1(n7804), .ip2(n9473), .op(n7805) );
  nor2_1 U9102 ( .ip1(n7828), .ip2(n7805), .op(n7806) );
  not_ab_or_c_or_d U9103 ( .ip1(n10902), .ip2(n9473), .ip3(n7807), .ip4(n7806), 
        .op(n7814) );
  nand2_1 U9104 ( .ip1(n7809), .ip2(n7808), .op(n7813) );
  inv_1 U9105 ( .ip(n11073), .op(n7864) );
  nand3_1 U9106 ( .ip1(n7810), .ip2(n11064), .ip3(n11071), .op(n7811) );
  nand2_1 U9107 ( .ip1(n7864), .ip2(n7811), .op(n7812) );
  nand3_1 U9108 ( .ip1(n7814), .ip2(n7813), .ip3(n7812), .op(n7821) );
  inv_1 U9109 ( .ip(n7823), .op(n7815) );
  nor2_1 U9110 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_rstrt_en_sync_inv), .ip2(
        n7815), .op(n7819) );
  nand2_1 U9111 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_10bit_mst_sync_inv), .ip2(
        i_i2c_U_DW_apb_i2c_mstfsm_addr_1byte_sent), .op(n7817) );
  inv_1 U9112 ( .ip(n7816), .op(n7824) );
  nor2_1 U9113 ( .ip1(n7817), .ip2(n7824), .op(n7912) );
  inv_1 U9114 ( .ip(n7912), .op(n7818) );
  nor2_1 U9115 ( .ip1(n7819), .ip2(n7818), .op(n7820) );
  nor2_1 U9116 ( .ip1(n7821), .ip2(n7820), .op(n7822) );
  nand2_1 U9117 ( .ip1(n7884), .ip2(n7822), .op(n8058) );
  nand2_1 U9118 ( .ip1(n7823), .ip2(
        i_i2c_U_DW_apb_i2c_sync_ic_rstrt_en_sync_inv), .op(n7826) );
  not_ab_or_c_or_d U9119 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_addr_1byte_sent), 
        .ip2(n7826), .ip3(n7825), .ip4(n7824), .op(n7843) );
  nand2_1 U9120 ( .ip1(n7864), .ip2(n10926), .op(n8108) );
  nand3_1 U9121 ( .ip1(n7895), .ip2(i_i2c_U_DW_apb_i2c_mstfsm_N252), .ip3(
        i_i2c_scl_s_hld_cmplt), .op(n7827) );
  nand2_1 U9122 ( .ip1(n7827), .ip2(n8745), .op(n7834) );
  nor2_1 U9123 ( .ip1(n7829), .ip2(n7828), .op(n10930) );
  and3_1 U9124 ( .ip1(n7832), .ip2(n7845), .ip3(i_i2c_mst_debug_cstate[3]), 
        .op(n7833) );
  nand2_1 U9125 ( .ip1(n11073), .ip2(n7917), .op(n7835) );
  nand3_1 U9126 ( .ip1(n8108), .ip2(n7836), .ip3(n7835), .op(n7842) );
  nor2_1 U9127 ( .ip1(i_i2c_ic_abort_sync), .ip2(n11861), .op(n7837) );
  and2_1 U9128 ( .ip1(n7864), .ip2(n7837), .op(n7886) );
  inv_1 U9129 ( .ip(n7886), .op(n7838) );
  inv_1 U9130 ( .ip(n9473), .op(n8993) );
  and3_1 U9131 ( .ip1(n7838), .ip2(n8993), .ip3(n10941), .op(n7841) );
  nor2_1 U9132 ( .ip1(n10942), .ip2(n8119), .op(n7839) );
  nor2_1 U9133 ( .ip1(n11055), .ip2(n7839), .op(n7840) );
  nor2_1 U9134 ( .ip1(n7845), .ip2(n7844), .op(n7849) );
  nor2_1 U9135 ( .ip1(n7847), .ip2(n7846), .op(n7848) );
  nor2_1 U9136 ( .ip1(n7849), .ip2(n7848), .op(n7885) );
  nor2_1 U9137 ( .ip1(n7852), .ip2(n7887), .op(n7850) );
  nand2_1 U9138 ( .ip1(n7888), .ip2(n7850), .op(n7861) );
  and2_1 U9139 ( .ip1(n10938), .ip2(n7851), .op(n11061) );
  nand3_1 U9140 ( .ip1(n11055), .ip2(i_i2c_mst_rxbyte_rdy), .ip3(n7852), .op(
        n7854) );
  nor2_1 U9141 ( .ip1(n7854), .ip2(n7853), .op(n7855) );
  nor2_1 U9142 ( .ip1(n7855), .ip2(n11021), .op(n7857) );
  ab_or_c_or_d U9143 ( .ip1(n7858), .ip2(n9333), .ip3(n7857), .ip4(n7856), 
        .op(n7859) );
  not_ab_or_c_or_d U9144 ( .ip1(n10938), .ip2(n11073), .ip3(n11061), .ip4(
        n7859), .op(n7860) );
  nand2_1 U9145 ( .ip1(n7861), .ip2(n7860), .op(n7911) );
  inv_1 U9146 ( .ip(n7911), .op(n7862) );
  nand3_1 U9147 ( .ip1(n7863), .ip2(n7885), .ip3(n7862), .op(n8989) );
  nand2_1 U9148 ( .ip1(n7864), .ip2(n10942), .op(n7867) );
  nand2_1 U9149 ( .ip1(n7865), .ip2(i_i2c_mst_rxbyte_rdy), .op(n7866) );
  nand2_1 U9150 ( .ip1(n7867), .ip2(n7866), .op(n7882) );
  inv_1 U9151 ( .ip(n10930), .op(n11074) );
  inv_1 U9152 ( .ip(n10926), .op(n10905) );
  nand2_1 U9153 ( .ip1(n11074), .ip2(n10905), .op(n7881) );
  or2_1 U9154 ( .ip1(i_i2c_ack_det), .ip2(n9473), .op(n11070) );
  inv_1 U9155 ( .ip(n11070), .op(n8111) );
  nand2_1 U9156 ( .ip1(n7868), .ip2(i_i2c_mst_debug_cstate[3]), .op(n7870) );
  nor3_1 U9157 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_10bit_mst_sync_inv), .ip2(
        n7871), .ip3(n8745), .op(n7872) );
  not_ab_or_c_or_d U9158 ( .ip1(n7874), .ip2(n7873), .ip3(n7896), .ip4(n7872), 
        .op(n7878) );
  nand2_1 U9159 ( .ip1(n9473), .ip2(n8968), .op(n7877) );
  nand3_1 U9160 ( .ip1(n10919), .ip2(i_i2c_ack_det), .ip3(n7875), .op(n7876)
         );
  nand3_1 U9161 ( .ip1(n7878), .ip2(n7877), .ip3(n7876), .op(n7880) );
  nor2_1 U9162 ( .ip1(n11064), .ip2(n8111), .op(n7879) );
  not_ab_or_c_or_d U9163 ( .ip1(n11055), .ip2(n7882), .ip3(n5248), .ip4(n7912), 
        .op(n7883) );
  nand3_1 U9164 ( .ip1(n7885), .ip2(n7884), .ip3(n7883), .op(n8053) );
  nor2_1 U9165 ( .ip1(n11068), .ip2(n7886), .op(n7913) );
  nand3_1 U9166 ( .ip1(n7888), .ip2(i_i2c_U_DW_apb_i2c_mstfsm_addr_1byte_sent), 
        .ip3(n7887), .op(n7909) );
  nor2_1 U9167 ( .ip1(i_i2c_tx_fifo_data_buf[8]), .ip2(n10917), .op(n7904) );
  nor2_1 U9168 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv), .ip2(n7889), 
        .op(n7903) );
  nand2_1 U9169 ( .ip1(i_i2c_ic_tar[10]), .ip2(i_i2c_U_DW_apb_i2c_mstfsm_N252), 
        .op(n11094) );
  nand2_1 U9170 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv), .ip2(n11094), 
        .op(n7890) );
  nand2_1 U9171 ( .ip1(n7890), .ip2(
        i_i2c_U_DW_apb_i2c_sync_ic_rstrt_en_sync_inv), .op(n7891) );
  inv_1 U9172 ( .ip(i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv), .op(n11091)
         );
  nand2_1 U9173 ( .ip1(n7891), .ip2(n11091), .op(n8113) );
  inv_1 U9174 ( .ip(i_i2c_U_DW_apb_i2c_mstfsm_N487), .op(n8121) );
  inv_1 U9175 ( .ip(i_i2c_U_DW_apb_i2c_mstfsm_tx_empty_hld), .op(n8101) );
  nor2_1 U9176 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_mst_tx_flush), .ip2(
        i_i2c_U_DW_apb_i2c_sync_tx_empty_int_inv), .op(n7893) );
  nand2_1 U9177 ( .ip1(n8105), .ip2(i_i2c_ic_bus_idle), .op(n7892) );
  not_ab_or_c_or_d U9178 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_mst_tx_flush), .ip2(
        n8101), .ip3(n7893), .ip4(n7892), .op(n7894) );
  nand2_1 U9179 ( .ip1(n8121), .ip2(n7894), .op(n11090) );
  nor2_1 U9180 ( .ip1(n8113), .ip2(n11090), .op(n7902) );
  nand2_1 U9181 ( .ip1(n7895), .ip2(n8337), .op(n7899) );
  inv_1 U9182 ( .ip(n11021), .op(n11126) );
  nand2_1 U9183 ( .ip1(n11126), .ip2(
        i_i2c_U_DW_apb_i2c_sync_ic_10bit_mst_sync_inv), .op(n7898) );
  nand2_1 U9184 ( .ip1(n7896), .ip2(i_i2c_mst_debug_cstate[0]), .op(n7897) );
  nand4_1 U9185 ( .ip1(n7900), .ip2(n7899), .ip3(n7898), .ip4(n7897), .op(
        n7901) );
  or4_1 U9186 ( .ip1(n7904), .ip2(n7903), .ip3(n7902), .ip4(n7901), .op(n7906)
         );
  nor2_1 U9187 ( .ip1(n7905), .ip2(n9473), .op(n8112) );
  not_ab_or_c_or_d U9188 ( .ip1(n8109), .ip2(n8993), .ip3(n7906), .ip4(n8112), 
        .op(n7908) );
  nand2_1 U9189 ( .ip1(n11070), .ip2(n10926), .op(n7907) );
  nand4_1 U9190 ( .ip1(n7909), .ip2(n7908), .ip3(n11035), .ip4(n7907), .op(
        n7910) );
  not_ab_or_c_or_d U9191 ( .ip1(i_i2c_ic_bus_idle), .ip2(n5225), .ip3(
        i_i2c_start_en), .ip4(n7914), .op(n7915) );
  or2_1 U9192 ( .ip1(n7916), .ip2(n7915), .op(n7920) );
  ab_or_c_or_d U9193 ( .ip1(n7919), .ip2(n7918), .ip3(n7917), .ip4(n10926), 
        .op(n8967) );
  not_ab_or_c_or_d U9194 ( .ip1(n7921), .ip2(n7920), .ip3(n8109), .ip4(n8967), 
        .op(n5110) );
  nor2_1 U9195 ( .ip1(i_i2c_byte_wait_scl), .ip2(n7922), .op(n11863) );
  and2_1 U9196 ( .ip1(i_i2c_rx_scl_lcnt_en), .ip2(i_i2c_rx_scl_hcnt_en), .op(
        n7923) );
  nand2_1 U9197 ( .ip1(n7776), .ip2(n7923), .op(n7925) );
  nor2_1 U9198 ( .ip1(i_i2c_mst_rx_bit_count[3]), .ip2(n7925), .op(n7942) );
  nor2_1 U9199 ( .ip1(i_i2c_mst_rx_bit_count[2]), .ip2(
        i_i2c_mst_rx_bit_count[1]), .op(n7924) );
  inv_1 U9200 ( .ip(i_i2c_mst_rx_bit_count[0]), .op(n7926) );
  and2_1 U9201 ( .ip1(n7924), .ip2(n7926), .op(n11038) );
  nand2_1 U9202 ( .ip1(n11038), .ip2(i_i2c_mst_rx_bit_count[3]), .op(n8973) );
  or2_1 U9203 ( .ip1(n7925), .ip2(n8973), .op(n7944) );
  nand2_1 U9204 ( .ip1(n7944), .ip2(n11863), .op(n9314) );
  nor2_1 U9205 ( .ip1(n7942), .ip2(n9314), .op(n7936) );
  and2_1 U9206 ( .ip1(n7942), .ip2(n11863), .op(n10890) );
  nand2_1 U9207 ( .ip1(n10890), .ip2(n7926), .op(n10878) );
  inv_1 U9208 ( .ip(n10878), .op(n10882) );
  nor2_1 U9209 ( .ip1(n7936), .ip2(n10882), .op(n7938) );
  inv_1 U9210 ( .ip(i_i2c_mst_rx_bit_count[1]), .op(n10881) );
  nand2_1 U9211 ( .ip1(n10890), .ip2(n10881), .op(n7927) );
  nand2_1 U9212 ( .ip1(n7938), .ip2(n7927), .op(n7928) );
  nand2_1 U9213 ( .ip1(n7928), .ip2(i_i2c_mst_rx_bit_count[2]), .op(n7929) );
  and2_1 U9214 ( .ip1(i_i2c_mst_rx_bit_count[0]), .ip2(
        i_i2c_mst_rx_bit_count[1]), .op(n7940) );
  inv_1 U9215 ( .ip(i_i2c_mst_rx_bit_count[2]), .op(n10887) );
  nand3_1 U9216 ( .ip1(n10890), .ip2(n7940), .ip3(n10887), .op(n10884) );
  nand2_1 U9217 ( .ip1(n7929), .ip2(n10884), .op(n5107) );
  inv_1 U9218 ( .ip(n11038), .op(n11041) );
  nor2_1 U9219 ( .ip1(n11041), .ip2(n5591), .op(n7931) );
  nor2_1 U9220 ( .ip1(i_i2c_mst_rx_bit_count[3]), .ip2(n7776), .op(n7930) );
  nor2_1 U9221 ( .ip1(n7931), .ip2(n7930), .op(n7933) );
  nand2_1 U9222 ( .ip1(n7936), .ip2(n7933), .op(n9312) );
  inv_1 U9223 ( .ip(n9312), .op(n7932) );
  nand2_1 U9224 ( .ip1(n7932), .ip2(i_i2c_rx_scl_lcnt_en), .op(n7935) );
  inv_1 U9225 ( .ip(n11863), .op(n10876) );
  or2_1 U9226 ( .ip1(n10876), .ip2(n7933), .op(n7934) );
  nand2_1 U9227 ( .ip1(n7935), .ip2(n7934), .op(n5194) );
  nand2_1 U9228 ( .ip1(n7936), .ip2(i_i2c_mst_rx_bit_count[0]), .op(n7937) );
  nand2_1 U9229 ( .ip1(n7937), .ip2(n10878), .op(n5109) );
  nor2_1 U9230 ( .ip1(n7938), .ip2(n10881), .op(n7939) );
  and3_1 U9231 ( .ip1(n10890), .ip2(i_i2c_mst_rx_bit_count[0]), .ip3(n10881), 
        .op(n10888) );
  or2_1 U9232 ( .ip1(n7939), .ip2(n10888), .op(n5108) );
  and2_1 U9233 ( .ip1(n7940), .ip2(i_i2c_mst_rx_bit_count[2]), .op(n7941) );
  nand2_1 U9234 ( .ip1(n7942), .ip2(n7941), .op(n10875) );
  inv_1 U9235 ( .ip(n10875), .op(n9616) );
  nor2_1 U9236 ( .ip1(i_i2c_mst_rx_bit_count[3]), .ip2(n9616), .op(n7943) );
  nor2_1 U9237 ( .ip1(n9314), .ip2(n7943), .op(n5106) );
  nor2_1 U9238 ( .ip1(n10876), .ip2(n7944), .op(n4931) );
  inv_1 U9239 ( .ip(i_i2c_scl_lcnt_cmplt), .op(n11040) );
  or2_1 U9240 ( .ip1(n5591), .ip2(n11040), .op(n8976) );
  nand2_1 U9241 ( .ip1(n9312), .ip2(n8976), .op(n9313) );
  nand2_1 U9242 ( .ip1(n9313), .ip2(i_i2c_rx_scl_hcnt_en), .op(n7947) );
  inv_1 U9243 ( .ip(n8976), .op(n7945) );
  nand3_1 U9244 ( .ip1(n9312), .ip2(n6352), .ip3(n7945), .op(n7946) );
  nand2_1 U9245 ( .ip1(n7947), .ip2(n7946), .op(n7948) );
  and2_1 U9246 ( .ip1(n7948), .ip2(n11863), .op(n5195) );
  and2_1 U9247 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[0]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[1]), .op(n9067) );
  and2_1 U9248 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_data_scl_lcnt_en), .ip2(
        i_i2c_scl_hcnt_en), .op(n7949) );
  nand2_1 U9249 ( .ip1(n7776), .ip2(n7949), .op(n9322) );
  nor2_1 U9250 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[3]), .ip2(n9322), .op(n9618) );
  nand3_1 U9251 ( .ip1(n11834), .ip2(n9618), .ip3(i_i2c_debug_wr), .op(n7955)
         );
  nor2_1 U9252 ( .ip1(n9067), .ip2(n7955), .op(n7954) );
  inv_1 U9253 ( .ip(i_i2c_debug_wr), .op(n7950) );
  nand2_1 U9254 ( .ip1(n11834), .ip2(n7950), .op(n10947) );
  nor2_1 U9255 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[1]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[0]), .op(n7951) );
  inv_1 U9256 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[2]), .op(n9068)
         );
  nand2_1 U9257 ( .ip1(n7951), .ip2(n9068), .op(n11046) );
  and2_1 U9258 ( .ip1(n11046), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[3]), .op(n8156) );
  nand2_1 U9259 ( .ip1(n11834), .ip2(n8156), .op(n7952) );
  and2_1 U9260 ( .ip1(n10947), .ip2(n7952), .op(n8154) );
  nand2_1 U9261 ( .ip1(n11834), .ip2(n9322), .op(n7953) );
  nand2_1 U9262 ( .ip1(n8154), .ip2(n7953), .op(n8149) );
  or2_1 U9263 ( .ip1(n7954), .ip2(n8149), .op(n8146) );
  inv_1 U9264 ( .ip(n7955), .op(n8151) );
  nand2_1 U9265 ( .ip1(n8151), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[0]), .op(n7956) );
  inv_1 U9266 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[1]), .op(n9064)
         );
  nand2_1 U9267 ( .ip1(n7956), .ip2(n9064), .op(n7957) );
  and2_1 U9268 ( .ip1(n8146), .ip2(n7957), .op(n4139) );
  inv_1 U9269 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_3_), .op(
        n9560) );
  nand2_1 U9270 ( .ip1(n11835), .ip2(n9560), .op(n8044) );
  inv_1 U9271 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[0]), .op(
        n11304) );
  inv_1 U9272 ( .ip(i_i2c_slv_rxbyte_rdy), .op(n11673) );
  nor2_1 U9273 ( .ip1(n11673), .ip2(n11083), .op(n10871) );
  inv_1 U9274 ( .ip(i_i2c_slv_debug_cstate[0]), .op(n7958) );
  nor2_1 U9275 ( .ip1(n7958), .ip2(n9592), .op(n11289) );
  inv_1 U9276 ( .ip(i_i2c_slv_debug_cstate[2]), .op(n9594) );
  nand2_1 U9277 ( .ip1(n11289), .ip2(n9594), .op(n9590) );
  or2_1 U9278 ( .ip1(n10871), .ip2(n9590), .op(n11299) );
  inv_1 U9279 ( .ip(n11299), .op(n11305) );
  nor2_1 U9280 ( .ip1(n7959), .ip2(n9585), .op(n11288) );
  inv_1 U9281 ( .ip(n11288), .op(n8136) );
  nand2_1 U9282 ( .ip1(n11289), .ip2(i_i2c_slv_debug_cstate[2]), .op(n11296)
         );
  nand2_1 U9283 ( .ip1(n8136), .ip2(n11296), .op(n7960) );
  nor2_1 U9284 ( .ip1(i_i2c_slv_rxbyte_rdy), .ip2(n11083), .op(n11235) );
  and2_1 U9285 ( .ip1(n7960), .ip2(n11235), .op(n11301) );
  or2_1 U9286 ( .ip1(n11305), .ip2(n11301), .op(n11311) );
  inv_1 U9287 ( .ip(n11311), .op(n11669) );
  nor2_1 U9288 ( .ip1(n11304), .ip2(n8044), .op(n9604) );
  not_ab_or_c_or_d U9289 ( .ip1(n8044), .ip2(n11304), .ip3(n11669), .ip4(n9604), .op(n4169) );
  nor2_1 U9290 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[1]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[2]), .op(n7961) );
  nand4_1 U9291 ( .ip1(n11305), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[3]), .ip3(n7961), .ip4(
        n11304), .op(n11312) );
  and3_1 U9292 ( .ip1(n11312), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[3]), .ip3(n11311), .op(
        n5074) );
  nand2_1 U9293 ( .ip1(i_i2c_tx_push), .ip2(i_i2c_tx_full), .op(n10195) );
  and4_1 U9294 ( .ip1(i_i2c_tx_push), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[1]), .ip3(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[0]), .ip4(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[2]), .op(n7962) );
  nor2_1 U9295 ( .ip1(i_i2c_tx_full), .ip2(n7962), .op(n7963) );
  not_ab_or_c_or_d U9296 ( .ip1(i_i2c_tx_pop_sync), .ip2(n10195), .ip3(n7963), 
        .ip4(n11026), .op(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N37) );
  nor2_1 U9297 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[0]), .ip2(n7964), 
        .op(n7965) );
  nor2_1 U9298 ( .ip1(n7966), .ip2(n7965), .op(n7967) );
  xor2_1 U9299 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_wrdc_tx_unconn[1]), .ip2(n7967), 
        .op(n11029) );
  and2_1 U9300 ( .ip1(i_i2c_tx_fifo_rst_n), .ip2(n11029), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N48) );
  or4_1 U9301 ( .ip1(n11867), .ip2(n11866), .ip3(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N37), .ip4(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N48), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N33) );
  or2_1 U9302 ( .ip1(i_i2c_ic_enable_sync), .ip2(i_i2c_slv_activity), .op(
        n7968) );
  nand2_1 U9303 ( .ip1(n7968), .ip2(i_i2c_ic_slave_en_sync), .op(n11236) );
  nor2_1 U9304 ( .ip1(n11236), .ip2(n7969), .op(i_i2c_U_DW_apb_i2c_slvfsm_N39)
         );
  inv_1 U9305 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[2]), .op(
        n8025) );
  inv_1 U9306 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[0]), 
        .op(n7970) );
  nand2_1 U9307 ( .ip1(n9560), .ip2(i_i2c_sda_vld), .op(n8004) );
  nor2_1 U9308 ( .ip1(n8004), .ip2(n11835), .op(n8041) );
  inv_1 U9309 ( .ip(n8041), .op(n7973) );
  nor2_1 U9310 ( .ip1(n7970), .ip2(n7973), .op(n9506) );
  inv_1 U9311 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[1]), 
        .op(n9505) );
  nand2_1 U9312 ( .ip1(n9505), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[2]), .op(n7974) );
  inv_1 U9313 ( .ip(n7974), .op(n7977) );
  nand2_1 U9314 ( .ip1(n9506), .ip2(n7977), .op(n7972) );
  inv_1 U9315 ( .ip(n11833), .op(n8096) );
  nand2_1 U9316 ( .ip1(n8096), .ip2(n9506), .op(n9507) );
  nor2_1 U9317 ( .ip1(n7974), .ip2(n9507), .op(n7971) );
  not_ab_or_c_or_d U9318 ( .ip1(n8025), .ip2(n7972), .ip3(n11669), .ip4(n7971), 
        .op(n5071) );
  or2_1 U9319 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[0]), 
        .ip2(n7973), .op(n9511) );
  nor2_1 U9320 ( .ip1(n11833), .ip2(n9511), .op(n9515) );
  nor2_1 U9321 ( .ip1(n7974), .ip2(n9511), .op(n7975) );
  nor2_1 U9322 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[3]), .ip2(
        n7975), .op(n7976) );
  not_ab_or_c_or_d U9323 ( .ip1(n7977), .ip2(n9515), .ip3(n11669), .ip4(n7976), 
        .op(n5070) );
  inv_1 U9324 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[0]), .op(
        n9554) );
  nand2_1 U9325 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[2]), 
        .ip2(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[1]), .op(n7980)
         );
  inv_1 U9326 ( .ip(n7980), .op(n7983) );
  nand2_1 U9327 ( .ip1(n9506), .ip2(n7983), .op(n7979) );
  nor2_1 U9328 ( .ip1(n7980), .ip2(n9507), .op(n7978) );
  not_ab_or_c_or_d U9329 ( .ip1(n9554), .ip2(n7979), .ip3(n11669), .ip4(n7978), 
        .op(n5073) );
  nor2_1 U9330 ( .ip1(n7980), .ip2(n9511), .op(n7981) );
  nor2_1 U9331 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[1]), .ip2(
        n7981), .op(n7982) );
  not_ab_or_c_or_d U9332 ( .ip1(n7983), .ip2(n9515), .ip3(n11669), .ip4(n7982), 
        .op(n5072) );
  inv_1 U9333 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[4]), .op(
        n7986) );
  inv_1 U9334 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[2]), 
        .op(n9504) );
  nand2_1 U9335 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[1]), 
        .ip2(n9504), .op(n7987) );
  inv_1 U9336 ( .ip(n7987), .op(n7990) );
  nand2_1 U9337 ( .ip1(n9506), .ip2(n7990), .op(n7985) );
  nor2_1 U9338 ( .ip1(n7987), .ip2(n9507), .op(n7984) );
  not_ab_or_c_or_d U9339 ( .ip1(n7986), .ip2(n7985), .ip3(n11669), .ip4(n7984), 
        .op(n5069) );
  nor2_1 U9340 ( .ip1(n7987), .ip2(n9511), .op(n7988) );
  nor2_1 U9341 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[5]), .ip2(
        n7988), .op(n7989) );
  not_ab_or_c_or_d U9342 ( .ip1(n7990), .ip2(n9515), .ip3(n11669), .ip4(n7989), 
        .op(n5068) );
  inv_1 U9343 ( .ip(i_i2c_ic_10bit_slv), .op(n11868) );
  nor4_1 U9344 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[1]), 
        .ip2(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[2]), .ip3(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_bit_count_2to0[0]), .ip4(n9560), 
        .op(n8037) );
  and2_1 U9345 ( .ip1(n11288), .ip2(n8037), .op(n8019) );
  inv_1 U9346 ( .ip(n8037), .op(n7991) );
  nor2_1 U9347 ( .ip1(n7991), .ip2(n11299), .op(n8038) );
  nor2_1 U9348 ( .ip1(n8019), .ip2(n8038), .op(n8045) );
  xor2_1 U9349 ( .ip1(i_i2c_ic_sar[8]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[1]), .op(n7992) );
  nand4_1 U9350 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[5]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[4]), .ip3(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[6]), .ip4(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[7]), .op(n8021) );
  or2_1 U9351 ( .ip1(n8021), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[3]), .op(n9541) );
  nor2_1 U9352 ( .ip1(n7992), .ip2(n9541), .op(n7995) );
  nor2_1 U9353 ( .ip1(n8025), .ip2(i_i2c_ic_sar[9]), .op(n7993) );
  not_ab_or_c_or_d U9354 ( .ip1(i_i2c_ic_sar[9]), .ip2(n8025), .ip3(n7993), 
        .ip4(n11868), .op(n7994) );
  nand2_1 U9355 ( .ip1(n7995), .ip2(n7994), .op(n8003) );
  nor2_1 U9356 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[6]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[4]), .op(n7999) );
  inv_1 U9357 ( .ip(n7999), .op(n7998) );
  inv_1 U9358 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[5]), .op(
        n7996) );
  inv_1 U9359 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[7]), .op(
        n8026) );
  nand3_1 U9360 ( .ip1(n7996), .ip2(n8026), .ip3(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[3]), .op(n7997) );
  nor2_1 U9361 ( .ip1(n7998), .ip2(n7997), .op(n9517) );
  nor3_1 U9362 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[3]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[7]), .ip3(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[1]), .op(n8001) );
  nor2_1 U9363 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[5]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[2]), .op(n8000) );
  and3_1 U9364 ( .ip1(n8001), .ip2(n8000), .ip3(n7999), .op(n9555) );
  nor2_1 U9365 ( .ip1(n9517), .ip2(n9555), .op(n8002) );
  nand2_1 U9366 ( .ip1(n8038), .ip2(n8002), .op(n8020) );
  or2_1 U9367 ( .ip1(n8003), .ip2(n8020), .op(n9544) );
  or2_1 U9368 ( .ip1(n11078), .ip2(n9544), .op(n9536) );
  and2_1 U9369 ( .ip1(n8004), .ip2(i_i2c_rx_slv_read), .op(n8005) );
  inv_1 U9370 ( .ip(n8038), .op(n8042) );
  mux2_1 U9371 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[0]), .ip2(
        n8005), .s(n8042), .op(n11238) );
  or2_1 U9372 ( .ip1(n11238), .ip2(n9544), .op(n8006) );
  nand2_1 U9373 ( .ip1(n9536), .ip2(n8006), .op(n8036) );
  inv_1 U9374 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[6]), .op(
        n9510) );
  mux2_1 U9375 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[6]), .ip2(
        n9510), .s(i_i2c_ic_sar[6]), .op(n8017) );
  mux2_1 U9376 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[7]), .ip2(
        n8026), .s(i_i2c_ic_sar[7]), .op(n8016) );
  xor2_1 U9377 ( .ip1(i_i2c_ic_sar[5]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[5]), .op(n8010) );
  xor2_1 U9378 ( .ip1(i_i2c_ic_sar[4]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[4]), .op(n8009) );
  xor2_1 U9379 ( .ip1(i_i2c_ic_sar[1]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[1]), .op(n8008) );
  xor2_1 U9380 ( .ip1(i_i2c_ic_sar[2]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[2]), .op(n8007) );
  nor4_1 U9381 ( .ip1(n8010), .ip2(n8009), .ip3(n8008), .ip4(n8007), .op(n8014) );
  xor2_1 U9382 ( .ip1(i_i2c_ic_sar[3]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[3]), .op(n8012) );
  xor2_1 U9383 ( .ip1(i_i2c_ic_sar[0]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[0]), .op(n8011) );
  nor3_1 U9384 ( .ip1(n11868), .ip2(n8012), .ip3(n8011), .op(n8013) );
  nand2_1 U9385 ( .ip1(n8014), .ip2(n8013), .op(n8015) );
  nor3_1 U9386 ( .ip1(n8017), .ip2(n8016), .ip3(n8015), .op(n8018) );
  nand2_1 U9387 ( .ip1(n8019), .ip2(n8018), .op(n8043) );
  nor2_1 U9388 ( .ip1(i_i2c_ic_10bit_slv), .ip2(n8020), .op(n9543) );
  xor2_1 U9389 ( .ip1(i_i2c_ic_sar[4]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[5]), .op(n8034) );
  xor2_1 U9390 ( .ip1(i_i2c_ic_sar[3]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[4]), .op(n8033) );
  inv_1 U9391 ( .ip(i_i2c_ic_sar[2]), .op(n8022) );
  nand2_1 U9392 ( .ip1(n8021), .ip2(n8022), .op(n8023) );
  mux2_1 U9393 ( .ip1(n8023), .ip2(n8022), .s(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[3]), .op(n8032) );
  inv_1 U9394 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[1]), .op(
        n8024) );
  mux2_1 U9395 ( .ip1(n8024), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[1]), .s(i_i2c_ic_sar[0]), 
        .op(n8030) );
  mux2_1 U9396 ( .ip1(n8025), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[2]), .s(i_i2c_ic_sar[1]), 
        .op(n8029) );
  mux2_1 U9397 ( .ip1(n9510), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[6]), .s(i_i2c_ic_sar[5]), 
        .op(n8028) );
  mux2_1 U9398 ( .ip1(n8026), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[7]), .s(i_i2c_ic_sar[6]), 
        .op(n8027) );
  nand4_1 U9399 ( .ip1(n8030), .ip2(n8029), .ip3(n8028), .ip4(n8027), .op(
        n8031) );
  nor4_1 U9400 ( .ip1(n8034), .ip2(n8033), .ip3(n8032), .ip4(n8031), .op(n8035) );
  nand2_1 U9401 ( .ip1(n9543), .ip2(n8035), .op(n9546) );
  nand2_1 U9402 ( .ip1(n8043), .ip2(n9546), .op(n9538) );
  not_ab_or_c_or_d U9403 ( .ip1(n8037), .ip2(n8045), .ip3(n8036), .ip4(n9538), 
        .op(n8040) );
  nand4_1 U9404 ( .ip1(n8038), .ip2(n9555), .ip3(
        i_i2c_ic_ack_general_call_sync), .ip4(n9554), .op(n8039) );
  nand2_1 U9405 ( .ip1(n8040), .ip2(n8039), .op(n8047) );
  nor2_1 U9406 ( .ip1(n11669), .ip2(n8041), .op(n9553) );
  nor2_1 U9407 ( .ip1(n8042), .ip2(n11835), .op(n9556) );
  nor2_1 U9408 ( .ip1(n8043), .ip2(n11835), .op(n9550) );
  not_ab_or_c_or_d U9409 ( .ip1(n8045), .ip2(n8044), .ip3(n9556), .ip4(n9550), 
        .op(n8046) );
  nand2_1 U9410 ( .ip1(n9553), .ip2(n8046), .op(n8048) );
  nand3_1 U9411 ( .ip1(n8047), .ip2(n11311), .ip3(n8048), .op(n8051) );
  inv_1 U9412 ( .ip(n8048), .op(n8049) );
  nand2_1 U9413 ( .ip1(n8049), .ip2(i_i2c_slv_rx_ack_vld), .op(n8050) );
  nand2_1 U9414 ( .ip1(n8051), .ip2(n8050), .op(n5082) );
  and2_1 U9415 ( .ip1(i_i2c_slv_rx_ack_vld), .ip2(
        i_i2c_U_DW_apb_i2c_slvfsm_ic_enable_sync_vld), .op(n8138) );
  or2_1 U9416 ( .ip1(i_i2c_ic_enable_sync), .ip2(n8138), .op(n5081) );
  nand3_1 U9417 ( .ip1(n11068), .ip2(i_i2c_U_DW_apb_i2c_mstfsm_old_is_read), 
        .ip3(i_i2c_U_DW_apb_i2c_mstfsm_N487), .op(n8052) );
  nand2_1 U9418 ( .ip1(n8052), .ip2(n11021), .op(n5201) );
  inv_1 U9419 ( .ip(i_i2c_U_DW_apb_i2c_mstfsm_byte_waiting_q), .op(n8064) );
  inv_1 U9420 ( .ip(n8058), .op(n9502) );
  nor2_1 U9421 ( .ip1(n9502), .ip2(n8987), .op(n8966) );
  inv_1 U9422 ( .ip(n8053), .op(n8988) );
  and2_1 U9423 ( .ip1(n8988), .ip2(n8989), .op(n8059) );
  nand2_1 U9424 ( .ip1(n8966), .ip2(n8059), .op(n8063) );
  nand2_1 U9425 ( .ip1(n10932), .ip2(n8126), .op(n8054) );
  nand2_1 U9426 ( .ip1(n8054), .ip2(i_i2c_U_DW_apb_i2c_sync_tx_empty_int_inv), 
        .op(n8057) );
  nand3_1 U9427 ( .ip1(n11126), .ip2(i_i2c_U_DW_apb_i2c_mstfsm_byte_waiting_q), 
        .ip3(n8055), .op(n8056) );
  nand3_1 U9428 ( .ip1(n8058), .ip2(n8057), .ip3(n8056), .op(n8061) );
  inv_1 U9429 ( .ip(n8059), .op(n8060) );
  nor3_1 U9430 ( .ip1(n8061), .ip2(n8987), .ip3(n8060), .op(n8062) );
  not_ab_or_c_or_d U9431 ( .ip1(n8064), .ip2(n8063), .ip3(n8062), .ip4(n8121), 
        .op(n5184) );
  nand2_1 U9432 ( .ip1(n6352), .ip2(n8065), .op(n11045) );
  inv_1 U9433 ( .ip(i_i2c_mst_tx_ack_vld), .op(n8067) );
  nor2_1 U9434 ( .ip1(n11045), .ip2(n8096), .op(n8066) );
  not_ab_or_c_or_d U9435 ( .ip1(n8068), .ip2(n11045), .ip3(n8067), .ip4(n8066), 
        .op(n4161) );
  inv_1 U9436 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly1), .op(n9055)
         );
  inv_1 U9437 ( .ip(n11859), .op(n9497) );
  nor2_1 U9438 ( .ip1(n9055), .ip2(n9497), .op(n11860) );
  and2_1 U9439 ( .ip1(n11859), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly2), .op(
        i_i2c_U_DW_apb_i2c_tx_shift_N402) );
  inv_1 U9440 ( .ip(n11045), .op(n8070) );
  nor2_1 U9441 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_q), .ip2(n11835), 
        .op(n8069) );
  nor2_1 U9442 ( .ip1(n8070), .ip2(n8069), .op(n4170) );
  inv_1 U9443 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[0]), .op(
        n9052) );
  inv_1 U9444 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_q), .op(n8071) );
  nor2_1 U9445 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_scl_is_low_qq), .ip2(n8071), 
        .op(n8074) );
  and2_1 U9446 ( .ip1(n8072), .ip2(i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv), 
        .op(n8073) );
  mux2_1 U9447 ( .ip1(n8074), .ip2(n11835), .s(n8073), .op(n9037) );
  nand2_1 U9448 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly1), .ip2(
        i_i2c_slv_tx_ready_unconn), .op(n8087) );
  nor2_1 U9449 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[3]), .ip2(
        n8087), .op(n8075) );
  nand2_1 U9450 ( .ip1(n9037), .ip2(n8075), .op(n8077) );
  nor2_1 U9451 ( .ip1(n9052), .ip2(n8077), .op(n8078) );
  nor2_1 U9452 ( .ip1(n9497), .ip2(n8078), .op(n8082) );
  nand2_1 U9453 ( .ip1(n8077), .ip2(n9052), .op(n8076) );
  and2_1 U9454 ( .ip1(n8082), .ip2(n8076), .op(n5101) );
  nand2_1 U9455 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[0]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[1]), .op(n9047) );
  nor2_1 U9456 ( .ip1(n9047), .ip2(n8077), .op(n8080) );
  nor2_1 U9457 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[1]), .ip2(
        n8078), .op(n8079) );
  nor3_1 U9458 ( .ip1(n8080), .ip2(n9497), .ip3(n8079), .op(n5100) );
  nor2_1 U9459 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[2]), .ip2(
        n8080), .op(n8081) );
  ab_or_c_or_d U9460 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[2]), 
        .ip2(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[1]), .ip3(n9497), 
        .ip4(n8081), .op(n8084) );
  nand2_1 U9461 ( .ip1(n8082), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[2]), .op(n8083) );
  nand2_1 U9462 ( .ip1(n8084), .ip2(n8083), .op(n5099) );
  inv_1 U9463 ( .ip(n9047), .op(n9046) );
  and3_1 U9464 ( .ip1(n9037), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[2]), .ip3(n9046), .op(
        n9620) );
  nand3_1 U9465 ( .ip1(n9620), .ip2(i_i2c_slv_tx_ready_unconn), .ip3(n11860), 
        .op(n8086) );
  nand2_1 U9466 ( .ip1(n11859), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[3]), .op(n8085) );
  nand2_1 U9467 ( .ip1(n8086), .ip2(n8085), .op(n5098) );
  or2_1 U9468 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[0]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[1]), .op(n9049) );
  or2_1 U9469 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[2]), .ip2(
        n9049), .op(n9039) );
  inv_1 U9470 ( .ip(n9039), .op(n8089) );
  inv_1 U9471 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[3]), .op(
        n9619) );
  nor2_1 U9472 ( .ip1(n9619), .ip2(n8087), .op(n8088) );
  and2_1 U9473 ( .ip1(n8089), .ip2(n8088), .op(n9041) );
  and2_1 U9474 ( .ip1(n11859), .ip2(n9041), .op(n8090) );
  nor2_1 U9475 ( .ip1(i_i2c_slv_tx_ack_vld), .ip2(n9041), .op(n8092) );
  nor2_1 U9476 ( .ip1(n8092), .ip2(n9497), .op(n5104) );
  inv_1 U9477 ( .ip(i_i2c_slv_ack_det), .op(n8093) );
  nor2_1 U9478 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_scl_edg_hl_q), .ip2(n8093), 
        .op(n8095) );
  nand2_1 U9479 ( .ip1(i_i2c_slv_tx_ack_vld), .ip2(i_i2c_sda_vld), .op(n8094)
         );
  mux2_1 U9480 ( .ip1(n8096), .ip2(n8095), .s(n8094), .op(n5065) );
  nand2_1 U9481 ( .ip1(n11127), .ip2(i_i2c_ic_enable_sync), .op(n8123) );
  nand2_1 U9482 ( .ip1(n10871), .ip2(i_i2c_ic_data_oe), .op(n8097) );
  or2_1 U9483 ( .ip1(n8097), .ip2(n9590), .op(n9572) );
  nor2_1 U9484 ( .ip1(i_i2c_rx_gen_call), .ip2(n9572), .op(n11230) );
  and2_1 U9485 ( .ip1(i_i2c_rx_addr_match), .ip2(i_i2c_rx_slv_read), .op(n8098) );
  and2_1 U9486 ( .ip1(n11230), .ip2(n8098), .op(n10142) );
  nor4_1 U9487 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_N487), .ip2(n11861), .ip3(
        n8099), .ip4(n10142), .op(n8103) );
  nor2_1 U9488 ( .ip1(i_i2c_U_DW_apb_i2c_sync_tx_empty_int_inv), .ip2(n9567), 
        .op(n8100) );
  nor2_1 U9489 ( .ip1(n8100), .ip2(n10142), .op(n11318) );
  inv_1 U9490 ( .ip(n11318), .op(n11319) );
  nor2_1 U9491 ( .ip1(n8101), .ip2(n11319), .op(n8102) );
  nor2_1 U9492 ( .ip1(n8103), .ip2(n8102), .op(n8104) );
  nor2_1 U9493 ( .ip1(n8123), .ip2(n8104), .op(n5029) );
  inv_1 U9494 ( .ip(i_i2c_mst_activity), .op(n11017) );
  not_ab_or_c_or_d U9495 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_sync_d), 
        .ip2(n11017), .ip3(n8105), .ip4(i_i2c_U_DW_apb_i2c_mstfsm_N487), .op(
        n11054) );
  inv_1 U9496 ( .ip(n11054), .op(n8107) );
  nand2_1 U9497 ( .ip1(n11127), .ip2(i_i2c_U_DW_apb_i2c_mstfsm_abrt_in_idle), 
        .op(n8106) );
  nand2_1 U9498 ( .ip1(n8107), .ip2(n8106), .op(n5197) );
  inv_1 U9499 ( .ip(n8108), .op(n11076) );
  nor2_1 U9500 ( .ip1(n10943), .ip2(n8109), .op(n8333) );
  nand2_1 U9501 ( .ip1(n11068), .ip2(n8333), .op(n8110) );
  nand2_1 U9502 ( .ip1(n8111), .ip2(n8110), .op(n8117) );
  inv_1 U9503 ( .ip(n8985), .op(n11096) );
  not_ab_or_c_or_d U9504 ( .ip1(n11096), .ip2(i_i2c_U_DW_apb_i2c_mstfsm_N487), 
        .ip3(n11054), .ip4(n11061), .op(n8116) );
  inv_1 U9505 ( .ip(n8112), .op(n8115) );
  inv_1 U9506 ( .ip(n11090), .op(n8114) );
  nand2_1 U9507 ( .ip1(n8114), .ip2(n8113), .op(n11093) );
  not_ab_or_c_or_d U9508 ( .ip1(n8119), .ip2(n10145), .ip3(n11076), .ip4(n8118), .op(n10147) );
  nor2_1 U9509 ( .ip1(n8121), .ip2(n10147), .op(n8120) );
  not_ab_or_c_or_d U9510 ( .ip1(n8121), .ip2(
        i_i2c_U_DW_apb_i2c_mstfsm_abrt_in_idle), .ip3(
        i_i2c_U_DW_apb_i2c_mstfsm_mst_tx_flush), .ip4(n8120), .op(n8122) );
  nor3_1 U9511 ( .ip1(n11319), .ip2(n8123), .ip3(n8122), .op(n4857) );
  inv_1 U9512 ( .ip(i_i2c_ic_rstrt_en), .op(
        i_i2c_U_DW_apb_i2c_sync_U_ic_rstrt_en_1_sync_N2) );
  nand3_1 U9513 ( .ip1(n10147), .ip2(
        i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_chk_win), .ip3(n10875), .op(n8125)
         );
  nand2_1 U9514 ( .ip1(n9616), .ip2(i_i2c_ic_abort_sync), .op(n8124) );
  nand2_1 U9515 ( .ip1(n8125), .ip2(n8124), .op(n4174) );
  nor2_1 U9516 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(n8126), .op(n11858) );
  inv_1 U9517 ( .ip(i_i2c_mst_rx_ack_vld), .op(n8127) );
  nor2_1 U9518 ( .ip1(i_i2c_scl_lcnt_cmplt), .ip2(i_i2c_mst_rx_bit_count[3]), 
        .op(n11037) );
  nor2_1 U9519 ( .ip1(n8127), .ip2(n11037), .op(n8129) );
  nor2_1 U9520 ( .ip1(n8973), .ip2(n5591), .op(n8128) );
  nor2_1 U9521 ( .ip1(n8129), .ip2(n8128), .op(n8130) );
  nor2_1 U9522 ( .ip1(n10876), .ip2(n8130), .op(n8131) );
  or2_1 U9523 ( .ip1(n8131), .ip2(n4931), .op(n4952) );
  inv_1 U9524 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_data_scl_lcnt_en), .op(n8132)
         );
  inv_1 U9525 ( .ip(n11834), .op(n8141) );
  nor2_1 U9526 ( .ip1(n8132), .ip2(n8141), .op(n8144) );
  nand3_1 U9527 ( .ip1(i_i2c_scl_lcnt_cmplt), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_data_scl_lcnt_en), .ip3(i_i2c_scl_hcnt_en), 
        .op(n8133) );
  nand2_1 U9528 ( .ip1(n5591), .ip2(n8133), .op(n8157) );
  inv_1 U9529 ( .ip(n11046), .op(n11047) );
  nand4_1 U9530 ( .ip1(n8157), .ip2(n11047), .ip3(i_i2c_debug_wr), .ip4(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[3]), .op(n8134) );
  nor2_1 U9531 ( .ip1(n8134), .ip2(n8141), .op(n8982) );
  and2_1 U9532 ( .ip1(i_i2c_U_DW_apb_i2c_mstfsm_mst_gen_ack_en_r), .ip2(
        i_i2c_mst_rx_ack_vld), .op(n8135) );
  nand2_1 U9533 ( .ip1(n11858), .ip2(n8135), .op(n8140) );
  and2_1 U9534 ( .ip1(n8136), .ip2(n9590), .op(n11244) );
  nand2_1 U9535 ( .ip1(n11289), .ip2(n9583), .op(n8137) );
  nand2_1 U9536 ( .ip1(n11244), .ip2(n8137), .op(n9080) );
  nand2_1 U9537 ( .ip1(n9080), .ip2(n8138), .op(n8139) );
  and2_1 U9538 ( .ip1(n8140), .ip2(n8139), .op(n9470) );
  inv_1 U9539 ( .ip(n9470), .op(n9336) );
  inv_1 U9540 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[3]), .op(n8977)
         );
  nand3_1 U9541 ( .ip1(n8145), .ip2(i_i2c_debug_wr), .ip3(n8977), .op(n9320)
         );
  not_ab_or_c_or_d U9542 ( .ip1(n11040), .ip2(n9336), .ip3(n9320), .ip4(n8141), 
        .op(n8142) );
  nor3_1 U9543 ( .ip1(n8982), .ip2(n8142), .ip3(n8151), .op(n8143) );
  mux2_1 U9544 ( .ip1(n8145), .ip2(n8144), .s(n8143), .op(n4141) );
  mux2_1 U9545 ( .ip1(n8151), .ip2(n8149), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[0]), .op(n4140) );
  nand2_1 U9546 ( .ip1(n8146), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[2]), .op(n8148) );
  nand3_1 U9547 ( .ip1(n8151), .ip2(n9067), .ip3(n9068), .op(n8147) );
  nand2_1 U9548 ( .ip1(n8148), .ip2(n8147), .op(n4138) );
  nand2_1 U9549 ( .ip1(n8149), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[3]), .op(n8153) );
  inv_1 U9550 ( .ip(n9067), .op(n8150) );
  nor2_1 U9551 ( .ip1(n9068), .ip2(n8150), .op(n9617) );
  nand2_1 U9552 ( .ip1(n8151), .ip2(n9617), .op(n8152) );
  nand2_1 U9553 ( .ip1(n8153), .ip2(n8152), .op(n4137) );
  inv_1 U9554 ( .ip(n8154), .op(n8155) );
  nand2_1 U9555 ( .ip1(n8155), .ip2(i_i2c_scl_hcnt_en), .op(n8164) );
  nor2_1 U9556 ( .ip1(n8156), .ip2(n8976), .op(n9325) );
  inv_1 U9557 ( .ip(n9325), .op(n8158) );
  nand2_1 U9558 ( .ip1(n8158), .ip2(n8157), .op(n8159) );
  nand2_1 U9559 ( .ip1(n8159), .ip2(i_i2c_scl_hcnt_en), .op(n8161) );
  nand3_1 U9560 ( .ip1(n9325), .ip2(n6352), .ip3(i_i2c_debug_wr), .op(n8160)
         );
  nand2_1 U9561 ( .ip1(n8161), .ip2(n8160), .op(n8162) );
  nand2_1 U9562 ( .ip1(n8162), .ip2(n11834), .op(n8163) );
  nand2_1 U9563 ( .ip1(n8164), .ip2(n8163), .op(n4142) );
  nand2_1 U9564 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[4]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[5]), .op(n8290) );
  nand2_1 U9565 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[1]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[2]), .op(n8289) );
  nor2_1 U9566 ( .ip1(n8188), .ip2(n8186), .op(n8174) );
  inv_1 U9567 ( .ip(n8174), .op(n8169) );
  nor2_1 U9568 ( .ip1(n8169), .ip2(n8189), .op(n8170) );
  nand2_1 U9569 ( .ip1(n5267), .ip2(n8170), .op(n8171) );
  xnor2_1 U9570 ( .ip1(n8172), .ip2(n8171), .op(n8197) );
  nand2_1 U9571 ( .ip1(n8174), .ip2(n8173), .op(n8175) );
  nor2_1 U9572 ( .ip1(n8175), .ip2(n8189), .op(n8176) );
  nand2_1 U9573 ( .ip1(n5267), .ip2(n8176), .op(n8177) );
  xnor2_1 U9574 ( .ip1(n8178), .ip2(n8177), .op(n8181) );
  inv_1 U9575 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[15]), .op(n8179)
         );
  nand2_1 U9576 ( .ip1(n8181), .ip2(n8179), .op(n8198) );
  inv_1 U9577 ( .ip(n8198), .op(n8180) );
  nor3_1 U9578 ( .ip1(n8196), .ip2(n8197), .ip3(n8180), .op(n8183) );
  nor2_1 U9579 ( .ip1(n8181), .ip2(n8179), .op(n8182) );
  nand2_1 U9580 ( .ip1(n5267), .ip2(n8184), .op(n8185) );
  inv_1 U9581 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[12]), .op(n8270)
         );
  inv_1 U9582 ( .ip(n8189), .op(n8190) );
  nand2_1 U9583 ( .ip1(n5267), .ip2(n8190), .op(n8191) );
  xnor2_1 U9584 ( .ip1(n8188), .ip2(n8191), .op(n8271) );
  nor2_1 U9585 ( .ip1(n8192), .ip2(n8193), .op(n8195) );
  nor2_1 U9586 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[13]), .ip2(
        n5460), .op(n8194) );
  or2_1 U9587 ( .ip1(n8195), .ip2(n8194), .op(n8200) );
  nand2_1 U9588 ( .ip1(n8197), .ip2(n8196), .op(n8199) );
  nand2_1 U9589 ( .ip1(n8199), .ip2(n8198), .op(n8269) );
  nor2_1 U9590 ( .ip1(n5454), .ip2(n8203), .op(n8206) );
  nand2_1 U9591 ( .ip1(n5454), .ip2(n8203), .op(n8204) );
  inv_1 U9592 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[4]), .op(n8240)
         );
  inv_1 U9593 ( .ip(n8215), .op(n8212) );
  nand2_1 U9594 ( .ip1(n5261), .ip2(n8212), .op(n8213) );
  xor2_1 U9595 ( .ip1(n5261), .ip2(n8215), .op(n8239) );
  nor2_1 U9596 ( .ip1(n8219), .ip2(n5468), .op(n8218) );
  nand2_1 U9597 ( .ip1(n5561), .ip2(n8219), .op(n8221) );
  nand2_1 U9598 ( .ip1(n5468), .ip2(n8219), .op(n8220) );
  xnor2_1 U9599 ( .ip1(n5469), .ip2(n5561), .op(n8231) );
  inv_1 U9600 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[2]), .op(n8233)
         );
  xnor2_1 U9601 ( .ip1(n8229), .ip2(n5464), .op(n8228) );
  inv_1 U9602 ( .ip(n8228), .op(n8230) );
  nor3_1 U9603 ( .ip1(n8233), .ip2(n8232), .ip3(n8231), .op(n8234) );
  not_ab_or_c_or_d U9604 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[3]), 
        .ip2(n8236), .ip3(n8235), .ip4(n8234), .op(n8237) );
  ab_or_c_or_d U9605 ( .ip1(n8240), .ip2(n8239), .ip3(n8238), .ip4(n8237), 
        .op(n8241) );
  inv_1 U9606 ( .ip(n8247), .op(n8243) );
  nor2_1 U9607 ( .ip1(n5459), .ip2(n8243), .op(n8244) );
  nand2_1 U9608 ( .ip1(n8244), .ip2(n5261), .op(n8245) );
  xnor2_1 U9609 ( .ip1(n5270), .ip2(n8245), .op(n8246) );
  inv_1 U9610 ( .ip(n8246), .op(n8254) );
  nor2_1 U9611 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[7]), .ip2(n8254), .op(n8251) );
  nand2_1 U9612 ( .ip1(n5261), .ip2(n8247), .op(n8248) );
  xnor2_1 U9613 ( .ip1(n5459), .ip2(n8248), .op(n8252) );
  inv_1 U9614 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[6]), .op(n8253)
         );
  nor3_1 U9615 ( .ip1(n8253), .ip2(n8252), .ip3(n8251), .op(n8255) );
  inv_1 U9616 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[8]), .op(n8274)
         );
  nand2_1 U9617 ( .ip1(n5267), .ip2(n8260), .op(n8259) );
  xnor2_1 U9618 ( .ip1(n8262), .ip2(n8259), .op(n8278) );
  inv_1 U9619 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[10]), .op(n8279)
         );
  nand2_1 U9620 ( .ip1(n8278), .ip2(n8279), .op(n8267) );
  inv_1 U9621 ( .ip(n8260), .op(n8261) );
  nor2_1 U9622 ( .ip1(n8262), .ip2(n8261), .op(n8263) );
  nand2_1 U9623 ( .ip1(n5267), .ip2(n8263), .op(n8264) );
  inv_1 U9624 ( .ip(n8266), .op(n8282) );
  nand2_1 U9625 ( .ip1(n8267), .ip2(n5546), .op(n8275) );
  ab_or_c_or_d U9626 ( .ip1(n8271), .ip2(n8270), .ip3(n8269), .ip4(n8268), 
        .op(n8283) );
  nor2_1 U9627 ( .ip1(n8275), .ip2(n8276), .op(n8281) );
  nor3_1 U9628 ( .ip1(n8279), .ip2(n8278), .ip3(n8277), .op(n8280) );
  not_ab_or_c_or_d U9629 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[11]), 
        .ip2(n8282), .ip3(n8281), .ip4(n8280), .op(n8284) );
  nor2_1 U9630 ( .ip1(n8284), .ip2(n8283), .op(n8285) );
  nand2_1 U9631 ( .ip1(n8304), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[0]), .op(n8306) );
  nor2_1 U9632 ( .ip1(n8289), .ip2(n8306), .op(n8308) );
  nand2_1 U9633 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[7]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[8]), .op(n8291) );
  nand2_1 U9634 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[10]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[11]), .op(n8292) );
  nor2_1 U9635 ( .ip1(n8319), .ip2(n8292), .op(n8321) );
  nand2_1 U9636 ( .ip1(n8321), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[12]), .op(n8323) );
  inv_1 U9637 ( .ip(n8323), .op(n8293) );
  nand2_1 U9638 ( .ip1(n8293), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[13]), .op(n8295) );
  nand2_1 U9639 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[13]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[14]), .op(n8294) );
  nor2_1 U9640 ( .ip1(n8294), .ip2(n8323), .op(n8325) );
  not_ab_or_c_or_d U9641 ( .ip1(n8196), .ip2(n8295), .ip3(n9335), .ip4(n8325), 
        .op(n4144) );
  inv_1 U9642 ( .ip(n8319), .op(n8296) );
  nand2_1 U9643 ( .ip1(n8296), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[10]), .op(n8297) );
  not_ab_or_c_or_d U9644 ( .ip1(n5547), .ip2(n8297), .ip3(n9335), .ip4(n8321), 
        .op(n4147) );
  inv_1 U9645 ( .ip(n8314), .op(n8298) );
  nand2_1 U9646 ( .ip1(n8298), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[7]), .op(n8299) );
  not_ab_or_c_or_d U9647 ( .ip1(n8274), .ip2(n8299), .ip3(n8316), .ip4(n9335), 
        .op(n4150) );
  inv_1 U9648 ( .ip(n8310), .op(n8300) );
  nand2_1 U9649 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[4]), .ip2(
        n8300), .op(n8301) );
  not_ab_or_c_or_d U9650 ( .ip1(n5545), .ip2(n8301), .ip3(n8312), .ip4(n9335), 
        .op(n4153) );
  inv_1 U9651 ( .ip(n8306), .op(n8302) );
  nand2_1 U9652 ( .ip1(n8302), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[1]), .op(n8303) );
  not_ab_or_c_or_d U9653 ( .ip1(n8233), .ip2(n8303), .ip3(n8308), .ip4(n9335), 
        .op(n4156) );
  nor2_1 U9654 ( .ip1(n9335), .ip2(n8305), .op(n4158) );
  xor2_1 U9655 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[1]), .ip2(n8306), .op(n8307) );
  nor2_1 U9656 ( .ip1(n9335), .ip2(n8307), .op(n4157) );
  xor2_1 U9657 ( .ip1(n8224), .ip2(n8308), .op(n8309) );
  xor2_1 U9658 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[4]), .ip2(n8310), .op(n8311) );
  xor2_1 U9659 ( .ip1(n8253), .ip2(n8312), .op(n8313) );
  xor2_1 U9660 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[7]), .ip2(n8314), .op(n8315) );
  inv_1 U9661 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[9]), .op(n8317)
         );
  nor2_1 U9662 ( .ip1(n9335), .ip2(n8318), .op(n4149) );
  nor2_1 U9663 ( .ip1(n9335), .ip2(n8320), .op(n4148) );
  nor2_1 U9664 ( .ip1(n9335), .ip2(n8322), .op(n4146) );
  xor2_1 U9665 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[13]), .ip2(
        n8323), .op(n8324) );
  nor2_1 U9666 ( .ip1(n9335), .ip2(n8324), .op(n4145) );
  xnor2_1 U9667 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_high_cntr[15]), .ip2(
        n8325), .op(n8326) );
  nor2_1 U9668 ( .ip1(n9335), .ip2(n8326), .op(n4143) );
  nand2_1 U9669 ( .ip1(n8328), .ip2(n8327), .op(n8329) );
  nand2_1 U9670 ( .ip1(n8333), .ip2(n8332), .op(i_i2c_U_DW_apb_i2c_mstfsm_N421) );
  inv_1 U9671 ( .ip(n11857), .op(n8335) );
  nor2_1 U9672 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_stop_scl_lcnt_en), .ip2(
        n9473), .op(n8334) );
  nor2_1 U9673 ( .ip1(n8335), .ip2(n8334), .op(n5041) );
  nor3_1 U9674 ( .ip1(i_i2c_scl_s_setup_en), .ip2(i_i2c_scl_s_setup_cmplt), 
        .ip3(n6352), .op(n8338) );
  and2_1 U9675 ( .ip1(i_i2c_re_start_en), .ip2(i_i2c_scl_lcnt_cmplt), .op(
        n8336) );
  and2_1 U9676 ( .ip1(n9473), .ip2(n8336), .op(n8339) );
  nand2_1 U9677 ( .ip1(n8339), .ip2(n8337), .op(n8526) );
  nor2_1 U9678 ( .ip1(n8338), .ip2(n8526), .op(n8344) );
  inv_1 U9679 ( .ip(i_i2c_scl_s_setup_en), .op(n8388) );
  inv_1 U9680 ( .ip(i_i2c_re_start_en), .op(n8994) );
  nand2_1 U9681 ( .ip1(n8339), .ip2(i_i2c_scl_s_setup_cmplt), .op(n8340) );
  nand2_1 U9682 ( .ip1(n8526), .ip2(n8340), .op(n8992) );
  nor2_1 U9683 ( .ip1(n8994), .ip2(n8992), .op(n9319) );
  nor2_1 U9684 ( .ip1(i_i2c_scl_lcnt_cmplt), .ip2(i_i2c_scl_s_hld_cmplt), .op(
        n8342) );
  inv_1 U9685 ( .ip(i_i2c_scl_s_setup_cmplt), .op(n8341) );
  nand2_1 U9686 ( .ip1(n8342), .ip2(n8341), .op(n9317) );
  nand2_1 U9687 ( .ip1(n9319), .ip2(n9317), .op(n8524) );
  nor2_1 U9688 ( .ip1(n8388), .ip2(n8524), .op(n8343) );
  or2_1 U9689 ( .ip1(n8344), .ip2(n8343), .op(n5191) );
  xor2_1 U9690 ( .ip1(n8345), .ip2(n8385), .op(n8346) );
  nor2_1 U9691 ( .ip1(n8388), .ip2(n8346), .op(n5146) );
  nand2_1 U9692 ( .ip1(n8385), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[0]), .op(n8348) );
  xor2_1 U9693 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[1]), .ip2(
        n8348), .op(n8347) );
  nor2_1 U9694 ( .ip1(n8388), .ip2(n8347), .op(n5145) );
  inv_1 U9695 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[2]), .op(n8353) );
  inv_1 U9696 ( .ip(n8348), .op(n8349) );
  nand2_1 U9697 ( .ip1(n8349), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[1]), .op(n8352) );
  nand2_1 U9698 ( .ip1(n8385), .ip2(n8350), .op(n8354) );
  inv_1 U9699 ( .ip(n8354), .op(n8351) );
  not_ab_or_c_or_d U9700 ( .ip1(n8353), .ip2(n8352), .ip3(n8351), .ip4(n8388), 
        .op(n5144) );
  xor2_1 U9701 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[3]), .ip2(
        n8354), .op(n8355) );
  nor2_1 U9702 ( .ip1(n8388), .ip2(n8355), .op(n5143) );
  nand2_1 U9703 ( .ip1(n8385), .ip2(n7152), .op(n8357) );
  xor2_1 U9704 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[4]), .ip2(
        n8357), .op(n8356) );
  nor2_1 U9705 ( .ip1(n8388), .ip2(n8356), .op(n5142) );
  inv_1 U9706 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[5]), .op(n8360) );
  inv_1 U9707 ( .ip(n8357), .op(n8358) );
  nand2_1 U9708 ( .ip1(n8358), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[4]), .op(n8359) );
  not_ab_or_c_or_d U9709 ( .ip1(n8360), .ip2(n8359), .ip3(n5594), .ip4(n8388), 
        .op(n5141) );
  inv_1 U9710 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[6]), .op(n8361) );
  xor2_1 U9711 ( .ip1(n8361), .ip2(n5594), .op(n8362) );
  xor2_1 U9712 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[7]), .ip2(
        n8364), .op(n8363) );
  nor2_1 U9713 ( .ip1(n8388), .ip2(n8363), .op(n5139) );
  inv_1 U9714 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[8]), .op(n8367) );
  inv_1 U9715 ( .ip(n8364), .op(n8365) );
  nand2_1 U9716 ( .ip1(n8365), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[7]), .op(n8366) );
  not_ab_or_c_or_d U9717 ( .ip1(n8367), .ip2(n8366), .ip3(n8368), .ip4(n8388), 
        .op(n5138) );
  inv_1 U9718 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[9]), .op(n8369) );
  xor2_1 U9719 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[10]), .ip2(
        n8372), .op(n8371) );
  nor2_1 U9720 ( .ip1(n8388), .ip2(n8371), .op(n5136) );
  inv_1 U9721 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[11]), .op(
        n8375) );
  inv_1 U9722 ( .ip(n8372), .op(n8373) );
  nand2_1 U9723 ( .ip1(n8373), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[10]), .op(n8374) );
  not_ab_or_c_or_d U9724 ( .ip1(n8375), .ip2(n8374), .ip3(n8376), .ip4(n8388), 
        .op(n5135) );
  inv_1 U9725 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[12]), .op(
        n8377) );
  xor2_1 U9726 ( .ip1(n8377), .ip2(n8376), .op(n8378) );
  xor2_1 U9727 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[13]), .ip2(
        n8380), .op(n8379) );
  nor2_1 U9728 ( .ip1(n8388), .ip2(n8379), .op(n5133) );
  inv_1 U9729 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[14]), .op(
        n8384) );
  inv_1 U9730 ( .ip(n8380), .op(n8381) );
  nand2_1 U9731 ( .ip1(n8381), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_setup_cntr[13]), .op(n8383) );
  not_ab_or_c_or_d U9732 ( .ip1(n8384), .ip2(n8383), .ip3(n8382), .ip4(n8388), 
        .op(n5132) );
  inv_1 U9733 ( .ip(n8385), .op(n8386) );
  nor2_1 U9734 ( .ip1(i_i2c_scl_s_setup_cmplt), .ip2(n8386), .op(n8387) );
  nor2_1 U9735 ( .ip1(n8388), .ip2(n8387), .op(n5190) );
  inv_1 U9736 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl_lcnt_en), .op(
        n8389) );
  nand2_1 U9737 ( .ip1(n9317), .ip2(n8389), .op(n8390) );
  nand2_1 U9738 ( .ip1(n9319), .ip2(n8390), .op(n8391) );
  nand2_1 U9739 ( .ip1(n8391), .ip2(n8526), .op(n4955) );
  inv_1 U9740 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[14]), .op(n8477)
         );
  nand2_1 U9741 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[10]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[11]), .op(n8473) );
  nand2_1 U9742 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[7]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[8]), .op(n8472) );
  nand2_1 U9743 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[4]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[5]), .op(n8471) );
  nand2_1 U9744 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[1]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[2]), .op(n8470) );
  nand2_1 U9745 ( .ip1(n5277), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[15]), .op(n8395) );
  nor2_1 U9746 ( .ip1(n5277), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[15]), .op(n8396) );
  nand2_1 U9747 ( .ip1(n5276), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[14]), .op(n8393) );
  or2_1 U9748 ( .ip1(n8396), .ip2(n8393), .op(n8394) );
  nand2_1 U9749 ( .ip1(n8395), .ip2(n8394), .op(n8403) );
  nor2_1 U9750 ( .ip1(n5276), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[14]), .op(n8397) );
  nor2_1 U9751 ( .ip1(n8397), .ip2(n8396), .op(n8406) );
  nand2_1 U9752 ( .ip1(n5268), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[13]), .op(n8400) );
  nand2_1 U9753 ( .ip1(n5275), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[12]), .op(n8398) );
  or2_1 U9754 ( .ip1(n8404), .ip2(n8398), .op(n8399) );
  nand2_1 U9755 ( .ip1(n8400), .ip2(n8399), .op(n8401) );
  and2_1 U9756 ( .ip1(n8406), .ip2(n8401), .op(n8402) );
  nor2_1 U9757 ( .ip1(n8403), .ip2(n8402), .op(n8422) );
  nor2_1 U9758 ( .ip1(n5275), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[12]), .op(n8405) );
  nor2_1 U9759 ( .ip1(n8405), .ip2(n8404), .op(n8407) );
  nand2_1 U9760 ( .ip1(n8407), .ip2(n8406), .op(n8427) );
  nand2_1 U9761 ( .ip1(n5269), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[11]), .op(n8411) );
  nor2_1 U9762 ( .ip1(n5269), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[11]), .op(n8412) );
  nand2_1 U9763 ( .ip1(n8408), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[10]), .op(n8409) );
  or2_1 U9764 ( .ip1(n8412), .ip2(n8409), .op(n8410) );
  nand2_1 U9765 ( .ip1(n8411), .ip2(n8410), .op(n8419) );
  nor2_1 U9766 ( .ip1(n8408), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[10]), .op(n8413) );
  nor2_1 U9767 ( .ip1(n8413), .ip2(n8412), .op(n8425) );
  nand2_1 U9768 ( .ip1(n8858), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[9]), .op(n8416) );
  nand2_1 U9769 ( .ip1(n5259), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[8]), .op(n8414) );
  or2_1 U9770 ( .ip1(n8423), .ip2(n8414), .op(n8415) );
  nand2_1 U9771 ( .ip1(n8416), .ip2(n8415), .op(n8417) );
  and2_1 U9772 ( .ip1(n8425), .ip2(n8417), .op(n8418) );
  nor2_1 U9773 ( .ip1(n8419), .ip2(n8418), .op(n8420) );
  or2_1 U9774 ( .ip1(n8427), .ip2(n8420), .op(n8421) );
  nand2_1 U9775 ( .ip1(n8422), .ip2(n8421), .op(n8469) );
  nor2_1 U9776 ( .ip1(n5259), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[8]), 
        .op(n8424) );
  nor2_1 U9777 ( .ip1(n8424), .ip2(n8423), .op(n8426) );
  nand2_1 U9778 ( .ip1(n8426), .ip2(n8425), .op(n8428) );
  nor2_1 U9779 ( .ip1(n8428), .ip2(n8427), .op(n8467) );
  nand2_1 U9780 ( .ip1(n5266), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[7]), .op(n8432) );
  nor2_1 U9781 ( .ip1(n5266), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[7]), 
        .op(n8433) );
  nand2_1 U9782 ( .ip1(n5278), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[6]), .op(n8430) );
  or2_1 U9783 ( .ip1(n8433), .ip2(n8430), .op(n8431) );
  nand2_1 U9784 ( .ip1(n8432), .ip2(n8431), .op(n8441) );
  nor2_1 U9785 ( .ip1(n5278), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[6]), 
        .op(n8434) );
  nor2_1 U9786 ( .ip1(n8434), .ip2(n8433), .op(n8460) );
  nand2_1 U9787 ( .ip1(n8879), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[5]), .op(n8438) );
  nor2_1 U9788 ( .ip1(n8879), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[5]), 
        .op(n8458) );
  nand2_1 U9789 ( .ip1(n8457), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[4]), .op(n8436) );
  or2_1 U9790 ( .ip1(n8458), .ip2(n8436), .op(n8437) );
  nand2_1 U9791 ( .ip1(n8438), .ip2(n8437), .op(n8439) );
  and2_1 U9792 ( .ip1(n8460), .ip2(n8439), .op(n8440) );
  nor2_1 U9793 ( .ip1(n8441), .ip2(n8440), .op(n8465) );
  nand2_1 U9794 ( .ip1(n8442), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[3]), .op(n8446) );
  nor2_1 U9795 ( .ip1(n8442), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[3]), 
        .op(n8451) );
  nand2_1 U9796 ( .ip1(n5280), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[2]), .op(n8444) );
  or2_1 U9797 ( .ip1(n8451), .ip2(n8444), .op(n8445) );
  nand2_1 U9798 ( .ip1(n8446), .ip2(n8445), .op(n8456) );
  nand2_1 U9799 ( .ip1(n5245), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[1]), .op(n8450) );
  nor2_1 U9800 ( .ip1(n7121), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[0]), 
        .op(n8448) );
  nor2_1 U9801 ( .ip1(n5245), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[1]), 
        .op(n8447) );
  or2_1 U9802 ( .ip1(n8448), .ip2(n8447), .op(n8449) );
  nand2_1 U9803 ( .ip1(n8450), .ip2(n8449), .op(n8454) );
  nor2_1 U9804 ( .ip1(n5280), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[2]), 
        .op(n8452) );
  nor2_1 U9805 ( .ip1(n8452), .ip2(n8451), .op(n8453) );
  and2_1 U9806 ( .ip1(n8454), .ip2(n8453), .op(n8455) );
  nor2_1 U9807 ( .ip1(n8456), .ip2(n8455), .op(n8463) );
  nor2_1 U9808 ( .ip1(n8457), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[4]), 
        .op(n8459) );
  nor2_1 U9809 ( .ip1(n8459), .ip2(n8458), .op(n8461) );
  nand2_1 U9810 ( .ip1(n8461), .ip2(n8460), .op(n8462) );
  or2_1 U9811 ( .ip1(n8463), .ip2(n8462), .op(n8464) );
  nand2_1 U9812 ( .ip1(n8465), .ip2(n8464), .op(n8466) );
  and2_1 U9813 ( .ip1(n8467), .ip2(n8466), .op(n8468) );
  nand2_1 U9814 ( .ip1(n8490), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[0]), .op(n8492) );
  nor2_1 U9815 ( .ip1(n8470), .ip2(n8492), .op(n8494) );
  nand2_1 U9816 ( .ip1(n8494), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[3]), .op(n8497) );
  nor2_1 U9817 ( .ip1(n8471), .ip2(n8497), .op(n8499) );
  nand2_1 U9818 ( .ip1(n8499), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[6]), .op(n8502) );
  nor2_1 U9819 ( .ip1(n8472), .ip2(n8502), .op(n8504) );
  nand2_1 U9820 ( .ip1(n8504), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[9]), .op(n8507) );
  nor2_1 U9821 ( .ip1(n8473), .ip2(n8507), .op(n8509) );
  and2_1 U9822 ( .ip1(n8509), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[12]), .op(n8512) );
  nand2_1 U9823 ( .ip1(n8512), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[13]), .op(n8476) );
  nor4_1 U9824 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_data_scl_lcnt_en), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl_lcnt_en), .ip3(
        i_i2c_rx_scl_lcnt_en), .ip4(
        i_i2c_U_DW_apb_i2c_tx_shift_stop_scl_lcnt_en), .op(n8474) );
  or2_1 U9825 ( .ip1(n8474), .ip2(n5591), .op(n8518) );
  nand3_1 U9826 ( .ip1(n8512), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[13]), .ip3(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[14]), .op(n8516) );
  inv_1 U9827 ( .ip(n8516), .op(n8475) );
  not_ab_or_c_or_d U9828 ( .ip1(n8477), .ip2(n8476), .ip3(n8518), .ip4(n8475), 
        .op(n5164) );
  inv_1 U9829 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[11]), .op(n8480)
         );
  inv_1 U9830 ( .ip(n8507), .op(n8478) );
  nand2_1 U9831 ( .ip1(n8478), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[10]), .op(n8479) );
  not_ab_or_c_or_d U9832 ( .ip1(n8480), .ip2(n8479), .ip3(n8509), .ip4(n8518), 
        .op(n5167) );
  inv_1 U9833 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[8]), .op(n8483) );
  inv_1 U9834 ( .ip(n8502), .op(n8481) );
  nand2_1 U9835 ( .ip1(n8481), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[7]), .op(n8482) );
  not_ab_or_c_or_d U9836 ( .ip1(n8483), .ip2(n8482), .ip3(n8504), .ip4(n8518), 
        .op(n5170) );
  inv_1 U9837 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[5]), .op(n8486) );
  inv_1 U9838 ( .ip(n8497), .op(n8484) );
  nand2_1 U9839 ( .ip1(n8484), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[4]), .op(n8485) );
  not_ab_or_c_or_d U9840 ( .ip1(n8486), .ip2(n8485), .ip3(n8499), .ip4(n8518), 
        .op(n5173) );
  inv_1 U9841 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[2]), .op(n8489) );
  inv_1 U9842 ( .ip(n8492), .op(n8487) );
  nand2_1 U9843 ( .ip1(n8487), .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[1]), .op(n8488) );
  not_ab_or_c_or_d U9844 ( .ip1(n8489), .ip2(n8488), .ip3(n8494), .ip4(n8518), 
        .op(n5176) );
  inv_1 U9845 ( .ip(n8490), .op(n8519) );
  nor2_1 U9846 ( .ip1(n8518), .ip2(n8491), .op(n5178) );
  xor2_1 U9847 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[1]), .ip2(n8492), 
        .op(n8493) );
  nor2_1 U9848 ( .ip1(n8518), .ip2(n8493), .op(n5177) );
  inv_1 U9849 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[3]), .op(n8495) );
  nor2_1 U9850 ( .ip1(n8518), .ip2(n8496), .op(n5175) );
  xor2_1 U9851 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[4]), .ip2(n8497), 
        .op(n8498) );
  nor2_1 U9852 ( .ip1(n8518), .ip2(n8498), .op(n5174) );
  inv_1 U9853 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[6]), .op(n8500) );
  nor2_1 U9854 ( .ip1(n8518), .ip2(n8501), .op(n5172) );
  xor2_1 U9855 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[7]), .ip2(n8502), 
        .op(n8503) );
  nor2_1 U9856 ( .ip1(n8518), .ip2(n8503), .op(n5171) );
  inv_1 U9857 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[9]), .op(n8505) );
  xor2_1 U9858 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[10]), .ip2(n8507), .op(n8508) );
  nor2_1 U9859 ( .ip1(n8518), .ip2(n8508), .op(n5168) );
  inv_1 U9860 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[12]), .op(n8510)
         );
  inv_1 U9861 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[13]), .op(n8513)
         );
  xnor2_1 U9862 ( .ip1(n8513), .ip2(n8512), .op(n8514) );
  inv_1 U9863 ( .ip(n8514), .op(n8515) );
  nor2_1 U9864 ( .ip1(n8518), .ip2(n8515), .op(n5165) );
  xor2_1 U9865 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_low_cntr[15]), .ip2(n8516), .op(n8517) );
  nor2_1 U9866 ( .ip1(n8518), .ip2(n8517), .op(n5163) );
  inv_1 U9867 ( .ip(n8518), .op(n8522) );
  inv_1 U9868 ( .ip(n8519), .op(n8520) );
  nand2_1 U9869 ( .ip1(n11040), .ip2(n8520), .op(n8521) );
  inv_1 U9870 ( .ip(n8524), .op(n8525) );
  nand2_1 U9871 ( .ip1(n8525), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_re_scl_s_hld_en), .op(n8529) );
  inv_1 U9872 ( .ip(n8526), .op(n8527) );
  nand2_1 U9873 ( .ip1(n8527), .ip2(i_i2c_scl_s_setup_cmplt), .op(n8528) );
  nand2_1 U9874 ( .ip1(n8529), .ip2(n8528), .op(n5189) );
  nor2_1 U9875 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_re_scl_s_hld_en), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_st_scl_s_hld_en), .op(n9331) );
  inv_1 U9876 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[0]), .op(n8684)
         );
  nand2_1 U9877 ( .ip1(n5277), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[15]), .op(n8533) );
  nor2_1 U9878 ( .ip1(n5277), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[15]), .op(n8534) );
  nand2_1 U9879 ( .ip1(n5276), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[14]), .op(n8531) );
  or2_1 U9880 ( .ip1(n8534), .ip2(n8531), .op(n8532) );
  nand2_1 U9881 ( .ip1(n8533), .ip2(n8532), .op(n8543) );
  nor2_1 U9882 ( .ip1(n5276), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[14]), .op(n8535) );
  nor2_1 U9883 ( .ip1(n8535), .ip2(n8534), .op(n8546) );
  nand2_1 U9884 ( .ip1(n5268), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[13]), .op(n8540) );
  nand2_1 U9885 ( .ip1(n5275), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[12]), .op(n8538) );
  or2_1 U9886 ( .ip1(n8544), .ip2(n8538), .op(n8539) );
  nand2_1 U9887 ( .ip1(n8540), .ip2(n8539), .op(n8541) );
  and2_1 U9888 ( .ip1(n8546), .ip2(n8541), .op(n8542) );
  nor2_1 U9889 ( .ip1(n8543), .ip2(n8542), .op(n8564) );
  nor2_1 U9890 ( .ip1(n5275), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[12]), .op(n8545) );
  nor2_1 U9891 ( .ip1(n8545), .ip2(n8544), .op(n8547) );
  nand2_1 U9892 ( .ip1(n8547), .ip2(n8546), .op(n8569) );
  nand2_1 U9893 ( .ip1(n5269), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[11]), .op(n8553) );
  xor2_1 U9894 ( .ip1(n8550), .ip2(n8549), .op(n8855) );
  nand2_1 U9895 ( .ip1(n8855), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[10]), .op(n8551) );
  or2_1 U9896 ( .ip1(n8554), .ip2(n8551), .op(n8552) );
  nand2_1 U9897 ( .ip1(n8553), .ip2(n8552), .op(n8561) );
  nor2_1 U9898 ( .ip1(n8855), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[10]), .op(n8555) );
  nor2_1 U9899 ( .ip1(n8555), .ip2(n8554), .op(n8567) );
  nand2_1 U9900 ( .ip1(n8858), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[9]), .op(n8558) );
  nor2_1 U9901 ( .ip1(n8858), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[9]), .op(n8566) );
  nand2_1 U9902 ( .ip1(n5259), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[8]), .op(n8556) );
  or2_1 U9903 ( .ip1(n8566), .ip2(n8556), .op(n8557) );
  nand2_1 U9904 ( .ip1(n8558), .ip2(n8557), .op(n8559) );
  and2_1 U9905 ( .ip1(n8567), .ip2(n8559), .op(n8560) );
  nor2_1 U9906 ( .ip1(n8561), .ip2(n8560), .op(n8562) );
  or2_1 U9907 ( .ip1(n8569), .ip2(n8562), .op(n8563) );
  nand2_1 U9908 ( .ip1(n8564), .ip2(n8563), .op(n8607) );
  nor2_1 U9909 ( .ip1(n5259), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[8]), .op(n8565) );
  nor2_1 U9910 ( .ip1(n8566), .ip2(n8565), .op(n8568) );
  nand2_1 U9911 ( .ip1(n8568), .ip2(n8567), .op(n8570) );
  nor2_1 U9912 ( .ip1(n8570), .ip2(n8569), .op(n8605) );
  nand2_1 U9913 ( .ip1(n5266), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[7]), .op(n8574) );
  nand2_1 U9914 ( .ip1(n5278), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[6]), .op(n8572) );
  or2_1 U9915 ( .ip1(n8575), .ip2(n8572), .op(n8573) );
  nand2_1 U9916 ( .ip1(n8574), .ip2(n8573), .op(n8582) );
  nor2_1 U9917 ( .ip1(n5278), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[6]), .op(n8576) );
  nor2_1 U9918 ( .ip1(n8576), .ip2(n8575), .op(n8598) );
  nand2_1 U9919 ( .ip1(n8879), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[5]), .op(n8579) );
  nor2_1 U9920 ( .ip1(n8879), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[5]), .op(n8596) );
  nand2_1 U9921 ( .ip1(n8457), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[4]), .op(n8577) );
  or2_1 U9922 ( .ip1(n8596), .ip2(n8577), .op(n8578) );
  nand2_1 U9923 ( .ip1(n8579), .ip2(n8578), .op(n8580) );
  and2_1 U9924 ( .ip1(n8598), .ip2(n8580), .op(n8581) );
  nor2_1 U9925 ( .ip1(n8582), .ip2(n8581), .op(n8603) );
  nand2_1 U9926 ( .ip1(n8442), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[3]), .op(n8585) );
  nor2_1 U9927 ( .ip1(n8442), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[3]), .op(n8590) );
  nand2_1 U9928 ( .ip1(n5280), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[2]), .op(n8583) );
  or2_1 U9929 ( .ip1(n8590), .ip2(n8583), .op(n8584) );
  nand2_1 U9930 ( .ip1(n8585), .ip2(n8584), .op(n8595) );
  nand2_1 U9931 ( .ip1(n5245), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[1]), .op(n8589) );
  nor2_1 U9932 ( .ip1(n5245), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[1]), .op(n8587) );
  or2_1 U9933 ( .ip1(n8586), .ip2(n8587), .op(n8588) );
  nand2_1 U9934 ( .ip1(n8589), .ip2(n8588), .op(n8593) );
  nor2_1 U9935 ( .ip1(n5280), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[2]), .op(n8591) );
  nor2_1 U9936 ( .ip1(n8591), .ip2(n8590), .op(n8592) );
  and2_1 U9937 ( .ip1(n8593), .ip2(n8592), .op(n8594) );
  nor2_1 U9938 ( .ip1(n8595), .ip2(n8594), .op(n8601) );
  nor2_1 U9939 ( .ip1(n8457), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[4]), .op(n8597) );
  nor2_1 U9940 ( .ip1(n8597), .ip2(n8596), .op(n8599) );
  nand2_1 U9941 ( .ip1(n8599), .ip2(n8598), .op(n8600) );
  or2_1 U9942 ( .ip1(n8601), .ip2(n8600), .op(n8602) );
  nand2_1 U9943 ( .ip1(n8603), .ip2(n8602), .op(n8604) );
  and2_1 U9944 ( .ip1(n8605), .ip2(n8604), .op(n8606) );
  nor2_1 U9945 ( .ip1(n8607), .ip2(n8606), .op(n8608) );
  nand2_1 U9946 ( .ip1(n8608), .ip2(n8911), .op(n8683) );
  nand2_1 U9947 ( .ip1(n8772), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[15]), .op(n8611) );
  nand2_1 U9948 ( .ip1(n8773), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[14]), .op(n8609) );
  or2_1 U9949 ( .ip1(n8612), .ip2(n8609), .op(n8610) );
  nand2_1 U9950 ( .ip1(n8611), .ip2(n8610), .op(n8619) );
  nand2_1 U9951 ( .ip1(n8778), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[13]), .op(n8616) );
  nand2_1 U9952 ( .ip1(n8620), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[12]), .op(n8614) );
  or2_1 U9953 ( .ip1(n8621), .ip2(n8614), .op(n8615) );
  nand2_1 U9954 ( .ip1(n8616), .ip2(n8615), .op(n8617) );
  and2_1 U9955 ( .ip1(n8623), .ip2(n8617), .op(n8618) );
  nor2_1 U9956 ( .ip1(n8619), .ip2(n8618), .op(n8640) );
  nor2_1 U9957 ( .ip1(n8620), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[12]), .op(n8622) );
  nor2_1 U9958 ( .ip1(n8622), .ip2(n8621), .op(n8624) );
  nand2_1 U9959 ( .ip1(n8624), .ip2(n8623), .op(n8645) );
  inv_1 U9960 ( .ip(n8645), .op(n8638) );
  inv_1 U9961 ( .ip(n8757), .op(n8626) );
  nor2_1 U9962 ( .ip1(n8626), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[11]), .op(n8629) );
  nand2_1 U9963 ( .ip1(n8761), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[10]), .op(n8625) );
  nor2_1 U9964 ( .ip1(n8629), .ip2(n8625), .op(n8628) );
  nor2_1 U9965 ( .ip1(n8628), .ip2(n8627), .op(n8636) );
  nor2_1 U9966 ( .ip1(n8630), .ip2(n8629), .op(n8643) );
  nor2_1 U9967 ( .ip1(n5265), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[9]), .op(n8641) );
  nand2_1 U9968 ( .ip1(n5264), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[8]), .op(n8631) );
  or2_1 U9969 ( .ip1(n8641), .ip2(n8631), .op(n8633) );
  nand2_1 U9970 ( .ip1(n5265), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[9]), .op(n8632) );
  nand2_1 U9971 ( .ip1(n8633), .ip2(n8632), .op(n8634) );
  nand2_1 U9972 ( .ip1(n8643), .ip2(n8634), .op(n8635) );
  nand2_1 U9973 ( .ip1(n8636), .ip2(n8635), .op(n8637) );
  nand2_1 U9974 ( .ip1(n8638), .ip2(n8637), .op(n8639) );
  nand2_1 U9975 ( .ip1(n8640), .ip2(n8639), .op(n8681) );
  nor2_1 U9976 ( .ip1(n5264), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[8]), .op(n8642) );
  nor2_1 U9977 ( .ip1(n8642), .ip2(n8641), .op(n8644) );
  nand2_1 U9978 ( .ip1(n8644), .ip2(n8643), .op(n8646) );
  nor2_1 U9979 ( .ip1(n8646), .ip2(n8645), .op(n8680) );
  nand2_1 U9980 ( .ip1(n5597), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[7]), .op(n8649) );
  nand2_1 U9981 ( .ip1(n5598), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[6]), .op(n8647) );
  or2_1 U9982 ( .ip1(n8650), .ip2(n8647), .op(n8648) );
  nand2_1 U9983 ( .ip1(n8649), .ip2(n8648), .op(n8657) );
  nor2_1 U9984 ( .ip1(n5598), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[6]), .op(n8651) );
  nand2_1 U9985 ( .ip1(n8800), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[5]), .op(n8654) );
  nand2_1 U9986 ( .ip1(n8822), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[4]), .op(n8652) );
  or2_1 U9987 ( .ip1(n8671), .ip2(n8652), .op(n8653) );
  nand2_1 U9988 ( .ip1(n8654), .ip2(n8653), .op(n8655) );
  and2_1 U9989 ( .ip1(n8673), .ip2(n8655), .op(n8656) );
  nor2_1 U9990 ( .ip1(n8657), .ip2(n8656), .op(n8678) );
  nand2_1 U9991 ( .ip1(n5274), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[3]), .op(n8660) );
  nor2_1 U9992 ( .ip1(n5274), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[3]), .op(n8665) );
  nand2_1 U9993 ( .ip1(n8807), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[2]), .op(n8658) );
  or2_1 U9994 ( .ip1(n8665), .ip2(n8658), .op(n8659) );
  nand2_1 U9995 ( .ip1(n8660), .ip2(n8659), .op(n8670) );
  nand2_1 U9996 ( .ip1(n8811), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[1]), .op(n8664) );
  nor2_1 U9997 ( .ip1(n8811), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[1]), .op(n8662) );
  or2_1 U9998 ( .ip1(n8661), .ip2(n8662), .op(n8663) );
  nand2_1 U9999 ( .ip1(n8664), .ip2(n8663), .op(n8668) );
  nor2_1 U10000 ( .ip1(n8807), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[2]), .op(n8666) );
  nor2_1 U10001 ( .ip1(n8666), .ip2(n8665), .op(n8667) );
  and2_1 U10002 ( .ip1(n8668), .ip2(n8667), .op(n8669) );
  nor2_1 U10003 ( .ip1(n8670), .ip2(n8669), .op(n8676) );
  nor2_1 U10004 ( .ip1(n8822), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[4]), .op(n8672) );
  nor2_1 U10005 ( .ip1(n8672), .ip2(n8671), .op(n8674) );
  nand2_1 U10006 ( .ip1(n8674), .ip2(n8673), .op(n8675) );
  or2_1 U10007 ( .ip1(n8676), .ip2(n8675), .op(n8677) );
  nand2_1 U10008 ( .ip1(n8678), .ip2(n8677), .op(n8679) );
  xor2_1 U10009 ( .ip1(n8684), .ip2(n8730), .op(n8685) );
  nor2_1 U10010 ( .ip1(n9331), .ip2(n8685), .op(n5162) );
  xor2_1 U10011 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[1]), .ip2(
        n8688), .op(n8686) );
  inv_1 U10012 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[2]), .op(n8691)
         );
  inv_1 U10013 ( .ip(n8688), .op(n8687) );
  nand2_1 U10014 ( .ip1(n8687), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[1]), .op(n8690) );
  nand2_1 U10015 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[1]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[2]), .op(n8689) );
  not_ab_or_c_or_d U10016 ( .ip1(n8691), .ip2(n8690), .ip3(n9331), .ip4(n8693), 
        .op(n5160) );
  inv_1 U10017 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[3]), .op(n8692)
         );
  nor2_1 U10018 ( .ip1(n9331), .ip2(n5262), .op(n5159) );
  xor2_1 U10019 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[4]), .ip2(
        n8696), .op(n8694) );
  nor2_1 U10020 ( .ip1(n9331), .ip2(n8694), .op(n5158) );
  inv_1 U10021 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[5]), .op(n8699)
         );
  inv_1 U10022 ( .ip(n8696), .op(n8695) );
  nand2_1 U10023 ( .ip1(n8695), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[4]), .op(n8698) );
  nand2_1 U10024 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[4]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[5]), .op(n8697) );
  not_ab_or_c_or_d U10025 ( .ip1(n8699), .ip2(n8698), .ip3(n9331), .ip4(n8702), 
        .op(n5157) );
  inv_1 U10026 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[6]), .op(n8700)
         );
  xor2_1 U10027 ( .ip1(n8700), .ip2(n8702), .op(n8701) );
  xor2_1 U10028 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[7]), .ip2(
        n8705), .op(n8703) );
  inv_1 U10029 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[8]), .op(n8708)
         );
  inv_1 U10030 ( .ip(n8705), .op(n8704) );
  nand2_1 U10031 ( .ip1(n8704), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[7]), .op(n8707) );
  nand2_1 U10032 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[7]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[8]), .op(n8706) );
  not_ab_or_c_or_d U10033 ( .ip1(n8708), .ip2(n8707), .ip3(n9331), .ip4(n8711), 
        .op(n5154) );
  inv_1 U10034 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[9]), .op(n8709)
         );
  xor2_1 U10035 ( .ip1(n8709), .ip2(n8711), .op(n8710) );
  nor2_1 U10036 ( .ip1(n9331), .ip2(n5538), .op(n5152) );
  inv_1 U10037 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[11]), .op(n8716) );
  inv_1 U10038 ( .ip(n8713), .op(n8712) );
  nand2_1 U10039 ( .ip1(n8712), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[10]), .op(n8715) );
  nand2_1 U10040 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[10]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[11]), .op(n8714) );
  nor2_1 U10041 ( .ip1(n8714), .ip2(n8713), .op(n8720) );
  not_ab_or_c_or_d U10042 ( .ip1(n8716), .ip2(n8715), .ip3(n9331), .ip4(n8720), 
        .op(n5151) );
  inv_1 U10043 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[12]), .op(n8717) );
  xnor2_1 U10044 ( .ip1(n8717), .ip2(n8720), .op(n8718) );
  inv_1 U10045 ( .ip(n8718), .op(n8719) );
  nor2_1 U10046 ( .ip1(n9331), .ip2(n8719), .op(n5150) );
  inv_1 U10047 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[13]), .op(n8721) );
  and2_1 U10048 ( .ip1(n8720), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[12]), .op(n8724) );
  xnor2_1 U10049 ( .ip1(n8721), .ip2(n8724), .op(n8722) );
  inv_1 U10050 ( .ip(n8722), .op(n8723) );
  nor2_1 U10051 ( .ip1(n9331), .ip2(n8723), .op(n5149) );
  inv_1 U10052 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[14]), .op(n8727) );
  nand2_1 U10053 ( .ip1(n8724), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[13]), .op(n8726) );
  nand3_1 U10054 ( .ip1(n8724), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[13]), .ip3(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[14]), .op(n8728) );
  inv_1 U10055 ( .ip(n8728), .op(n8725) );
  not_ab_or_c_or_d U10056 ( .ip1(n8727), .ip2(n8726), .ip3(n9331), .ip4(n8725), 
        .op(n5148) );
  xor2_1 U10057 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_s_hld_cntr[15]), .ip2(
        n8728), .op(n8729) );
  nor2_1 U10058 ( .ip1(n9331), .ip2(n8729), .op(n5147) );
  inv_1 U10059 ( .ip(n8730), .op(n8731) );
  nor2_1 U10060 ( .ip1(i_i2c_scl_s_hld_cmplt), .ip2(n8731), .op(n8732) );
  nor2_1 U10061 ( .ip1(n9331), .ip2(n8732), .op(n5188) );
  inv_1 U10062 ( .ip(i_i2c_tx_rd_addr[1]), .op(n8733) );
  nor3_1 U10063 ( .ip1(i_i2c_tx_rd_addr[2]), .ip2(i_i2c_tx_rd_addr[0]), .ip3(
        n8733), .op(n10178) );
  nand2_1 U10064 ( .ip1(n10178), .ip2(i_i2c_U_dff_tx_mem[53]), .op(n8743) );
  inv_1 U10065 ( .ip(i_i2c_tx_rd_addr[2]), .op(n8734) );
  nor3_1 U10066 ( .ip1(i_i2c_tx_rd_addr[0]), .ip2(i_i2c_tx_rd_addr[1]), .ip3(
        n8734), .op(n10180) );
  inv_1 U10067 ( .ip(i_i2c_tx_rd_addr[0]), .op(n11228) );
  nor3_1 U10068 ( .ip1(n8734), .ip2(n11228), .ip3(n8733), .op(n11214) );
  and2_1 U10069 ( .ip1(n11214), .ip2(i_i2c_U_dff_tx_mem[8]), .op(n8740) );
  nor3_1 U10070 ( .ip1(i_i2c_tx_rd_addr[1]), .ip2(n11228), .ip3(n8734), .op(
        n10179) );
  nand2_1 U10071 ( .ip1(n10179), .ip2(i_i2c_U_dff_tx_mem[26]), .op(n8738) );
  nor3_1 U10072 ( .ip1(i_i2c_tx_rd_addr[2]), .ip2(i_i2c_tx_rd_addr[1]), .ip3(
        n11228), .op(n10181) );
  nand2_1 U10073 ( .ip1(n10181), .ip2(i_i2c_U_dff_tx_mem[62]), .op(n8737) );
  nor3_1 U10074 ( .ip1(i_i2c_tx_rd_addr[2]), .ip2(i_i2c_tx_rd_addr[0]), .ip3(
        i_i2c_tx_rd_addr[1]), .op(n10182) );
  nand2_1 U10075 ( .ip1(n10182), .ip2(i_i2c_U_dff_tx_mem[71]), .op(n8736) );
  nor3_1 U10076 ( .ip1(i_i2c_tx_rd_addr[0]), .ip2(n8734), .ip3(n8733), .op(
        n10189) );
  nand2_1 U10077 ( .ip1(n10189), .ip2(i_i2c_U_dff_tx_mem[17]), .op(n8735) );
  nand4_1 U10078 ( .ip1(n8738), .ip2(n8737), .ip3(n8736), .ip4(n8735), .op(
        n8739) );
  not_ab_or_c_or_d U10079 ( .ip1(n10180), .ip2(i_i2c_U_dff_tx_mem[35]), .ip3(
        n8740), .ip4(n8739), .op(n8742) );
  nand2_1 U10080 ( .ip1(i_i2c_tx_rd_addr[0]), .ip2(i_i2c_tx_rd_addr[1]), .op(
        n11209) );
  nor2_1 U10081 ( .ip1(i_i2c_tx_rd_addr[2]), .ip2(n11209), .op(n10190) );
  nand2_1 U10082 ( .ip1(n10190), .ip2(i_i2c_U_dff_tx_mem[44]), .op(n8741) );
  nand3_1 U10083 ( .ip1(n8743), .ip2(n8742), .ip3(n8741), .op(n8744) );
  mux2_1 U10084 ( .ip1(i_i2c_tx_fifo_data_buf[8]), .ip2(n8744), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .op(n5214) );
  nand3_1 U10085 ( .ip1(n8745), .ip2(i_i2c_U_DW_apb_i2c_mstfsm_addr_1byte_sent), .ip3(i_i2c_U_DW_apb_i2c_mstfsm_N487), .op(n8747) );
  nand2_1 U10086 ( .ip1(n8747), .ip2(n8746), .op(n5200) );
  nand2_1 U10087 ( .ip1(n6352), .ip2(i_i2c_scl_lcnt_cmplt), .op(n8748) );
  inv_1 U10088 ( .ip(i_i2c_scl_p_setup_cmplt), .op(n9474) );
  nand2_1 U10089 ( .ip1(n8748), .ip2(n9474), .op(n8749) );
  nand2_1 U10090 ( .ip1(n9473), .ip2(n8749), .op(n8751) );
  nand2_1 U10091 ( .ip1(n9474), .ip2(n11040), .op(n9309) );
  nand2_1 U10092 ( .ip1(n9309), .ip2(i_i2c_scl_p_setup_en), .op(n8750) );
  nand2_1 U10093 ( .ip1(n8751), .ip2(n8750), .op(n8752) );
  and2_1 U10094 ( .ip1(n8752), .ip2(n11857), .op(n5061) );
  inv_1 U10095 ( .ip(i_i2c_scl_p_setup_en), .op(n8965) );
  inv_1 U10096 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[0]), .op(
        n8915) );
  nor2_1 U10097 ( .ip1(n8620), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[12]), .op(n8753) );
  nor2_1 U10098 ( .ip1(n8778), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[13]), .op(n8780) );
  nor2_1 U10099 ( .ip1(n8753), .ip2(n8780), .op(n8756) );
  nor2_1 U10100 ( .ip1(n8773), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[14]), .op(n8755) );
  nor2_1 U10101 ( .ip1(n8754), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[15]), .op(n8775) );
  nor2_1 U10102 ( .ip1(n8755), .ip2(n8775), .op(n8784) );
  nand2_1 U10103 ( .ip1(n8756), .ip2(n8784), .op(n8793) );
  nand2_1 U10104 ( .ip1(n5273), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[11]), .op(n8760) );
  nor2_1 U10105 ( .ip1(n5273), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[11]), .op(n8762) );
  nand2_1 U10106 ( .ip1(n8761), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[10]), .op(n8758) );
  or2_1 U10107 ( .ip1(n8762), .ip2(n8758), .op(n8759) );
  nand2_1 U10108 ( .ip1(n8760), .ip2(n8759), .op(n8770) );
  nor2_1 U10109 ( .ip1(n8761), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[10]), .op(n8763) );
  nor2_1 U10110 ( .ip1(n8763), .ip2(n8762), .op(n8791) );
  nand2_1 U10111 ( .ip1(n5265), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[9]), .op(n8767) );
  nor2_1 U10112 ( .ip1(n5265), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[9]), .op(n8789) );
  nand2_1 U10113 ( .ip1(n5264), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[8]), .op(n8765) );
  or2_1 U10114 ( .ip1(n8789), .ip2(n8765), .op(n8766) );
  nand2_1 U10115 ( .ip1(n8767), .ip2(n8766), .op(n8768) );
  and2_1 U10116 ( .ip1(n8791), .ip2(n8768), .op(n8769) );
  nor2_1 U10117 ( .ip1(n8770), .ip2(n8769), .op(n8771) );
  or2_1 U10118 ( .ip1(n8793), .ip2(n8771), .op(n8788) );
  nand2_1 U10119 ( .ip1(n8772), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[15]), .op(n8777) );
  nand2_1 U10120 ( .ip1(n8773), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[14]), .op(n8774) );
  or2_1 U10121 ( .ip1(n8775), .ip2(n8774), .op(n8776) );
  nand2_1 U10122 ( .ip1(n8777), .ip2(n8776), .op(n8786) );
  nand2_1 U10123 ( .ip1(n8778), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[13]), .op(n8782) );
  nand2_1 U10124 ( .ip1(n8620), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[12]), .op(n8779) );
  or2_1 U10125 ( .ip1(n8780), .ip2(n8779), .op(n8781) );
  nand2_1 U10126 ( .ip1(n8782), .ip2(n8781), .op(n8783) );
  and2_1 U10127 ( .ip1(n8784), .ip2(n8783), .op(n8785) );
  nor2_1 U10128 ( .ip1(n8786), .ip2(n8785), .op(n8787) );
  nand2_1 U10129 ( .ip1(n8788), .ip2(n8787), .op(n8834) );
  nor2_1 U10130 ( .ip1(n5264), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[8]), .op(n8790) );
  nor2_1 U10131 ( .ip1(n8790), .ip2(n8789), .op(n8792) );
  nand2_1 U10132 ( .ip1(n8792), .ip2(n8791), .op(n8794) );
  nor2_1 U10133 ( .ip1(n8794), .ip2(n8793), .op(n8832) );
  nand2_1 U10134 ( .ip1(n5597), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[7]), .op(n8797) );
  nor2_1 U10135 ( .ip1(n5597), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[7]), .op(n8798) );
  nand2_1 U10136 ( .ip1(n5598), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[6]), .op(n8795) );
  or2_1 U10137 ( .ip1(n8798), .ip2(n8795), .op(n8796) );
  nand2_1 U10138 ( .ip1(n8797), .ip2(n8796), .op(n8806) );
  nor2_1 U10139 ( .ip1(n5598), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[6]), .op(n8799) );
  nor2_1 U10140 ( .ip1(n8799), .ip2(n8798), .op(n8825) );
  nand2_1 U10141 ( .ip1(n8800), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[5]), .op(n8803) );
  nor2_1 U10142 ( .ip1(n8800), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[5]), .op(n8823) );
  nand2_1 U10143 ( .ip1(n8822), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[4]), .op(n8801) );
  or2_1 U10144 ( .ip1(n8823), .ip2(n8801), .op(n8802) );
  nand2_1 U10145 ( .ip1(n8803), .ip2(n8802), .op(n8804) );
  and2_1 U10146 ( .ip1(n8825), .ip2(n8804), .op(n8805) );
  nor2_1 U10147 ( .ip1(n8806), .ip2(n8805), .op(n8830) );
  nand2_1 U10148 ( .ip1(n5274), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[3]), .op(n8810) );
  nor2_1 U10149 ( .ip1(n5274), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[3]), .op(n8816) );
  nand2_1 U10150 ( .ip1(n8807), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[2]), .op(n8808) );
  or2_1 U10151 ( .ip1(n8816), .ip2(n8808), .op(n8809) );
  nand2_1 U10152 ( .ip1(n8810), .ip2(n8809), .op(n8821) );
  nand2_1 U10153 ( .ip1(n8811), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[1]), .op(n8815) );
  nor2_1 U10154 ( .ip1(n6994), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[0]), .op(n8813) );
  nor2_1 U10155 ( .ip1(n8811), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[1]), .op(n8812) );
  or2_1 U10156 ( .ip1(n8813), .ip2(n8812), .op(n8814) );
  nand2_1 U10157 ( .ip1(n8815), .ip2(n8814), .op(n8819) );
  nor2_1 U10158 ( .ip1(n8807), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[2]), .op(n8817) );
  nor2_1 U10159 ( .ip1(n8817), .ip2(n8816), .op(n8818) );
  and2_1 U10160 ( .ip1(n8819), .ip2(n8818), .op(n8820) );
  nor2_1 U10161 ( .ip1(n8821), .ip2(n8820), .op(n8828) );
  nor2_1 U10162 ( .ip1(n8822), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[4]), .op(n8824) );
  nor2_1 U10163 ( .ip1(n8824), .ip2(n8823), .op(n8826) );
  nand2_1 U10164 ( .ip1(n8826), .ip2(n8825), .op(n8827) );
  or2_1 U10165 ( .ip1(n8828), .ip2(n8827), .op(n8829) );
  nand2_1 U10166 ( .ip1(n8830), .ip2(n8829), .op(n8831) );
  and2_1 U10167 ( .ip1(n8832), .ip2(n8831), .op(n8833) );
  nor2_1 U10168 ( .ip1(n8834), .ip2(n8833), .op(n8836) );
  nand2_1 U10169 ( .ip1(n8836), .ip2(n8835), .op(n8914) );
  nand2_1 U10170 ( .ip1(n5277), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[15]), .op(n8839) );
  nor2_1 U10171 ( .ip1(n5277), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[15]), .op(n8840) );
  nand2_1 U10172 ( .ip1(n5276), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[14]), .op(n8837) );
  or2_1 U10173 ( .ip1(n8840), .ip2(n8837), .op(n8838) );
  nand2_1 U10174 ( .ip1(n8839), .ip2(n8838), .op(n8847) );
  nor2_1 U10175 ( .ip1(n5276), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[14]), .op(n8841) );
  nor2_1 U10176 ( .ip1(n8841), .ip2(n8840), .op(n8850) );
  nand2_1 U10177 ( .ip1(n5268), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[13]), .op(n8844) );
  nor2_1 U10178 ( .ip1(n5268), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[13]), .op(n8848) );
  nand2_1 U10179 ( .ip1(n5275), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[12]), .op(n8842) );
  or2_1 U10180 ( .ip1(n8848), .ip2(n8842), .op(n8843) );
  nand2_1 U10181 ( .ip1(n8844), .ip2(n8843), .op(n8845) );
  and2_1 U10182 ( .ip1(n8850), .ip2(n8845), .op(n8846) );
  nor2_1 U10183 ( .ip1(n8847), .ip2(n8846), .op(n8867) );
  nor2_1 U10184 ( .ip1(n5275), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[12]), .op(n8849) );
  nor2_1 U10185 ( .ip1(n8849), .ip2(n8848), .op(n8851) );
  nand2_1 U10186 ( .ip1(n8851), .ip2(n8850), .op(n8872) );
  nand2_1 U10187 ( .ip1(n5269), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[11]), .op(n8854) );
  nor2_1 U10188 ( .ip1(n5269), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[11]), .op(n8856) );
  nand2_1 U10189 ( .ip1(n8855), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[10]), .op(n8852) );
  or2_1 U10190 ( .ip1(n8856), .ip2(n8852), .op(n8853) );
  nand2_1 U10191 ( .ip1(n8854), .ip2(n8853), .op(n8864) );
  nor2_1 U10192 ( .ip1(n8855), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[10]), .op(n8857) );
  nor2_1 U10193 ( .ip1(n8857), .ip2(n8856), .op(n8870) );
  nand2_1 U10194 ( .ip1(n8858), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[9]), .op(n8861) );
  nor2_1 U10195 ( .ip1(n8858), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[9]), .op(n8868) );
  nand2_1 U10196 ( .ip1(n5259), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[8]), .op(n8859) );
  or2_1 U10197 ( .ip1(n8868), .ip2(n8859), .op(n8860) );
  nand2_1 U10198 ( .ip1(n8861), .ip2(n8860), .op(n8862) );
  and2_1 U10199 ( .ip1(n8870), .ip2(n8862), .op(n8863) );
  nor2_1 U10200 ( .ip1(n8864), .ip2(n8863), .op(n8865) );
  or2_1 U10201 ( .ip1(n8872), .ip2(n8865), .op(n8866) );
  nand2_1 U10202 ( .ip1(n8867), .ip2(n8866), .op(n8910) );
  nor2_1 U10203 ( .ip1(n5259), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[8]), .op(n8869) );
  nor2_1 U10204 ( .ip1(n8869), .ip2(n8868), .op(n8871) );
  nand2_1 U10205 ( .ip1(n8871), .ip2(n8870), .op(n8873) );
  nor2_1 U10206 ( .ip1(n8873), .ip2(n8872), .op(n8908) );
  nand2_1 U10207 ( .ip1(n5266), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[7]), .op(n8876) );
  nor2_1 U10208 ( .ip1(n5266), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[7]), .op(n8877) );
  nand2_1 U10209 ( .ip1(n5278), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[6]), .op(n8874) );
  or2_1 U10210 ( .ip1(n8877), .ip2(n8874), .op(n8875) );
  nand2_1 U10211 ( .ip1(n8876), .ip2(n8875), .op(n8885) );
  nor2_1 U10212 ( .ip1(n5278), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[6]), .op(n8878) );
  nor2_1 U10213 ( .ip1(n8878), .ip2(n8877), .op(n8901) );
  nand2_1 U10214 ( .ip1(n8879), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[5]), .op(n8882) );
  nor2_1 U10215 ( .ip1(n8879), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[5]), .op(n8899) );
  nand2_1 U10216 ( .ip1(n8457), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[4]), .op(n8880) );
  or2_1 U10217 ( .ip1(n8899), .ip2(n8880), .op(n8881) );
  nand2_1 U10218 ( .ip1(n8882), .ip2(n8881), .op(n8883) );
  and2_1 U10219 ( .ip1(n8901), .ip2(n8883), .op(n8884) );
  nor2_1 U10220 ( .ip1(n8885), .ip2(n8884), .op(n8906) );
  nand2_1 U10221 ( .ip1(n8442), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[3]), .op(n8888) );
  nor2_1 U10222 ( .ip1(n8442), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[3]), .op(n8893) );
  nand2_1 U10223 ( .ip1(n5280), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[2]), .op(n8886) );
  or2_1 U10224 ( .ip1(n8893), .ip2(n8886), .op(n8887) );
  nand2_1 U10225 ( .ip1(n8888), .ip2(n8887), .op(n8898) );
  nand2_1 U10226 ( .ip1(n5245), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[1]), .op(n8892) );
  nor2_1 U10227 ( .ip1(n5245), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[1]), .op(n8890) );
  or2_1 U10228 ( .ip1(n8889), .ip2(n8890), .op(n8891) );
  nand2_1 U10229 ( .ip1(n8892), .ip2(n8891), .op(n8896) );
  nor2_1 U10230 ( .ip1(n5280), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[2]), .op(n8894) );
  nor2_1 U10231 ( .ip1(n8894), .ip2(n8893), .op(n8895) );
  and2_1 U10232 ( .ip1(n8896), .ip2(n8895), .op(n8897) );
  nor2_1 U10233 ( .ip1(n8898), .ip2(n8897), .op(n8904) );
  nor2_1 U10234 ( .ip1(n8457), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[4]), .op(n8900) );
  nor2_1 U10235 ( .ip1(n8900), .ip2(n8899), .op(n8902) );
  nand2_1 U10236 ( .ip1(n8902), .ip2(n8901), .op(n8903) );
  or2_1 U10237 ( .ip1(n8904), .ip2(n8903), .op(n8905) );
  nand2_1 U10238 ( .ip1(n8906), .ip2(n8905), .op(n8907) );
  and2_1 U10239 ( .ip1(n8908), .ip2(n8907), .op(n8909) );
  nor2_1 U10240 ( .ip1(n8910), .ip2(n8909), .op(n8912) );
  nand2_1 U10241 ( .ip1(n8912), .ip2(n8911), .op(n8913) );
  nor2_1 U10242 ( .ip1(n8965), .ip2(n8916), .op(n5059) );
  nand2_1 U10243 ( .ip1(n8962), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[0]), .op(n8919) );
  xor2_1 U10244 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[1]), .ip2(
        n8919), .op(n8917) );
  nor2_1 U10245 ( .ip1(n8965), .ip2(n8917), .op(n5058) );
  inv_1 U10246 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[2]), .op(
        n8922) );
  inv_1 U10247 ( .ip(n8919), .op(n8918) );
  nand2_1 U10248 ( .ip1(n8918), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[1]), .op(n8921) );
  nand2_1 U10249 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[1]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[2]), .op(n8920) );
  not_ab_or_c_or_d U10250 ( .ip1(n8922), .ip2(n8921), .ip3(n8924), .ip4(n8965), 
        .op(n5057) );
  inv_1 U10251 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[3]), .op(
        n8923) );
  nor2_1 U10252 ( .ip1(n8965), .ip2(n5263), .op(n5056) );
  nand2_1 U10253 ( .ip1(n8924), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[3]), .op(n8927) );
  xor2_1 U10254 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[4]), .ip2(
        n8927), .op(n8925) );
  nor2_1 U10255 ( .ip1(n8965), .ip2(n8925), .op(n5055) );
  inv_1 U10256 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[5]), .op(
        n8930) );
  inv_1 U10257 ( .ip(n8927), .op(n8926) );
  nand2_1 U10258 ( .ip1(n8926), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[4]), .op(n8929) );
  nand2_1 U10259 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[4]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[5]), .op(n8928) );
  not_ab_or_c_or_d U10260 ( .ip1(n8930), .ip2(n8929), .ip3(n8933), .ip4(n8965), 
        .op(n5054) );
  inv_1 U10261 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[6]), .op(
        n8931) );
  xor2_1 U10262 ( .ip1(n8931), .ip2(n8933), .op(n8932) );
  xor2_1 U10263 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[7]), .ip2(
        n8936), .op(n8934) );
  inv_1 U10264 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[8]), .op(
        n8939) );
  inv_1 U10265 ( .ip(n8936), .op(n8935) );
  nand2_1 U10266 ( .ip1(n8935), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[7]), .op(n8938) );
  nand2_1 U10267 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[7]), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[8]), .op(n8937) );
  nor2_1 U10268 ( .ip1(n8937), .ip2(n8936), .op(n8942) );
  not_ab_or_c_or_d U10269 ( .ip1(n8939), .ip2(n8938), .ip3(n8942), .ip4(n8965), 
        .op(n5051) );
  inv_1 U10270 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[9]), .op(
        n8940) );
  nor2_1 U10271 ( .ip1(n8965), .ip2(n8941), .op(n5050) );
  nand2_1 U10272 ( .ip1(n8942), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[9]), .op(n8945) );
  xor2_1 U10273 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[10]), .ip2(
        n8945), .op(n8943) );
  nor2_1 U10274 ( .ip1(n8965), .ip2(n8943), .op(n5049) );
  inv_1 U10275 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[11]), .op(
        n8948) );
  inv_1 U10276 ( .ip(n8945), .op(n8944) );
  nand2_1 U10277 ( .ip1(n8944), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[10]), .op(n8947) );
  nand2_1 U10278 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[10]), 
        .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[11]), .op(n8946) );
  nor2_1 U10279 ( .ip1(n8946), .ip2(n8945), .op(n8952) );
  not_ab_or_c_or_d U10280 ( .ip1(n8948), .ip2(n8947), .ip3(n8952), .ip4(n8965), 
        .op(n5048) );
  inv_1 U10281 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[12]), .op(
        n8949) );
  xnor2_1 U10282 ( .ip1(n8949), .ip2(n8952), .op(n8950) );
  inv_1 U10283 ( .ip(n8950), .op(n8951) );
  nor2_1 U10284 ( .ip1(n8965), .ip2(n8951), .op(n5047) );
  nand2_1 U10285 ( .ip1(n8952), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[12]), .op(n8955) );
  xor2_1 U10286 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[13]), .ip2(
        n8955), .op(n8953) );
  nor2_1 U10287 ( .ip1(n8965), .ip2(n8953), .op(n5046) );
  inv_1 U10288 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[14]), .op(
        n8958) );
  inv_1 U10289 ( .ip(n8955), .op(n8954) );
  nand2_1 U10290 ( .ip1(n8954), .ip2(
        i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[13]), .op(n8957) );
  nand2_1 U10291 ( .ip1(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[13]), 
        .ip2(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[14]), .op(n8956) );
  nor2_1 U10292 ( .ip1(n8956), .ip2(n8955), .op(n8959) );
  not_ab_or_c_or_d U10293 ( .ip1(n8958), .ip2(n8957), .ip3(n8959), .ip4(n8965), 
        .op(n5045) );
  inv_1 U10294 ( .ip(i_i2c_U_DW_apb_i2c_clk_gen_scl_p_setup_cntr[15]), .op(
        n8960) );
  nor2_1 U10295 ( .ip1(n8965), .ip2(n8961), .op(n5060) );
  inv_1 U10296 ( .ip(n8962), .op(n8963) );
  nor2_1 U10297 ( .ip1(i_i2c_scl_p_setup_cmplt), .ip2(n8963), .op(n8964) );
  nor2_1 U10298 ( .ip1(n8965), .ip2(n8964), .op(n5044) );
  not_ab_or_c_or_d U10299 ( .ip1(n9502), .ip2(n8989), .ip3(n8988), .ip4(n8966), 
        .op(n8971) );
  or3_1 U10300 ( .ip1(n11126), .ip2(n8968), .ip3(n8967), .op(n8970) );
  nor2_1 U10301 ( .ip1(i_i2c_re_start_en), .ip2(n8971), .op(n8969) );
  not_ab_or_c_or_d U10302 ( .ip1(i_i2c_byte_wait_scl), .ip2(n8971), .ip3(n8970), .ip4(n8969), .op(n5192) );
  inv_1 U10303 ( .ip(i_i2c_mst_rx_bwen), .op(n8972) );
  nor2_1 U10304 ( .ip1(n8972), .ip2(n11037), .op(n8975) );
  nor2_1 U10305 ( .ip1(n8973), .ip2(n8976), .op(n8974) );
  mux2_1 U10306 ( .ip1(n8975), .ip2(i_i2c_rx_scl_hcnt_en), .s(n8974), .op(
        n4160) );
  inv_1 U10307 ( .ip(i_i2c_scl_hcnt_en), .op(n8981) );
  nand2_1 U10308 ( .ip1(n11047), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[3]), .op(n9323) );
  nor2_1 U10309 ( .ip1(n9323), .ip2(n8976), .op(n8980) );
  nand2_1 U10310 ( .ip1(n8977), .ip2(n11040), .op(n8978) );
  nor2_1 U10311 ( .ip1(n8978), .ip2(n5591), .op(n11048) );
  nor2_1 U10312 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_mst_tx_bwen), .ip2(n8980), 
        .op(n8979) );
  not_ab_or_c_or_d U10313 ( .ip1(n8981), .ip2(n8980), .ip3(n11048), .ip4(n8979), .op(n4127) );
  inv_1 U10314 ( .ip(n8982), .op(n9321) );
  nand2_1 U10315 ( .ip1(n11834), .ip2(i_i2c_mst_tx_ack_vld), .op(n8983) );
  nand2_1 U10316 ( .ip1(n9321), .ip2(n8983), .op(n4172) );
  nor2_1 U10317 ( .ip1(i_i2c_ic_enable_sync), .ip2(i_i2c_mst_activity), .op(
        n8984) );
  nor2_1 U10318 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv), .ip2(n8984), .op(n8986) );
  nand2_1 U10319 ( .ip1(n8986), .ip2(n8985), .op(n9503) );
  nor2_1 U10320 ( .ip1(n9503), .ip2(n8987), .op(i_i2c_U_DW_apb_i2c_mstfsm_N72)
         );
  nor2_1 U10321 ( .ip1(n9503), .ip2(n8988), .op(i_i2c_U_DW_apb_i2c_mstfsm_N75)
         );
  inv_1 U10322 ( .ip(n8989), .op(n8990) );
  nor2_1 U10323 ( .ip1(n9503), .ip2(n8990), .op(i_i2c_U_DW_apb_i2c_mstfsm_N74)
         );
  nor2_1 U10324 ( .ip1(n9503), .ip2(n8991), .op(i_i2c_U_DW_apb_i2c_mstfsm_N76)
         );
  inv_1 U10325 ( .ip(n8992), .op(n8996) );
  nor3_1 U10326 ( .ip1(i_i2c_scl_s_setup_cmplt), .ip2(i_i2c_scl_s_hld_cmplt), 
        .ip3(n8993), .op(n8995) );
  ab_or_c_or_d U10327 ( .ip1(n8996), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda), .ip3(n8995), .ip4(n8994), 
        .op(n4953) );
  nor2_1 U10328 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_st_scl_s_hld_en), .ip2(
        i_i2c_start_en), .op(n4956) );
  nand2_1 U10329 ( .ip1(i_i2c_U_dff_tx_mem[63]), .ip2(n10182), .op(n9005) );
  and2_1 U10330 ( .ip1(i_i2c_U_dff_tx_mem[0]), .ip2(n11214), .op(n9002) );
  nand2_1 U10331 ( .ip1(i_i2c_U_dff_tx_mem[36]), .ip2(n10190), .op(n9000) );
  nand2_1 U10332 ( .ip1(i_i2c_U_dff_tx_mem[9]), .ip2(n10189), .op(n8999) );
  nand2_1 U10333 ( .ip1(i_i2c_U_dff_tx_mem[18]), .ip2(n10179), .op(n8998) );
  nand2_1 U10334 ( .ip1(i_i2c_U_dff_tx_mem[27]), .ip2(n10180), .op(n8997) );
  nand4_1 U10335 ( .ip1(n9000), .ip2(n8999), .ip3(n8998), .ip4(n8997), .op(
        n9001) );
  not_ab_or_c_or_d U10336 ( .ip1(i_i2c_U_dff_tx_mem[45]), .ip2(n10178), .ip3(
        n9002), .ip4(n9001), .op(n9004) );
  nand2_1 U10337 ( .ip1(i_i2c_U_dff_tx_mem[54]), .ip2(n10181), .op(n9003) );
  nand3_1 U10338 ( .ip1(n9005), .ip2(n9004), .ip3(n9003), .op(n9006) );
  mux2_1 U10339 ( .ip1(i_i2c_tx_fifo_data_buf[0]), .ip2(n9006), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .op(n5222) );
  nand2_1 U10340 ( .ip1(i_i2c_U_dff_tx_mem[55]), .ip2(n10181), .op(n9015) );
  and2_1 U10341 ( .ip1(n11214), .ip2(i_i2c_U_dff_tx_mem[1]), .op(n9012) );
  nand2_1 U10342 ( .ip1(n10180), .ip2(i_i2c_U_dff_tx_mem[28]), .op(n9010) );
  nand2_1 U10343 ( .ip1(n10178), .ip2(i_i2c_U_dff_tx_mem[46]), .op(n9009) );
  nand2_1 U10344 ( .ip1(n10179), .ip2(i_i2c_U_dff_tx_mem[19]), .op(n9008) );
  nand2_1 U10345 ( .ip1(n10182), .ip2(i_i2c_U_dff_tx_mem[64]), .op(n9007) );
  nand4_1 U10346 ( .ip1(n9010), .ip2(n9009), .ip3(n9008), .ip4(n9007), .op(
        n9011) );
  not_ab_or_c_or_d U10347 ( .ip1(i_i2c_U_dff_tx_mem[37]), .ip2(n10190), .ip3(
        n9012), .ip4(n9011), .op(n9014) );
  nand2_1 U10348 ( .ip1(n10189), .ip2(i_i2c_U_dff_tx_mem[10]), .op(n9013) );
  nand3_1 U10349 ( .ip1(n9015), .ip2(n9014), .ip3(n9013), .op(n9016) );
  mux2_1 U10350 ( .ip1(i_i2c_tx_fifo_data_buf[1]), .ip2(n9016), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .op(n5221) );
  nand2_1 U10351 ( .ip1(i_i2c_U_dff_tx_mem[56]), .ip2(n10181), .op(n9025) );
  and2_1 U10352 ( .ip1(n11214), .ip2(i_i2c_U_dff_tx_mem[2]), .op(n9022) );
  nand2_1 U10353 ( .ip1(n10178), .ip2(i_i2c_U_dff_tx_mem[47]), .op(n9020) );
  nand2_1 U10354 ( .ip1(n10180), .ip2(i_i2c_U_dff_tx_mem[29]), .op(n9019) );
  nand2_1 U10355 ( .ip1(n10182), .ip2(i_i2c_U_dff_tx_mem[65]), .op(n9018) );
  nand2_1 U10356 ( .ip1(n10179), .ip2(i_i2c_U_dff_tx_mem[20]), .op(n9017) );
  nand4_1 U10357 ( .ip1(n9020), .ip2(n9019), .ip3(n9018), .ip4(n9017), .op(
        n9021) );
  not_ab_or_c_or_d U10358 ( .ip1(i_i2c_U_dff_tx_mem[11]), .ip2(n10189), .ip3(
        n9022), .ip4(n9021), .op(n9024) );
  nand2_1 U10359 ( .ip1(n10190), .ip2(i_i2c_U_dff_tx_mem[38]), .op(n9023) );
  nand3_1 U10360 ( .ip1(n9025), .ip2(n9024), .ip3(n9023), .op(n9026) );
  mux2_1 U10361 ( .ip1(i_i2c_tx_fifo_data_buf[2]), .ip2(n9026), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .op(n5220) );
  nand2_1 U10362 ( .ip1(i_i2c_U_dff_tx_mem[52]), .ip2(n10178), .op(n9035) );
  and2_1 U10363 ( .ip1(n11214), .ip2(i_i2c_U_dff_tx_mem[7]), .op(n9032) );
  nand2_1 U10364 ( .ip1(n10189), .ip2(i_i2c_U_dff_tx_mem[16]), .op(n9030) );
  nand2_1 U10365 ( .ip1(n10180), .ip2(i_i2c_U_dff_tx_mem[34]), .op(n9029) );
  nand2_1 U10366 ( .ip1(n10182), .ip2(i_i2c_U_dff_tx_mem[70]), .op(n9028) );
  nand2_1 U10367 ( .ip1(n10181), .ip2(i_i2c_U_dff_tx_mem[61]), .op(n9027) );
  nand4_1 U10368 ( .ip1(n9030), .ip2(n9029), .ip3(n9028), .ip4(n9027), .op(
        n9031) );
  not_ab_or_c_or_d U10369 ( .ip1(n10179), .ip2(i_i2c_U_dff_tx_mem[25]), .ip3(
        n9032), .ip4(n9031), .op(n9034) );
  nand2_1 U10370 ( .ip1(n10190), .ip2(i_i2c_U_dff_tx_mem[43]), .op(n9033) );
  nand3_1 U10371 ( .ip1(n9035), .ip2(n9034), .ip3(n9033), .op(n9036) );
  mux2_1 U10372 ( .ip1(i_i2c_tx_fifo_data_buf[7]), .ip2(n9036), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .op(n5215) );
  inv_1 U10373 ( .ip(i_i2c_slv_tx_ready_unconn), .op(n9038) );
  nor3_1 U10374 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[3]), .ip2(
        n9038), .ip3(n9037), .op(n9059) );
  nand2_1 U10375 ( .ip1(n9059), .ip2(n9039), .op(n9040) );
  nand3_1 U10376 ( .ip1(n9040), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_ready_dly1), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_data_sda), .op(n9062) );
  not_ab_or_c_or_d U10377 ( .ip1(i_i2c_tx_fifo_data_buf[7]), .ip2(n9055), 
        .ip3(n9041), .ip4(n9497), .op(n9061) );
  inv_1 U10378 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[2]), .op(
        n9045) );
  inv_1 U10379 ( .ip(i_i2c_tx_fifo_data_buf[1]), .op(n9043) );
  nor2_1 U10380 ( .ip1(i_i2c_tx_fifo_data_buf[2]), .ip2(n9052), .op(n9042) );
  not_ab_or_c_or_d U10381 ( .ip1(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[1]), .ip2(n9043), .ip3(
        n9042), .ip4(n9046), .op(n9044) );
  not_ab_or_c_or_d U10382 ( .ip1(i_i2c_tx_fifo_data_buf[0]), .ip2(n9046), 
        .ip3(n9045), .ip4(n9044), .op(n9057) );
  nor2_1 U10383 ( .ip1(i_i2c_tx_fifo_data_buf[3]), .ip2(n9049), .op(n9056) );
  inv_1 U10384 ( .ip(i_i2c_tx_fifo_data_buf[5]), .op(n10897) );
  nor2_1 U10385 ( .ip1(i_i2c_tx_fifo_data_buf[4]), .ip2(n9047), .op(n9051) );
  or2_1 U10386 ( .ip1(i_i2c_tx_fifo_data_buf[6]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[1]), .op(n9048) );
  nand2_1 U10387 ( .ip1(n9049), .ip2(n9048), .op(n9050) );
  not_ab_or_c_or_d U10388 ( .ip1(n9052), .ip2(n10897), .ip3(n9051), .ip4(n9050), .op(n9053) );
  nor2_1 U10389 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_slv_tx_bit_count[2]), .ip2(
        n9053), .op(n9054) );
  nor4_1 U10390 ( .ip1(n9057), .ip2(n9056), .ip3(n9055), .ip4(n9054), .op(
        n9058) );
  nand2_1 U10391 ( .ip1(n9059), .ip2(n9058), .op(n9060) );
  nand3_1 U10392 ( .ip1(n9062), .ip2(n9061), .ip3(n9060), .op(n5103) );
  mux2_1 U10393 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[7]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[5]), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[1]), .op(n9075) );
  nor2_1 U10394 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[2]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[0]), .op(n9074) );
  inv_1 U10395 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[1]), .op(n10914)
         );
  nor2_1 U10396 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[3]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[1]), .op(n9063) );
  not_ab_or_c_or_d U10397 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[1]), 
        .ip2(n10914), .ip3(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[0]), .ip4(
        n9063), .op(n9066) );
  and3_1 U10398 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[0]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[2]), .ip3(n9064), .op(n9065)
         );
  not_ab_or_c_or_d U10399 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[0]), 
        .ip2(n9067), .ip3(n9066), .ip4(n9065), .op(n9069) );
  nor2_1 U10400 ( .ip1(n9069), .ip2(n9068), .op(n9073) );
  mux2_1 U10401 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[6]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[4]), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[1]), .op(n9070) );
  nand2_1 U10402 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[0]), .ip2(
        n9070), .op(n9071) );
  nor2_1 U10403 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[2]), .ip2(
        n9071), .op(n9072) );
  not_ab_or_c_or_d U10404 ( .ip1(n9075), .ip2(n9074), .ip3(n9073), .ip4(n9072), 
        .op(n9078) );
  inv_1 U10405 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_data_sda), .op(n9077) );
  nand2_1 U10406 ( .ip1(n11048), .ip2(i_i2c_debug_wr), .op(n9076) );
  mux2_1 U10407 ( .ip1(n9078), .ip2(n9077), .s(n9076), .op(n9079) );
  nand3_1 U10408 ( .ip1(n9321), .ip2(n11834), .ip3(n9079), .op(n4116) );
  inv_1 U10409 ( .ip(i_i2c_ic_clk_oe), .op(n9344) );
  mux2_1 U10410 ( .ip1(n9344), .ip2(n6352), .s(
        i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv), .op(n9469) );
  nand2_1 U10411 ( .ip1(n11858), .ip2(
        i_i2c_U_DW_apb_i2c_mstfsm_mst_gen_ack_en_r), .op(n9082) );
  nand2_1 U10412 ( .ip1(n9080), .ip2(
        i_i2c_U_DW_apb_i2c_slvfsm_ic_enable_sync_vld), .op(n9081) );
  nand2_1 U10413 ( .ip1(n9082), .ip2(n9081), .op(n9341) );
  inv_1 U10414 ( .ip(n9469), .op(n9342) );
  inv_1 U10415 ( .ip(i_i2c_ic_sda_tx_hold_sync[0]), .op(n9108) );
  nand2_1 U10416 ( .ip1(n9469), .ip2(n9108), .op(n9091) );
  nor4_1 U10417 ( .ip1(i_i2c_ic_sda_tx_hold_sync[14]), .ip2(
        i_i2c_ic_sda_tx_hold_sync[13]), .ip3(i_i2c_ic_sda_tx_hold_sync[12]), 
        .ip4(i_i2c_ic_sda_tx_hold_sync[10]), .op(n9084) );
  nor3_1 U10418 ( .ip1(i_i2c_ic_sda_tx_hold_sync[11]), .ip2(
        i_i2c_ic_sda_tx_hold_sync[9]), .ip3(i_i2c_ic_sda_tx_hold_sync[15]), 
        .op(n9083) );
  and2_1 U10419 ( .ip1(n9084), .ip2(n9083), .op(n9097) );
  nor2_1 U10420 ( .ip1(i_i2c_ic_sda_tx_hold_sync[5]), .ip2(
        i_i2c_ic_sda_tx_hold_sync[6]), .op(n9087) );
  inv_1 U10421 ( .ip(i_i2c_ic_sda_tx_hold_sync[8]), .op(n9086) );
  nand2_1 U10422 ( .ip1(i_i2c_ic_sda_tx_hold_sync[0]), .ip2(
        i_i2c_ic_sda_tx_hold_sync[1]), .op(n9085) );
  nand3_1 U10423 ( .ip1(n9087), .ip2(n9086), .ip3(n9085), .op(n9089) );
  inv_1 U10424 ( .ip(i_i2c_ic_sda_tx_hold_sync[4]), .op(n9119) );
  inv_1 U10425 ( .ip(i_i2c_ic_sda_tx_hold_sync[3]), .op(n9114) );
  inv_1 U10426 ( .ip(i_i2c_ic_sda_tx_hold_sync[2]), .op(n9107) );
  inv_1 U10427 ( .ip(i_i2c_ic_sda_tx_hold_sync[7]), .op(n9102) );
  nand4_1 U10428 ( .ip1(n9119), .ip2(n9114), .ip3(n9107), .ip4(n9102), .op(
        n9088) );
  nor2_1 U10429 ( .ip1(n9089), .ip2(n9088), .op(n9090) );
  and2_1 U10430 ( .ip1(n9097), .ip2(n9090), .op(n9304) );
  nand2_1 U10431 ( .ip1(n9091), .ip2(n9304), .op(n9308) );
  mux2_1 U10432 ( .ip1(n9093), .ip2(n9092), .s(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r), .op(n9154) );
  mux2_1 U10433 ( .ip1(n9095), .ip2(n9094), .s(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r), .op(n9161) );
  mux2_1 U10434 ( .ip1(i_i2c_ic_fs_spklen[3]), .ip2(i_i2c_ic_hs_spklen[3]), 
        .s(i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r), .op(n9105) );
  nand2_1 U10435 ( .ip1(n9106), .ip2(n9105), .op(n9124) );
  mux2_1 U10436 ( .ip1(i_i2c_ic_fs_spklen[5]), .ip2(i_i2c_ic_hs_spklen[5]), 
        .s(i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r), .op(n9129) );
  nand2_1 U10437 ( .ip1(n9138), .ip2(n9101), .op(n9096) );
  nand2_1 U10438 ( .ip1(n9096), .ip2(i_i2c_ic_sda_tx_hold_sync[8]), .op(n9098)
         );
  nand2_1 U10439 ( .ip1(n9132), .ip2(n9154), .op(n9099) );
  nand2_1 U10440 ( .ip1(n9149), .ip2(i_i2c_ic_sda_tx_hold_sync[7]), .op(n9137)
         );
  nand2_1 U10441 ( .ip1(n9099), .ip2(n9137), .op(n9100) );
  nor2_1 U10442 ( .ip1(n9100), .ip2(n9138), .op(n9146) );
  nor2_1 U10443 ( .ip1(n9146), .ip2(n9104), .op(n9136) );
  inv_1 U10444 ( .ip(n9105), .op(n9165) );
  xnor2_1 U10445 ( .ip1(n9106), .ip2(n9165), .op(n9115) );
  nor2_1 U10446 ( .ip1(i_i2c_ic_sda_tx_hold_sync[2]), .ip2(n9106), .op(n9113)
         );
  mux2_1 U10447 ( .ip1(i_i2c_ic_fs_spklen[1]), .ip2(i_i2c_ic_hs_spklen[1]), 
        .s(i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r), .op(n9177) );
  inv_1 U10448 ( .ip(n9177), .op(n9111) );
  inv_1 U10449 ( .ip(n9106), .op(n9175) );
  mux2_1 U10450 ( .ip1(i_i2c_ic_fs_spklen[0]), .ip2(i_i2c_ic_hs_spklen[0]), 
        .s(i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r), .op(n9182) );
  not_ab_or_c_or_d U10451 ( .ip1(n5539), .ip2(n5572), .ip3(n9182), .ip4(n9108), 
        .op(n9109) );
  not_ab_or_c_or_d U10452 ( .ip1(i_i2c_ic_sda_tx_hold_sync[1]), .ip2(n9111), 
        .ip3(n9109), .ip4(n9110), .op(n9112) );
  ab_or_c_or_d U10453 ( .ip1(n9114), .ip2(n9115), .ip3(n9113), .ip4(n9112), 
        .op(n9118) );
  inv_1 U10454 ( .ip(n9115), .op(n9116) );
  nand2_1 U10455 ( .ip1(n9116), .ip2(i_i2c_ic_sda_tx_hold_sync[3]), .op(n9117)
         );
  nand2_1 U10456 ( .ip1(n9117), .ip2(n9118), .op(n9122) );
  xor2_1 U10457 ( .ip1(n9161), .ip2(n9124), .op(n9120) );
  nand2_1 U10458 ( .ip1(n9120), .ip2(n9119), .op(n9121) );
  inv_1 U10459 ( .ip(n9123), .op(n9130) );
  nand2_1 U10460 ( .ip1(n9124), .ip2(n9161), .op(n9125) );
  nand2_1 U10461 ( .ip1(n9130), .ip2(n9125), .op(n9126) );
  nand2_1 U10462 ( .ip1(n9126), .ip2(i_i2c_ic_sda_tx_hold_sync[4]), .op(n9127)
         );
  inv_1 U10463 ( .ip(n9129), .op(n9156) );
  nand2_1 U10464 ( .ip1(n9130), .ip2(n9156), .op(n9131) );
  nand2_1 U10465 ( .ip1(n9132), .ip2(n9131), .op(n9133) );
  fulladder U10466 ( .a(i_i2c_ic_sda_tx_hold_sync[5]), .b(n9134), .ci(n9133), 
        .co(n9135) );
  nor2_1 U10467 ( .ip1(n9136), .ip2(n9135), .op(n9145) );
  nor2_1 U10468 ( .ip1(i_i2c_ic_sda_tx_hold_sync[7]), .ip2(n9149), .op(n9142)
         );
  inv_1 U10469 ( .ip(n9137), .op(n9140) );
  inv_1 U10470 ( .ip(n9138), .op(n9139) );
  nor2_1 U10471 ( .ip1(n9140), .ip2(n9139), .op(n9141) );
  nor2_1 U10472 ( .ip1(n9142), .ip2(n9141), .op(n9143) );
  nor2_1 U10473 ( .ip1(i_i2c_ic_sda_tx_hold_sync[8]), .ip2(n9143), .op(n9144)
         );
  ab_or_c_or_d U10474 ( .ip1(n9146), .ip2(n5573), .ip3(n9145), .ip4(n9144), 
        .op(n9147) );
  nand2_2 U10475 ( .ip1(n5604), .ip2(n9147), .op(n9148) );
  nand2_4 U10476 ( .ip1(n9148), .ip2(
        i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv), .op(n9186) );
  or2_1 U10477 ( .ip1(n9149), .ip2(n9186), .op(n9153) );
  or2_1 U10478 ( .ip1(i_i2c_ic_sda_tx_hold_sync[7]), .ip2(n9153), .op(n9194)
         );
  nand2_1 U10479 ( .ip1(n9194), .ip2(i_i2c_ic_sda_tx_hold_sync[8]), .op(n9281)
         );
  or2_1 U10480 ( .ip1(i_i2c_ic_sda_tx_hold_sync[12]), .ip2(
        i_i2c_ic_sda_tx_hold_sync[11]), .op(n9150) );
  inv_1 U10481 ( .ip(i_i2c_ic_sda_tx_hold_sync[9]), .op(n9280) );
  nand2_1 U10482 ( .ip1(n5525), .ip2(n9280), .op(n9202) );
  nor2_1 U10483 ( .ip1(n9150), .ip2(n9202), .op(n9151) );
  nand2_1 U10484 ( .ip1(n9281), .ip2(n9151), .op(n9201) );
  nor2_1 U10485 ( .ip1(n9201), .ip2(i_i2c_ic_sda_tx_hold_sync[13]), .op(n9197)
         );
  inv_1 U10486 ( .ip(i_i2c_ic_sda_tx_hold_sync[14]), .op(n9152) );
  xnor2_1 U10487 ( .ip1(i_i2c_ic_sda_tx_hold_sync[7]), .ip2(n9153), .op(n9158)
         );
  or2_1 U10488 ( .ip1(n9154), .ip2(n9186), .op(n9155) );
  or2_1 U10489 ( .ip1(i_i2c_ic_sda_tx_hold_sync[6]), .ip2(n9155), .op(n9157)
         );
  nand2_1 U10490 ( .ip1(n9158), .ip2(n9157), .op(n9222) );
  xnor2_1 U10491 ( .ip1(i_i2c_ic_sda_tx_hold_sync[6]), .ip2(n9155), .op(n9168)
         );
  or2_1 U10492 ( .ip1(n9156), .ip2(n9186), .op(n9160) );
  or2_1 U10493 ( .ip1(i_i2c_ic_sda_tx_hold_sync[5]), .ip2(n9160), .op(n9167)
         );
  nand2_1 U10494 ( .ip1(n9168), .ip2(n9167), .op(n9229) );
  nor2_1 U10495 ( .ip1(n9158), .ip2(n9157), .op(n9221) );
  or2_1 U10496 ( .ip1(n9229), .ip2(n9221), .op(n9159) );
  nand2_1 U10497 ( .ip1(n9222), .ip2(n9159), .op(n9169) );
  or2_1 U10498 ( .ip1(n9161), .ip2(n9186), .op(n9164) );
  or2_1 U10499 ( .ip1(i_i2c_ic_sda_tx_hold_sync[4]), .ip2(n9164), .op(n9162)
         );
  nand2_1 U10500 ( .ip1(n9163), .ip2(n9162), .op(n9235) );
  xnor2_1 U10501 ( .ip1(i_i2c_ic_sda_tx_hold_sync[4]), .ip2(n9164), .op(n9171)
         );
  or2_1 U10502 ( .ip1(i_i2c_ic_sda_tx_hold_sync[3]), .ip2(n9174), .op(n9170)
         );
  nand2_1 U10503 ( .ip1(n9171), .ip2(n9170), .op(n9240) );
  inv_1 U10504 ( .ip(n9240), .op(n9234) );
  nor2_1 U10505 ( .ip1(n9168), .ip2(n9167), .op(n9217) );
  nor2_1 U10506 ( .ip1(n9217), .ip2(n9221), .op(n9173) );
  nor2_1 U10507 ( .ip1(n9171), .ip2(n9170), .op(n9239) );
  nor2_1 U10508 ( .ip1(n9239), .ip2(n9172), .op(n9216) );
  nand2_1 U10509 ( .ip1(n9216), .ip2(n9173), .op(n9192) );
  or2_1 U10510 ( .ip1(i_i2c_ic_sda_tx_hold_sync[2]), .ip2(n5564), .op(n9189)
         );
  nand2_1 U10511 ( .ip1(n9189), .ip2(n9188), .op(n9247) );
  xnor2_1 U10512 ( .ip1(i_i2c_ic_sda_tx_hold_sync[2]), .ip2(n5564), .op(n9187)
         );
  nand2_1 U10513 ( .ip1(n9187), .ip2(n9186), .op(n9250) );
  inv_1 U10514 ( .ip(n9186), .op(n9178) );
  nand2_1 U10515 ( .ip1(n9178), .ip2(n9177), .op(n9180) );
  or2_1 U10516 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv), .ip2(n9304), 
        .op(n9179) );
  nand2_1 U10517 ( .ip1(n9179), .ip2(n9180), .op(n9181) );
  nand2_1 U10518 ( .ip1(n9184), .ip2(i_i2c_ic_sda_tx_hold_sync[1]), .op(n9256)
         );
  inv_1 U10519 ( .ip(n9182), .op(n9183) );
  or2_1 U10520 ( .ip1(n9183), .ip2(n9186), .op(n9260) );
  nor2_1 U10521 ( .ip1(i_i2c_ic_sda_tx_hold_sync[0]), .ip2(n9260), .op(n9258)
         );
  or2_1 U10522 ( .ip1(n9258), .ip2(n9255), .op(n9185) );
  nor2_1 U10523 ( .ip1(n9186), .ip2(n5566), .op(n9244) );
  or2_1 U10524 ( .ip1(n9194), .ip2(i_i2c_ic_sda_tx_hold_sync[8]), .op(n9211)
         );
  xnor2_2 U10525 ( .ip1(i_i2c_ic_sda_tx_hold_sync[15]), .ip2(n9196), .op(n9348) );
  and2_1 U10526 ( .ip1(n9348), .ip2(n9347), .op(n9303) );
  inv_1 U10527 ( .ip(n9197), .op(n9198) );
  nor2_1 U10528 ( .ip1(n9348), .ip2(n9347), .op(n9200) );
  nor3_1 U10529 ( .ip1(n9349), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[14]), .ip3(n9200), .op(
        n9302) );
  and2_1 U10530 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[14]), 
        .ip2(n9349), .op(n9199) );
  or2_1 U10531 ( .ip1(n9200), .ip2(n9199), .op(n9296) );
  nand2_1 U10532 ( .ip1(n9441), .ip2(n5516), .op(n9207) );
  nor2_1 U10533 ( .ip1(n5516), .ip2(n9441), .op(n9297) );
  nor2_1 U10534 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[12]), 
        .ip2(n9297), .op(n9205) );
  inv_1 U10535 ( .ip(n9281), .op(n9214) );
  nor2_1 U10536 ( .ip1(n9214), .ip2(n9202), .op(n9209) );
  inv_1 U10537 ( .ip(i_i2c_ic_sda_tx_hold_sync[11]), .op(n9203) );
  nand2_1 U10538 ( .ip1(n9205), .ip2(n9415), .op(n9206) );
  and2_1 U10539 ( .ip1(n9207), .ip2(n9206), .op(n9208) );
  nor2_1 U10540 ( .ip1(n9296), .ip2(n9208), .op(n9301) );
  inv_1 U10541 ( .ip(n9209), .op(n9210) );
  nor2_1 U10542 ( .ip1(n9398), .ip2(n9461), .op(n9291) );
  nand2_1 U10543 ( .ip1(n9211), .ip2(n9281), .op(n9213) );
  nor2_1 U10544 ( .ip1(n9383), .ip2(n9382), .op(n9286) );
  inv_1 U10545 ( .ip(n9217), .op(n9230) );
  nand2_1 U10546 ( .ip1(n9228), .ip2(n9230), .op(n9215) );
  nand2_1 U10547 ( .ip1(n9229), .ip2(n9215), .op(n9220) );
  inv_1 U10548 ( .ip(n9216), .op(n9226) );
  nor2_1 U10549 ( .ip1(n9226), .ip2(n9217), .op(n9218) );
  inv_1 U10550 ( .ip(n9232), .op(n9242) );
  and2_1 U10551 ( .ip1(n9218), .ip2(n9242), .op(n9219) );
  nor2_1 U10552 ( .ip1(n9220), .ip2(n9219), .op(n9225) );
  inv_1 U10553 ( .ip(n9221), .op(n9223) );
  nand2_1 U10554 ( .ip1(n9223), .ip2(n9222), .op(n9224) );
  xor2_1 U10555 ( .ip1(n9225), .ip2(n9224), .op(n9379) );
  nand2_1 U10556 ( .ip1(n9230), .ip2(n9229), .op(n9231) );
  inv_1 U10557 ( .ip(n9375), .op(n9276) );
  nor2_1 U10558 ( .ip1(n9379), .ip2(n9434), .op(n9274) );
  nor3_1 U10559 ( .ip1(n9276), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[6]), .ip3(n9274), .op(
        n9278) );
  inv_1 U10560 ( .ip(n9239), .op(n9241) );
  nand2_1 U10561 ( .ip1(n9241), .ip2(n9240), .op(n9243) );
  xnor2_1 U10562 ( .ip1(n9243), .ip2(n9242), .op(n9368) );
  nor2_1 U10563 ( .ip1(n9374), .ip2(n9450), .op(n9271) );
  inv_1 U10564 ( .ip(n9244), .op(n9251) );
  nand2_1 U10565 ( .ip1(n9251), .ip2(n9252), .op(n9245) );
  nand2_1 U10566 ( .ip1(n9250), .ip2(n9245), .op(n9249) );
  nand2_1 U10567 ( .ip1(n5563), .ip2(n9247), .op(n9248) );
  nand2_1 U10568 ( .ip1(n9251), .ip2(n9250), .op(n9254) );
  inv_1 U10569 ( .ip(n9252), .op(n9253) );
  xnor2_1 U10570 ( .ip1(n9254), .ip2(n9253), .op(n9363) );
  inv_1 U10571 ( .ip(n9363), .op(n9360) );
  inv_1 U10572 ( .ip(n9255), .op(n9257) );
  nand2_1 U10573 ( .ip1(n9257), .ip2(n9256), .op(n9259) );
  xor2_1 U10574 ( .ip1(n9259), .ip2(n9258), .op(n9357) );
  inv_1 U10575 ( .ip(n9357), .op(n9262) );
  xnor2_1 U10576 ( .ip1(i_i2c_ic_sda_tx_hold_sync[0]), .ip2(n9260), .op(n9354)
         );
  inv_1 U10577 ( .ip(n9354), .op(n9261) );
  not_ab_or_c_or_d U10578 ( .ip1(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[1]), .ip2(n9262), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[0]), .ip4(n9261), .op(
        n9263) );
  nor2_1 U10579 ( .ip1(n9445), .ip2(n9263), .op(n9265) );
  nor2_1 U10580 ( .ip1(n9357), .ip2(n9263), .op(n9264) );
  or2_1 U10581 ( .ip1(n9265), .ip2(n9264), .op(n9266) );
  nor2_1 U10582 ( .ip1(n9365), .ip2(n9364), .op(n9267) );
  not_ab_or_c_or_d U10583 ( .ip1(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[2]), .ip2(n9363), .ip3(
        n9266), .ip4(n9267), .op(n9269) );
  nor3_1 U10584 ( .ip1(n9363), .ip2(n9267), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[2]), .op(n9268) );
  not_ab_or_c_or_d U10585 ( .ip1(n9365), .ip2(n9364), .ip3(n9269), .ip4(n9268), 
        .op(n9270) );
  not_ab_or_c_or_d U10586 ( .ip1(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[4]), .ip2(n9371), .ip3(
        n9271), .ip4(n9270), .op(n9273) );
  nor3_1 U10587 ( .ip1(n9371), .ip2(n9271), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[4]), .op(n9272) );
  not_ab_or_c_or_d U10588 ( .ip1(n9374), .ip2(n9450), .ip3(n9273), .ip4(n9272), 
        .op(n9275) );
  not_ab_or_c_or_d U10589 ( .ip1(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[6]), .ip2(n9276), .ip3(
        n9275), .ip4(n9274), .op(n9277) );
  not_ab_or_c_or_d U10590 ( .ip1(n9379), .ip2(n9434), .ip3(n9278), .ip4(n9277), 
        .op(n9279) );
  ab_or_c_or_d U10591 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[8]), 
        .ip2(n9389), .ip3(n9286), .ip4(n9279), .op(n9285) );
  nor2_1 U10592 ( .ip1(n9396), .ip2(n9438), .op(n9284) );
  nor3_1 U10593 ( .ip1(n9291), .ip2(n9285), .ip3(n9284), .op(n9295) );
  nor3_1 U10594 ( .ip1(n9286), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[8]), .ip3(n9389), .op(
        n9287) );
  nor2_1 U10595 ( .ip1(n9382), .ip2(n9287), .op(n9289) );
  nor2_1 U10596 ( .ip1(n9383), .ip2(n9287), .op(n9288) );
  or2_1 U10597 ( .ip1(n9289), .ip2(n9288), .op(n9293) );
  nor2_1 U10598 ( .ip1(n9293), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[10]), .op(n9290) );
  nor2_1 U10599 ( .ip1(n9396), .ip2(n9290), .op(n9292) );
  not_ab_or_c_or_d U10600 ( .ip1(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[10]), .ip2(n9293), .ip3(
        n9292), .ip4(n9291), .op(n9294) );
  not_ab_or_c_or_d U10601 ( .ip1(n9398), .ip2(n9461), .ip3(n9295), .ip4(n9294), 
        .op(n9299) );
  nor2_1 U10602 ( .ip1(n9415), .ip2(n9463), .op(n9298) );
  nand2_1 U10603 ( .ip1(n9304), .ip2(i_i2c_ic_sda_tx_hold_sync[1]), .op(n9305)
         );
  nand2_1 U10604 ( .ip1(n9306), .ip2(n9305), .op(n9307) );
  nand2_1 U10605 ( .ip1(n9308), .ip2(n9307), .op(n9471) );
  nor3_1 U10606 ( .ip1(n9469), .ip2(n9341), .ip3(n9471), .op(
        i_i2c_U_DW_apb_i2c_tx_shift_mst_slv_ack_ext) );
  or2_1 U10607 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_stop_scl), .ip2(n9473), .op(
        n9310) );
  nand2_1 U10608 ( .ip1(n9310), .ip2(n9309), .op(n9311) );
  nand2_1 U10609 ( .ip1(n9311), .ip2(n11857), .op(n5043) );
  nor2_1 U10610 ( .ip1(i_i2c_mst_rx_data_scl), .ip2(n9312), .op(n9316) );
  nor2_1 U10611 ( .ip1(n9314), .ip2(n9313), .op(n9315) );
  nor2_1 U10612 ( .ip1(n9316), .ip2(n9315), .op(n4930) );
  nand2_1 U10613 ( .ip1(n9317), .ip2(i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl), 
        .op(n9318) );
  nand2_1 U10614 ( .ip1(n9319), .ip2(n9318), .op(n4954) );
  nand3_1 U10615 ( .ip1(n9321), .ip2(i_i2c_U_DW_apb_i2c_tx_shift_data_scl), 
        .ip3(n9320), .op(n9328) );
  nor2_1 U10616 ( .ip1(n9323), .ip2(n9322), .op(n9324) );
  or2_1 U10617 ( .ip1(n9325), .ip2(n9324), .op(n9326) );
  nand2_1 U10618 ( .ip1(n9326), .ip2(i_i2c_debug_wr), .op(n9327) );
  nand3_1 U10619 ( .ip1(n9328), .ip2(n11834), .ip3(n9327), .op(n4117) );
  nor3_1 U10620 ( .ip1(n11251), .ip2(n11253), .ip3(n11259), .op(n11264) );
  nand2_1 U10621 ( .ip1(n11264), .ip2(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[3]), .op(n11268) );
  nor2_1 U10622 ( .ip1(n11268), .ip2(n9329), .op(n11273) );
  nand2_1 U10623 ( .ip1(n11273), .ip2(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[5]), .op(n11284) );
  nor2_1 U10624 ( .ip1(n11284), .ip2(n11283), .op(n11277) );
  nand2_1 U10625 ( .ip1(n11277), .ip2(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[7]), .op(n9330) );
  nand2_1 U10626 ( .ip1(n9330), .ip2(n11272), .op(n11282) );
  nand2_1 U10627 ( .ip1(n11242), .ip2(i_i2c_slv_debug_cstate[3]), .op(n11239)
         );
  nor2_1 U10628 ( .ip1(n11083), .ip2(n11239), .op(n11056) );
  inv_1 U10629 ( .ip(n11056), .op(n10144) );
  nand3_1 U10630 ( .ip1(n11282), .ip2(n10144), .ip3(n9565), .op(
        i_i2c_scl_hld_low_en) );
  nor4_1 U10631 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_scl_hld_low_en_r), .ip2(
        i_i2c_scl_s_setup_en), .ip3(i_i2c_scl_p_setup_en), .ip4(
        i_i2c_U_DW_apb_i2c_tx_shift_data_scl_lcnt_en), .op(n9332) );
  nand2_1 U10632 ( .ip1(n9332), .ip2(n9331), .op(n9338) );
  nor4_1 U10633 ( .ip1(i_i2c_rx_scl_lcnt_en), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl_lcnt_en), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_stop_scl_lcnt_en), .ip4(i_i2c_start_en), 
        .op(n9334) );
  nand3_1 U10634 ( .ip1(n9335), .ip2(n9334), .ip3(n9333), .op(n9337) );
  nand4_1 U10635 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_stop_scl), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_data_scl), .ip3(i_i2c_mst_rx_data_scl), 
        .ip4(i_i2c_U_DW_apb_i2c_tx_shift_re_start_scl), .op(n9339) );
  nor2_1 U10636 ( .ip1(n9339), .ip2(i_i2c_scl_hld_low_en), .op(n9340) );
  nor3_1 U10637 ( .ip1(n9480), .ip2(n11096), .ip3(n9340), .op(n9346) );
  inv_1 U10638 ( .ip(n9471), .op(n9478) );
  not_ab_or_c_or_d U10639 ( .ip1(n9342), .ip2(n9478), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_mst_slv_ack_ext_r), .ip4(n9341), .op(n9481) );
  inv_1 U10640 ( .ip(n9480), .op(n9343) );
  not_ab_or_c_or_d U10641 ( .ip1(n11096), .ip2(n9481), .ip3(n9344), .ip4(n9343), .op(n9345) );
  or2_1 U10642 ( .ip1(n9346), .ip2(n9345), .op(n4951) );
  inv_1 U10643 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[2]), .op(
        n9426) );
  inv_1 U10644 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[0]), .op(
        n9443) );
  inv_1 U10645 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[15]), .op(
        n9347) );
  nor2_1 U10646 ( .ip1(n9347), .ip2(n9348), .op(n9352) );
  inv_1 U10647 ( .ip(n9402), .op(n9349) );
  and2_1 U10648 ( .ip1(n9350), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[14]), .op(n9351) );
  nor2_1 U10649 ( .ip1(n9352), .ip2(n9351), .op(n9423) );
  inv_1 U10650 ( .ip(n9383), .op(n9353) );
  inv_1 U10651 ( .ip(n9379), .op(n9378) );
  inv_1 U10652 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[5]), .op(
        n9450) );
  inv_1 U10653 ( .ip(n9368), .op(n9371) );
  nor2_1 U10654 ( .ip1(n9450), .ip2(n9374), .op(n9370) );
  inv_1 U10655 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[4]), .op(
        n9430) );
  inv_1 U10656 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[3]), .op(
        n9364) );
  nor2_1 U10657 ( .ip1(n9364), .ip2(n9365), .op(n9362) );
  nand2_1 U10658 ( .ip1(n9354), .ip2(n9443), .op(n9356) );
  inv_1 U10659 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[1]), .op(
        n9445) );
  nor2_1 U10660 ( .ip1(n9445), .ip2(n9357), .op(n9355) );
  nor2_1 U10661 ( .ip1(n9356), .ip2(n9355), .op(n9359) );
  and2_1 U10662 ( .ip1(n9357), .ip2(n9445), .op(n9358) );
  not_ab_or_c_or_d U10663 ( .ip1(n9426), .ip2(n9360), .ip3(n9358), .ip4(n9359), 
        .op(n9361) );
  not_ab_or_c_or_d U10664 ( .ip1(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[2]), .ip2(n9363), .ip3(
        n9362), .ip4(n9361), .op(n9367) );
  and2_1 U10665 ( .ip1(n9365), .ip2(n9364), .op(n9366) );
  not_ab_or_c_or_d U10666 ( .ip1(n9430), .ip2(n9368), .ip3(n9366), .ip4(n9367), 
        .op(n9369) );
  not_ab_or_c_or_d U10667 ( .ip1(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[4]), .ip2(n9371), .ip3(
        n9369), .ip4(n9370), .op(n9373) );
  inv_1 U10668 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[6]), .op(
        n9431) );
  not_ab_or_c_or_d U10669 ( .ip1(n9374), .ip2(n9450), .ip3(n9372), .ip4(n9373), 
        .op(n9377) );
  nor2_1 U10670 ( .ip1(n9431), .ip2(n9375), .op(n9376) );
  ab_or_c_or_d U10671 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[7]), 
        .ip2(n9378), .ip3(n9377), .ip4(n9376), .op(n9387) );
  inv_1 U10672 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[7]), .op(
        n9434) );
  nand2_1 U10673 ( .ip1(n9379), .ip2(n9434), .op(n9381) );
  inv_1 U10674 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[8]), .op(
        n9455) );
  nand2_1 U10675 ( .ip1(n9388), .ip2(n9455), .op(n9380) );
  nand2_1 U10676 ( .ip1(n9381), .ip2(n9380), .op(n9385) );
  inv_1 U10677 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[9]), .op(
        n9382) );
  nand2_1 U10678 ( .ip1(n9383), .ip2(n9382), .op(n9384) );
  nand2_1 U10679 ( .ip1(n9386), .ip2(n9387), .op(n9391) );
  inv_1 U10680 ( .ip(n9388), .op(n9389) );
  inv_1 U10681 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[10]), .op(
        n9438) );
  nand2_1 U10682 ( .ip1(n9396), .ip2(n9438), .op(n9394) );
  inv_1 U10683 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[11]), .op(
        n9461) );
  nand2_1 U10684 ( .ip1(n9398), .ip2(n9461), .op(n9393) );
  nand2_1 U10685 ( .ip1(n5519), .ip2(n5556), .op(n9397) );
  nand2_1 U10686 ( .ip1(n9397), .ip2(n9461), .op(n9401) );
  nand2_1 U10687 ( .ip1(n5524), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[10]), .op(n9399) );
  nand2_1 U10688 ( .ip1(n9399), .ip2(n9398), .op(n9400) );
  nand2_1 U10689 ( .ip1(n9400), .ip2(n9401), .op(n9411) );
  inv_1 U10690 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[14]), .op(
        n9466) );
  inv_1 U10691 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[13]), .op(
        n9441) );
  inv_1 U10692 ( .ip(n5557), .op(n9416) );
  nand2_1 U10693 ( .ip1(n9407), .ip2(n9441), .op(n9409) );
  nand2_1 U10694 ( .ip1(n5516), .ip2(n5523), .op(n9408) );
  nand2_1 U10695 ( .ip1(n9408), .ip2(n9409), .op(n9410) );
  and2_1 U10696 ( .ip1(n9411), .ip2(n9414), .op(n9412) );
  nand2_1 U10697 ( .ip1(n9413), .ip2(n9412), .op(n9421) );
  inv_1 U10698 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[12]), .op(
        n9463) );
  nand2_1 U10699 ( .ip1(n9415), .ip2(n9463), .op(n9417) );
  nand2_1 U10700 ( .ip1(n9420), .ip2(n9421), .op(n9422) );
  nand2_1 U10701 ( .ip1(n9444), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[1]), .op(n9425) );
  and2_1 U10702 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[2]), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[1]), .op(n9424) );
  inv_1 U10703 ( .ip(n9447), .op(n9427) );
  not_ab_or_c_or_d U10704 ( .ip1(n9426), .ip2(n9425), .ip3(n9469), .ip4(n9427), 
        .op(n4948) );
  nand2_1 U10705 ( .ip1(n9427), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[3]), .op(n9429) );
  nand2_1 U10706 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[4]), 
        .ip2(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[3]), .op(n9428) );
  not_ab_or_c_or_d U10707 ( .ip1(n9430), .ip2(n9429), .ip3(n9449), .ip4(n9469), 
        .op(n4946) );
  or2_1 U10708 ( .ip1(n9431), .ip2(n9452), .op(n9433) );
  nand2_1 U10709 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[6]), 
        .ip2(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[7]), .op(n9432) );
  not_ab_or_c_or_d U10710 ( .ip1(n9434), .ip2(n9433), .ip3(n9454), .ip4(n9469), 
        .op(n4943) );
  inv_1 U10711 ( .ip(n9458), .op(n9435) );
  nand2_1 U10712 ( .ip1(n9435), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[9]), .op(n9437) );
  nand2_1 U10713 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[9]), 
        .ip2(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[10]), .op(n9436) );
  not_ab_or_c_or_d U10714 ( .ip1(n9438), .ip2(n9437), .ip3(n9460), .ip4(n9469), 
        .op(n4940) );
  nand2_1 U10715 ( .ip1(n9462), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[12]), .op(n9440) );
  nand3_1 U10716 ( .ip1(n9462), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[13]), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[12]), .op(n9465) );
  inv_1 U10717 ( .ip(n9465), .op(n9439) );
  not_ab_or_c_or_d U10718 ( .ip1(n9441), .ip2(n9440), .ip3(n9469), .ip4(n9439), 
        .op(n4937) );
  not_ab_or_c_or_d U10719 ( .ip1(n9443), .ip2(n9442), .ip3(n9469), .ip4(n9444), 
        .op(n4950) );
  xor2_1 U10720 ( .ip1(n9445), .ip2(n9444), .op(n9446) );
  nor2_1 U10721 ( .ip1(n9469), .ip2(n9446), .op(n4949) );
  xor2_1 U10722 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[3]), .ip2(
        n9447), .op(n9448) );
  xor2_1 U10723 ( .ip1(n9450), .ip2(n9449), .op(n9451) );
  xnor2_1 U10724 ( .ip1(n9455), .ip2(n9454), .op(n9456) );
  inv_1 U10725 ( .ip(n9456), .op(n9457) );
  nor2_1 U10726 ( .ip1(n9469), .ip2(n9457), .op(n4942) );
  xor2_1 U10727 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[14]), 
        .ip2(n9465), .op(n9464) );
  nor2_1 U10728 ( .ip1(n9469), .ip2(n9464), .op(n4936) );
  nor2_1 U10729 ( .ip1(n9466), .ip2(n9465), .op(n9467) );
  nor2_1 U10730 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_sda_hold_count_r[15]), 
        .ip2(n9467), .op(n9468) );
  nor2_1 U10731 ( .ip1(n9469), .ip2(n9468), .op(n4935) );
  and3_1 U10732 ( .ip1(n9470), .ip2(i_i2c_U_DW_apb_i2c_tx_shift_slv_data_sda), 
        .ip3(i_i2c_U_DW_apb_i2c_tx_shift_data_sda), .op(n9472) );
  mux2_1 U10733 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_data_sda_prev_r), .ip2(
        n9472), .s(n9471), .op(n4934) );
  inv_1 U10734 ( .ip(i_i2c_U_DW_apb_i2c_tx_shift_stop_sda), .op(n9476) );
  mux2_1 U10735 ( .ip1(n9476), .ip2(n9474), .s(n9473), .op(n9475) );
  nand2_1 U10736 ( .ip1(n9475), .ip2(n11857), .op(n5042) );
  nand2_1 U10737 ( .ip1(n9478), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_stop_sda_gate_r), .op(n9477) );
  nand2_1 U10738 ( .ip1(n9477), .ip2(n9476), .op(
        i_i2c_U_DW_apb_i2c_tx_shift_N281) );
  nand2_1 U10739 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_start_sda_gate_r), .ip2(
        n9478), .op(n9482) );
  and3_1 U10740 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_re_start_sda_r), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_start_sda), .op(n9483) );
  or3_1 U10741 ( .ip1(i_i2c_ic_clk_oe), .ip2(n9483), .ip3(
        i_i2c_U_DW_apb_i2c_tx_shift_start_sda_gate_r), .op(n9479) );
  nand2_1 U10742 ( .ip1(n9482), .ip2(n9479), .op(
        i_i2c_U_DW_apb_i2c_tx_shift_N272) );
  nand2_1 U10743 ( .ip1(n9481), .ip2(n9480), .op(n9486) );
  and4_1 U10744 ( .ip1(n9483), .ip2(i_i2c_U_DW_apb_i2c_tx_shift_N281), .ip3(
        n9482), .ip4(n4934), .op(n9485) );
  nor2_1 U10745 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_ic_data_oe_early), .ip2(
        n9486), .op(n9484) );
  not_ab_or_c_or_d U10746 ( .ip1(n9486), .ip2(n9485), .ip3(n9484), .ip4(n11096), .op(i_i2c_U_DW_apb_i2c_tx_shift_N85) );
  and2_1 U10747 ( .ip1(n11045), .ip2(i_i2c_U_DW_apb_i2c_rx_filter_mst_arb_lost), .op(n9494) );
  nor4_1 U10748 ( .ip1(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[0]), 
        .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[3]), 
        .ip3(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[2]), 
        .ip4(
        i_i2c_U_DW_apb_i2c_rx_filter_delay_re_start_en_or_split_start_en[1]), 
        .op(n9487) );
  nand2_1 U10749 ( .ip1(n9487), .ip2(n11083), .op(n9492) );
  or2_1 U10750 ( .ip1(i_i2c_mst_tx_ack_vld), .ip2(n9488), .op(n9490) );
  nand2_1 U10751 ( .ip1(n11863), .ip2(i_i2c_mst_rx_ack_vld), .op(n9489) );
  xor2_1 U10752 ( .ip1(i_i2c_ic_data_oe), .ip2(n11833), .op(n9496) );
  ab_or_c_or_d U10753 ( .ip1(n9490), .ip2(n9489), .ip3(n11045), .ip4(n9496), 
        .op(n9491) );
  not_ab_or_c_or_d U10754 ( .ip1(n9492), .ip2(n9491), .ip3(i_i2c_start_en), 
        .ip4(n11857), .op(n9493) );
  nor2_1 U10755 ( .ip1(n9494), .ip2(n9493), .op(n9495) );
  nor2_1 U10756 ( .ip1(n11017), .ip2(n9495), .op(n4932) );
  inv_1 U10757 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_slv_arb_lost), .op(n9501) );
  nor3_1 U10758 ( .ip1(i_i2c_slv_tx_ack_vld), .ip2(n9497), .ip3(n9496), .op(
        n9498) );
  nor2_1 U10759 ( .ip1(n11045), .ip2(n9498), .op(n9500) );
  inv_1 U10760 ( .ip(i_i2c_slv_activity), .op(n9499) );
  not_ab_or_c_or_d U10761 ( .ip1(n9501), .ip2(n11045), .ip3(n9500), .ip4(n9499), .op(n4164) );
  nor2_1 U10762 ( .ip1(n9503), .ip2(n9502), .op(i_i2c_U_DW_apb_i2c_mstfsm_N73)
         );
  nand2_1 U10763 ( .ip1(n9505), .ip2(n9504), .op(n9512) );
  inv_1 U10764 ( .ip(n9512), .op(n9516) );
  nand2_1 U10765 ( .ip1(n9506), .ip2(n9516), .op(n9509) );
  nor2_1 U10766 ( .ip1(n9512), .ip2(n9507), .op(n9508) );
  not_ab_or_c_or_d U10767 ( .ip1(n9510), .ip2(n9509), .ip3(n11669), .ip4(n9508), .op(n5067) );
  nor2_1 U10768 ( .ip1(n9512), .ip2(n9511), .op(n9513) );
  nor2_1 U10769 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[7]), .ip2(
        n9513), .op(n9514) );
  not_ab_or_c_or_d U10770 ( .ip1(n9516), .ip2(n9515), .ip3(n11669), .ip4(n9514), .op(n5066) );
  nand2_1 U10771 ( .ip1(n9553), .ip2(i_i2c_rx_hs_mcode), .op(n9519) );
  nand2_1 U10772 ( .ip1(n9556), .ip2(n9517), .op(n9518) );
  nand2_1 U10773 ( .ip1(n9519), .ip2(n9518), .op(n5083) );
  inv_1 U10774 ( .ip(i_i2c_rx_hs_mcode), .op(n9520) );
  nand2_1 U10775 ( .ip1(n9520), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_rx_hs_mcode_r), .op(n9523) );
  inv_1 U10776 ( .ip(i_i2c_hs_mcode_en), .op(n9521) );
  nand2_1 U10777 ( .ip1(n9521), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_hs_mcode_en_r), .op(n9522) );
  mux2_1 U10778 ( .ip1(n9523), .ip2(n9522), .s(n11091), .op(n9524) );
  mux2_1 U10779 ( .ip1(n9524), .ip2(n11864), .s(
        i_i2c_U_DW_apb_i2c_rx_filter_hs_mcode_fed_dtctd_r), .op(n9525) );
  inv_1 U10780 ( .ip(n9525), .op(i_i2c_U_DW_apb_i2c_rx_filter_N50) );
  inv_1 U10781 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_hs_mcode_fed_dtctd_r), .op(
        n9526) );
  nor3_1 U10782 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv), .ip2(n9526), 
        .ip3(n11045), .op(n9527) );
  nor2_1 U10783 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_ic_hs_r), .ip2(n9527), 
        .op(n9528) );
  nor2_1 U10784 ( .ip1(n9528), .ip2(n11864), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_ic_hs) );
  mux2_1 U10785 ( .ip1(n9530), .ip2(i_i2c_U_DW_apb_i2c_rx_filter_scl_clk_int), 
        .s(n9529), .op(n5130) );
  inv_1 U10786 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt[0]), .op(n9531) );
  nor2_1 U10787 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt[1]), .ip2(n9531), 
        .op(n9532) );
  nor2_1 U10788 ( .ip1(n9532), .ip2(n9533), .op(n5087) );
  nor2_1 U10789 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt[0]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt[1]), .op(n9534) );
  nor2_1 U10790 ( .ip1(n9534), .ip2(n9533), .op(n5088) );
  inv_1 U10791 ( .ip(i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt[1]), .op(n9535) );
  nor2_1 U10792 ( .ip1(i_i2c_U_DW_apb_i2c_rx_filter_sda_cnt[0]), .ip2(n9535), 
        .op(n5227) );
  or2_1 U10793 ( .ip1(i_i2c_rx_slv_read), .ip2(n9544), .op(n9537) );
  nand2_1 U10794 ( .ip1(n9537), .ip2(n9536), .op(n9539) );
  nor2_1 U10795 ( .ip1(n9539), .ip2(n9538), .op(n9540) );
  nor2_1 U10796 ( .ip1(n11669), .ip2(n9540), .op(n9552) );
  inv_1 U10797 ( .ip(n9541), .op(n9542) );
  nand2_1 U10798 ( .ip1(n9543), .ip2(n9542), .op(n9545) );
  and2_1 U10799 ( .ip1(n9545), .ip2(n9544), .op(n11086) );
  nand2_1 U10800 ( .ip1(n11086), .ip2(n9546), .op(n9548) );
  inv_1 U10801 ( .ip(n11835), .op(n9547) );
  nand2_1 U10802 ( .ip1(n9548), .ip2(n9547), .op(n9549) );
  nand2_1 U10803 ( .ip1(n9549), .ip2(n9553), .op(n11087) );
  nor2_1 U10804 ( .ip1(n9550), .ip2(n11087), .op(n9551) );
  mux2_1 U10805 ( .ip1(n9552), .ip2(i_i2c_rx_addr_match), .s(n9551), .op(n5085) );
  inv_1 U10806 ( .ip(n9553), .op(n9559) );
  and3_1 U10807 ( .ip1(n9556), .ip2(n9555), .ip3(n9554), .op(n9557) );
  nor2_1 U10808 ( .ip1(i_i2c_rx_gen_call), .ip2(n9557), .op(n9558) );
  nor2_1 U10809 ( .ip1(n9559), .ip2(n9558), .op(n5084) );
  nand2_1 U10810 ( .ip1(n9560), .ip2(n11673), .op(n9561) );
  and2_1 U10811 ( .ip1(n11311), .ip2(n9561), .op(n9562) );
  nor2_1 U10812 ( .ip1(n10145), .ip2(n11239), .op(n9564) );
  or2_1 U10813 ( .ip1(n9564), .ip2(n11859), .op(n9586) );
  nand2_1 U10814 ( .ip1(n9586), .ip2(n9577), .op(n9570) );
  or2_1 U10815 ( .ip1(n9566), .ip2(n9565), .op(n9569) );
  nand2_1 U10816 ( .ip1(i_i2c_tx_fifo_data_buf[8]), .ip2(n11056), .op(n9568)
         );
  nand4_1 U10817 ( .ip1(n9570), .ip2(n9569), .ip3(n9568), .ip4(n9567), .op(
        n9571) );
  or2_1 U10818 ( .ip1(n10142), .ip2(n9571), .op(n11233) );
  inv_1 U10819 ( .ip(n11233), .op(n9581) );
  inv_1 U10820 ( .ip(i_i2c_rx_slv_read), .op(n11077) );
  and4_1 U10821 ( .ip1(i_i2c_rx_addr_match), .ip2(n11230), .ip3(
        i_i2c_U_DW_apb_i2c_sync_ic_10bit_slv_sync_inv), .ip4(n11077), .op(
        n9575) );
  inv_1 U10822 ( .ip(i_i2c_ic_ack_general_call_sync), .op(n9573) );
  inv_1 U10823 ( .ip(i_i2c_rx_gen_call), .op(n11671) );
  nor3_1 U10824 ( .ip1(n9573), .ip2(n9572), .ip3(n11671), .op(n9574) );
  nor2_1 U10825 ( .ip1(n9575), .ip2(n9574), .op(n9599) );
  nand3_1 U10826 ( .ip1(n11288), .ip2(i_i2c_slv_rxbyte_rdy), .ip3(
        i_i2c_rx_addr_match), .op(n9576) );
  nand2_1 U10827 ( .ip1(n9576), .ip2(n11296), .op(n9587) );
  nand2_1 U10828 ( .ip1(n9587), .ip2(n9577), .op(n9580) );
  inv_1 U10829 ( .ip(n9590), .op(n9578) );
  nand2_1 U10830 ( .ip1(n9578), .ip2(i_i2c_s_det), .op(n9579) );
  and4_1 U10831 ( .ip1(n9581), .ip2(n9599), .ip3(n9580), .ip4(n9579), .op(
        n9582) );
  nor2_1 U10832 ( .ip1(n11236), .ip2(n9582), .op(i_i2c_U_DW_apb_i2c_slvfsm_N38) );
  not_ab_or_c_or_d U10833 ( .ip1(n11279), .ip2(n9585), .ip3(n9584), .ip4(n9583), .op(n9588) );
  nor3_1 U10834 ( .ip1(n9588), .ip2(n9587), .ip3(n9586), .op(n9589) );
  nor2_1 U10835 ( .ip1(i_i2c_p_det), .ip2(n9589), .op(n9597) );
  inv_1 U10836 ( .ip(n11235), .op(n9591) );
  nor2_1 U10837 ( .ip1(n9591), .ip2(n9590), .op(n9596) );
  nand2_1 U10838 ( .ip1(i_i2c_ic_enable_sync), .ip2(i_i2c_s_det), .op(n9593)
         );
  not_ab_or_c_or_d U10839 ( .ip1(n9594), .ip2(n9593), .ip3(
        i_i2c_slv_debug_cstate[0]), .ip4(n9592), .op(n9595) );
  nor4_1 U10840 ( .ip1(n9598), .ip2(n9597), .ip3(n9596), .ip4(n9595), .op(
        n9600) );
  nand2_1 U10841 ( .ip1(n9600), .ip2(n9599), .op(n9602) );
  inv_1 U10842 ( .ip(n11236), .op(n9601) );
  inv_1 U10843 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[1]), .op(
        n11307) );
  inv_1 U10844 ( .ip(n9604), .op(n9606) );
  nand2_1 U10845 ( .ip1(n9604), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[1]), .op(n11667) );
  inv_1 U10846 ( .ip(n11667), .op(n9605) );
  not_ab_or_c_or_d U10847 ( .ip1(n11307), .ip2(n9606), .ip3(n11669), .ip4(
        n9605), .op(n4168) );
  inv_1 U10848 ( .ip(i_apb_U_DW_apb_ahbsif_nextstate[1]), .op(n10097) );
  nand2_1 U10849 ( .ip1(n9607), .ip2(n10097), .op(n9608) );
  mux2_1 U10850 ( .ip1(i_apb_psel_en), .ip2(n9608), .s(i_apb_pclk_en), .op(
        n4205) );
  nand2_1 U10851 ( .ip1(n9684), .ip2(i_apb_U_DW_apb_ahbsif_state[2]), .op(
        n10089) );
  nand2_1 U10852 ( .ip1(n10089), .ip2(n9609), .op(n9610) );
  mux2_1 U10853 ( .ip1(i_apb_penable), .ip2(n9610), .s(i_apb_pclk_en), .op(
        n4204) );
  nand2_1 U10854 ( .ip1(n9611), .ip2(i_apb_pwrite), .op(n9612) );
  nand2_1 U10855 ( .ip1(n11117), .ip2(n9612), .op(n4818) );
  mux2_1 U10856 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[12]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[12]), .s(n9690), .op(n4839) );
  nand2_1 U10857 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[12]), 
        .op(n9615) );
  nand2_1 U10858 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[12]), 
        .op(n9614) );
  nand2_1 U10859 ( .ip1(n9692), .ip2(i_apb_U_DW_apb_ahbsif_piped_haddr_c[12]), 
        .op(n9613) );
  nand3_1 U10860 ( .ip1(n9615), .ip2(n9614), .ip3(n9613), .op(n4746) );
  nand3_1 U10861 ( .ip1(n9616), .ip2(i_i2c_tx_fifo_data_buf[8]), .ip3(n11863), 
        .op(n9623) );
  nand3_1 U10862 ( .ip1(n9618), .ip2(n10941), .ip3(n9617), .op(n9622) );
  nand3_1 U10863 ( .ip1(n9620), .ip2(n11859), .ip3(n9619), .op(n9621) );
  nand3_1 U10864 ( .ip1(n9623), .ip2(n9622), .ip3(n9621), .op(
        i_i2c_U_DW_apb_i2c_tx_shift_N74) );
  xor2_1 U10865 ( .ip1(i_i2c_set_tx_empty_en), .ip2(i_i2c_set_tx_empty_en_flg), 
        .op(n4136) );
  xor2_1 U10866 ( .ip1(i_i2c_U_DW_apb_i2c_intctl_set_tx_empty_en_flg_sync_q), 
        .ip2(i_i2c_U_DW_apb_i2c_intctl_set_tx_empty_en_flg_sync), .op(n9629)
         );
  and2_1 U10867 ( .ip1(n9629), .ip2(i_i2c_tx_fifo_rst_n), .op(n9655) );
  xor2_1 U10868 ( .ip1(n9655), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[7]), .op(n9624) );
  xor2_1 U10869 ( .ip1(n9625), .ip2(n9624), .op(n9628) );
  nor2_1 U10870 ( .ip1(n11026), .ip2(n9626), .op(n9627) );
  or2_1 U10871 ( .ip1(n9655), .ip2(n9627), .op(n9657) );
  nand2_1 U10872 ( .ip1(n9628), .ip2(n9657), .op(n9631) );
  nor3_1 U10873 ( .ip1(n9629), .ip2(n11026), .ip3(i_i2c_tx_push), .op(n9658)
         );
  nand2_1 U10874 ( .ip1(n9658), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[7]), .op(n9630) );
  nand2_1 U10875 ( .ip1(n9631), .ip2(n9630), .op(n4128) );
  fulladder U10876 ( .a(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[6]), .b(n9655), .ci(n9632), .co(n9625), .s(n9633) );
  nand2_1 U10877 ( .ip1(n9633), .ip2(n9657), .op(n9635) );
  nand2_1 U10878 ( .ip1(n9658), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[6]), .op(n9634) );
  nand2_1 U10879 ( .ip1(n9635), .ip2(n9634), .op(n4129) );
  fulladder U10880 ( .a(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[5]), .b(n9655), .ci(n9636), .co(n9632), .s(n9637) );
  nand2_1 U10881 ( .ip1(n9637), .ip2(n9657), .op(n9639) );
  nand2_1 U10882 ( .ip1(n9658), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[5]), .op(n9638) );
  nand2_1 U10883 ( .ip1(n9639), .ip2(n9638), .op(n4130) );
  fulladder U10884 ( .a(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[4]), .b(n9655), .ci(n9640), .co(n9636), .s(n9641) );
  nand2_1 U10885 ( .ip1(n9641), .ip2(n9657), .op(n9643) );
  nand2_1 U10886 ( .ip1(n9658), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[4]), .op(n9642) );
  nand2_1 U10887 ( .ip1(n9643), .ip2(n9642), .op(n4131) );
  fulladder U10888 ( .a(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[3]), .b(n9655), .ci(n9644), .co(n9640), .s(n9645) );
  nand2_1 U10889 ( .ip1(n9645), .ip2(n9657), .op(n9647) );
  nand2_1 U10890 ( .ip1(n9658), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[3]), .op(n9646) );
  nand2_1 U10891 ( .ip1(n9647), .ip2(n9646), .op(n4132) );
  fulladder U10892 ( .a(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[2]), .b(n9655), .ci(n9648), .co(n9644), .s(n9649) );
  nand2_1 U10893 ( .ip1(n9649), .ip2(n9657), .op(n9651) );
  nand2_1 U10894 ( .ip1(n9658), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[2]), .op(n9650) );
  nand2_1 U10895 ( .ip1(n9651), .ip2(n9650), .op(n4133) );
  inv_1 U10896 ( .ip(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[0]), .op(n9652)
         );
  nand2_1 U10897 ( .ip1(n9657), .ip2(n9652), .op(n9654) );
  nand2_1 U10898 ( .ip1(n9658), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[0]), .op(n9653) );
  nand2_1 U10899 ( .ip1(n9654), .ip2(n9653), .op(n4135) );
  fulladder U10900 ( .a(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[1]), .b(n9655), .ci(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[0]), .co(n9648), .s(n9656) );
  nand2_1 U10901 ( .ip1(n9657), .ip2(n9656), .op(n9660) );
  nand2_1 U10902 ( .ip1(n9658), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[1]), .op(n9659) );
  nand2_1 U10903 ( .ip1(n9660), .ip2(n9659), .op(n4134) );
  inv_1 U10904 ( .ip(n11162), .op(n11160) );
  nor3_1 U10905 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[12]), .ip2(n9661), 
        .ip3(n11160), .op(ex_i_ahb_AHB_Slave_PWM_hsel) );
  mux2_1 U10906 ( .ip1(i_ahb_U_mux_hsel_prev[3]), .ip2(
        ex_i_ahb_AHB_Slave_PWM_hsel), .s(ex_i_ahb_AHB_MASTER_CORTEXM0_hready), 
        .op(n4851) );
  nand3_1 U10907 ( .ip1(n11162), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hready), 
        .ip3(n9661), .op(n9664) );
  nand2_1 U10908 ( .ip1(n9662), .ip2(i_ahb_U_mux_hsel_prev[2]), .op(n9663) );
  nand2_1 U10909 ( .ip1(n9664), .ip2(n9663), .op(n4850) );
  mux2_1 U10910 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[6]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[6]), .s(n9690), .op(n4841) );
  nand2_1 U10911 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[6]), 
        .op(n9667) );
  nand2_1 U10912 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[6]), 
        .op(n9666) );
  nand2_1 U10913 ( .ip1(n9692), .ip2(i_apb_U_DW_apb_ahbsif_piped_haddr_c[6]), 
        .op(n9665) );
  nand3_1 U10914 ( .ip1(n9667), .ip2(n9666), .ip3(n9665), .op(n4748) );
  mux2_1 U10915 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[7]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[7]), .s(n9690), .op(n4840) );
  nand2_1 U10916 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[7]), 
        .op(n9670) );
  nand2_1 U10917 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[7]), 
        .op(n9669) );
  nand2_1 U10918 ( .ip1(n9692), .ip2(i_apb_U_DW_apb_ahbsif_piped_haddr_c[7]), 
        .op(n9668) );
  nand3_1 U10919 ( .ip1(n9670), .ip2(n9669), .ip3(n9668), .op(n4747) );
  mux2_1 U10920 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[5]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[5]), .s(n9690), .op(n4842) );
  nand2_1 U10921 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[5]), 
        .op(n9673) );
  nand2_1 U10922 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[5]), 
        .op(n9672) );
  nand2_1 U10923 ( .ip1(n9692), .ip2(i_apb_U_DW_apb_ahbsif_piped_haddr_c[5]), 
        .op(n9671) );
  nand3_1 U10924 ( .ip1(n9673), .ip2(n9672), .ip3(n9671), .op(n4749) );
  mux2_1 U10925 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[3]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[3]), .s(n9690), .op(n4844) );
  nand2_1 U10926 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[3]), 
        .op(n9676) );
  nand2_1 U10927 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[3]), 
        .op(n9675) );
  nand2_1 U10928 ( .ip1(n9692), .ip2(i_apb_U_DW_apb_ahbsif_piped_haddr_c[3]), 
        .op(n9674) );
  nand3_1 U10929 ( .ip1(n9676), .ip2(n9675), .ip3(n9674), .op(n4751) );
  mux2_1 U10930 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[4]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[4]), .s(n9690), .op(n4843) );
  nand2_1 U10931 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[4]), 
        .op(n9679) );
  nand2_1 U10932 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[4]), 
        .op(n9678) );
  nand2_1 U10933 ( .ip1(n9692), .ip2(i_apb_U_DW_apb_ahbsif_piped_haddr_c[4]), 
        .op(n9677) );
  nand3_1 U10934 ( .ip1(n9679), .ip2(n9678), .ip3(n9677), .op(n4750) );
  inv_1 U10935 ( .ip(i_apb_U_DW_apb_ahbsif_use_saved_c), .op(n9680) );
  nor2_1 U10936 ( .ip1(n9680), .ip2(i_apb_pclk_en), .op(
        i_apb_U_DW_apb_ahbsif_N727) );
  nor2_1 U10937 ( .ip1(n9684), .ip2(n9681), .op(n9682) );
  or2_1 U10938 ( .ip1(i_apb_U_DW_apb_ahbsif_use_saved_data), .ip2(n9682), .op(
        n9683) );
  mux2_1 U10939 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[5]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[5]), .s(n11107), .op(n4810) );
  nand2_1 U10940 ( .ip1(n9684), .ip2(i_apb_U_DW_apb_ahbsif_use_saved_data), 
        .op(n9685) );
  nand2_1 U10941 ( .ip1(n5592), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[5]), .op(n9689) );
  nand2_1 U10942 ( .ip1(n9685), .ip2(n6858), .op(n9686) );
  nand2_1 U10943 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[5]), 
        .op(n9688) );
  nand2_1 U10944 ( .ip1(n11117), .ip2(i_apb_pwdata_int[5]), .op(n9687) );
  nand3_1 U10945 ( .ip1(n9689), .ip2(n9688), .ip3(n9687), .op(n4779) );
  mux2_1 U10946 ( .ip1(i_apb_U_DW_apb_ahbsif_piped_haddr_c[2]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[2]), .s(n9690), .op(n4845) );
  nand2_1 U10947 ( .ip1(n7201), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[2]), 
        .op(n9695) );
  nand2_1 U10948 ( .ip1(n9691), .ip2(i_apb_U_DW_apb_ahbsif_saved_haddr_c[2]), 
        .op(n9694) );
  nand2_1 U10949 ( .ip1(n9692), .ip2(i_apb_U_DW_apb_ahbsif_piped_haddr_c[2]), 
        .op(n9693) );
  nand3_1 U10950 ( .ip1(n9695), .ip2(n9694), .ip3(n9693), .op(n4752) );
  mux2_1 U10951 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[0]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[0]), .s(n11107), .op(n4815) );
  nand2_1 U10952 ( .ip1(n5592), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[0]), .op(n9698) );
  nand2_1 U10953 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[0]), 
        .op(n9697) );
  nand2_1 U10954 ( .ip1(n11117), .ip2(i_apb_pwdata_int[0]), .op(n9696) );
  nand3_1 U10955 ( .ip1(n9698), .ip2(n9697), .ip3(n9696), .op(n4784) );
  mux2_1 U10956 ( .ip1(n10802), .ip2(i_apb_pwdata_int[0]), .s(n9699), .op(
        n4631) );
  nor2_1 U10957 ( .ip1(n10802), .ip2(n10139), .op(n9811) );
  nand2_1 U10958 ( .ip1(n9811), .ip2(n11635), .op(n9746) );
  inv_1 U10959 ( .ip(n9700), .op(n9701) );
  nor2_1 U10960 ( .ip1(n9702), .ip2(n9701), .op(n4638) );
  or2_1 U10961 ( .ip1(n9988), .ip2(n10982), .op(n9703) );
  nand2_1 U10962 ( .ip1(n10802), .ip2(n9703), .op(i_ssi_U_mstfsm_N219) );
  mux2_1 U10963 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[1]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[1]), .s(n11107), .op(n4814) );
  nand2_1 U10964 ( .ip1(n5592), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[1]), .op(n9706) );
  nand2_1 U10965 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[1]), 
        .op(n9705) );
  nand2_1 U10966 ( .ip1(n11117), .ip2(i_apb_pwdata_int[1]), .op(n9704) );
  nand3_1 U10967 ( .ip1(n9706), .ip2(n9705), .ip3(n9704), .op(n4783) );
  mux2_1 U10968 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[2]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[2]), .s(n11107), .op(n4813) );
  nand2_1 U10969 ( .ip1(n5592), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[2]), .op(n9709) );
  nand2_1 U10970 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[2]), 
        .op(n9708) );
  nand2_1 U10971 ( .ip1(n11117), .ip2(i_apb_pwdata_int[2]), .op(n9707) );
  nand3_1 U10972 ( .ip1(n9709), .ip2(n9708), .ip3(n9707), .op(n4782) );
  mux2_1 U10973 ( .ip1(i_apb_pwdata_int[2]), .ip2(i_ssi_baudr[2]), .s(n9746), 
        .op(n4625) );
  mux2_1 U10974 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[3]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[3]), .s(n11107), .op(n4812) );
  nand2_1 U10975 ( .ip1(n5592), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[3]), .op(n9712) );
  nand2_1 U10976 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[3]), 
        .op(n9711) );
  nand2_1 U10977 ( .ip1(n11117), .ip2(i_apb_pwdata_int[3]), .op(n9710) );
  nand3_1 U10978 ( .ip1(n9712), .ip2(n9711), .ip3(n9710), .op(n4781) );
  mux2_1 U10979 ( .ip1(i_apb_pwdata_int[3]), .ip2(i_ssi_baudr[3]), .s(n9746), 
        .op(n4624) );
  mux2_1 U10980 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[4]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[4]), .s(n11107), .op(n4811) );
  nand2_1 U10981 ( .ip1(n5592), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[4]), .op(n9715) );
  nand2_1 U10982 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[4]), 
        .op(n9714) );
  nand2_1 U10983 ( .ip1(n11117), .ip2(i_apb_pwdata_int[4]), .op(n9713) );
  nand3_1 U10984 ( .ip1(n9715), .ip2(n9714), .ip3(n9713), .op(n4780) );
  mux2_1 U10985 ( .ip1(i_apb_pwdata_int[4]), .ip2(i_ssi_baudr[4]), .s(n9746), 
        .op(n4623) );
  mux2_1 U10986 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[15]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[15]), .s(n11107), .op(n4800) );
  nand2_1 U10987 ( .ip1(n5592), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[15]), .op(n9718) );
  nand2_1 U10988 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[15]), 
        .op(n9717) );
  nand2_1 U10989 ( .ip1(n11117), .ip2(i_apb_pwdata_int[15]), .op(n9716) );
  nand3_1 U10990 ( .ip1(n9718), .ip2(n9717), .ip3(n9716), .op(n4769) );
  mux2_1 U10991 ( .ip1(i_apb_pwdata_int[15]), .ip2(i_ssi_baudr[15]), .s(n9746), 
        .op(n4612) );
  mux2_1 U10992 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[14]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[14]), .s(n11107), .op(n4801) );
  nand2_1 U10993 ( .ip1(n5592), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[14]), .op(n9721) );
  nand2_1 U10994 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[14]), 
        .op(n9720) );
  nand2_1 U10995 ( .ip1(n11117), .ip2(i_apb_pwdata_int[14]), .op(n9719) );
  nand3_1 U10996 ( .ip1(n9721), .ip2(n9720), .ip3(n9719), .op(n4770) );
  mux2_1 U10997 ( .ip1(i_apb_pwdata_int[14]), .ip2(i_ssi_baudr[14]), .s(n9746), 
        .op(n4613) );
  mux2_1 U10998 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[13]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[13]), .s(n11107), .op(n4802) );
  nand2_1 U10999 ( .ip1(n5592), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[13]), .op(n9724) );
  nand2_1 U11000 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[13]), 
        .op(n9723) );
  nand2_1 U11001 ( .ip1(n11117), .ip2(i_apb_pwdata_int[13]), .op(n9722) );
  nand3_1 U11002 ( .ip1(n9724), .ip2(n9723), .ip3(n9722), .op(n4771) );
  mux2_1 U11003 ( .ip1(i_apb_pwdata_int[13]), .ip2(i_ssi_baudr[13]), .s(n9746), 
        .op(n4614) );
  mux2_1 U11004 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[12]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[12]), .s(n11107), .op(n4803) );
  nand2_1 U11005 ( .ip1(n5592), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[12]), .op(n9727) );
  nand2_1 U11006 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[12]), 
        .op(n9726) );
  nand2_1 U11007 ( .ip1(n11117), .ip2(i_apb_pwdata_int[12]), .op(n9725) );
  nand3_1 U11008 ( .ip1(n9727), .ip2(n9726), .ip3(n9725), .op(n4772) );
  mux2_1 U11009 ( .ip1(i_apb_pwdata_int[12]), .ip2(i_ssi_baudr[12]), .s(n9746), 
        .op(n4615) );
  mux2_1 U11010 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[11]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[11]), .s(n11107), .op(n4804) );
  nand2_1 U11011 ( .ip1(n5592), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[11]), .op(n9730) );
  nand2_1 U11012 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[11]), 
        .op(n9729) );
  nand2_1 U11013 ( .ip1(n11117), .ip2(i_apb_pwdata_int[11]), .op(n9728) );
  nand3_1 U11014 ( .ip1(n9730), .ip2(n9729), .ip3(n9728), .op(n4773) );
  mux2_1 U11015 ( .ip1(i_apb_pwdata_int[11]), .ip2(i_ssi_baudr[11]), .s(n9746), 
        .op(n4616) );
  mux2_1 U11016 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[10]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[10]), .s(n11107), .op(n4805) );
  nand2_1 U11017 ( .ip1(n5592), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[10]), .op(n9733) );
  nand2_1 U11018 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[10]), 
        .op(n9732) );
  nand2_1 U11019 ( .ip1(n11117), .ip2(i_apb_pwdata_int[10]), .op(n9731) );
  nand3_1 U11020 ( .ip1(n9733), .ip2(n9732), .ip3(n9731), .op(n4774) );
  mux2_1 U11021 ( .ip1(i_apb_pwdata_int[10]), .ip2(i_ssi_baudr[10]), .s(n9746), 
        .op(n4617) );
  mux2_1 U11022 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[9]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[9]), .s(n11107), .op(n4806) );
  nand2_1 U11023 ( .ip1(n5592), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[9]), .op(n9736) );
  nand2_1 U11024 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[9]), 
        .op(n9735) );
  nand2_1 U11025 ( .ip1(n11117), .ip2(i_apb_pwdata_int[9]), .op(n9734) );
  nand3_1 U11026 ( .ip1(n9736), .ip2(n9735), .ip3(n9734), .op(n4775) );
  mux2_1 U11027 ( .ip1(i_apb_pwdata_int[9]), .ip2(i_ssi_baudr[9]), .s(n9746), 
        .op(n4618) );
  mux2_1 U11028 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[8]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[8]), .s(n11107), .op(n4807) );
  nand2_1 U11029 ( .ip1(n5592), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[8]), .op(n9739) );
  nand2_1 U11030 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[8]), 
        .op(n9738) );
  nand2_1 U11031 ( .ip1(n11117), .ip2(i_apb_pwdata_int[8]), .op(n9737) );
  nand3_1 U11032 ( .ip1(n9739), .ip2(n9738), .ip3(n9737), .op(n4776) );
  mux2_1 U11033 ( .ip1(i_apb_pwdata_int[8]), .ip2(i_ssi_baudr[8]), .s(n9746), 
        .op(n4619) );
  mux2_1 U11034 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[7]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[7]), .s(n11107), .op(n4808) );
  nand2_1 U11035 ( .ip1(n5592), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[7]), .op(n9742) );
  nand2_1 U11036 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[7]), 
        .op(n9741) );
  nand2_1 U11037 ( .ip1(n11117), .ip2(i_apb_pwdata_int[7]), .op(n9740) );
  nand3_1 U11038 ( .ip1(n9742), .ip2(n9741), .ip3(n9740), .op(n4777) );
  mux2_1 U11039 ( .ip1(i_apb_pwdata_int[7]), .ip2(i_ssi_baudr[7]), .s(n9746), 
        .op(n4620) );
  mux2_1 U11040 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[6]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[6]), .s(n11107), .op(n4809) );
  nand2_1 U11041 ( .ip1(n5592), .ip2(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[6]), .op(n9745) );
  nand2_1 U11042 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[6]), 
        .op(n9744) );
  nand2_1 U11043 ( .ip1(n11117), .ip2(i_apb_pwdata_int[6]), .op(n9743) );
  nand3_1 U11044 ( .ip1(n9745), .ip2(n9744), .ip3(n9743), .op(n4778) );
  inv_1 U11045 ( .ip(n9747), .op(n9753) );
  or2_1 U11046 ( .ip1(i_ssi_baudr[10]), .ip2(i_ssi_baudr[14]), .op(n9751) );
  nor4_1 U11047 ( .ip1(i_ssi_baudr[13]), .ip2(i_ssi_baudr[8]), .ip3(
        i_ssi_baudr[11]), .ip4(i_ssi_baudr[12]), .op(n9749) );
  nor3_1 U11048 ( .ip1(i_ssi_baudr[5]), .ip2(i_ssi_baudr[15]), .ip3(
        i_ssi_baudr[9]), .op(n9748) );
  nand2_1 U11049 ( .ip1(n9749), .ip2(n9748), .op(n9750) );
  and2_1 U11050 ( .ip1(n10972), .ip2(i_ssi_baudr[1]), .op(n5234) );
  nand2_1 U11051 ( .ip1(n11855), .ip2(i_ssi_U_sclkgen_ssi_cnt[1]), .op(n9757)
         );
  or3_1 U11052 ( .ip1(n9755), .ip2(n9764), .ip3(i_ssi_U_sclkgen_ssi_cnt[1]), 
        .op(n9756) );
  nand2_1 U11053 ( .ip1(n9757), .ip2(n9756), .op(i_ssi_U_sclkgen_N41) );
  nand2_1 U11054 ( .ip1(n11855), .ip2(i_ssi_U_sclkgen_ssi_cnt[2]), .op(n9762)
         );
  nor2_1 U11055 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[2]), .ip2(n9764), .op(n9758) );
  mux2_1 U11056 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[2]), .ip2(n9758), .s(
        i_ssi_U_sclkgen_ssi_cnt[1]), .op(n9759) );
  nand2_1 U11057 ( .ip1(n9760), .ip2(n9759), .op(n9761) );
  nand2_1 U11058 ( .ip1(n9762), .ip2(n9761), .op(i_ssi_U_sclkgen_N42) );
  or2_1 U11059 ( .ip1(n9764), .ip2(n9763), .op(n9766) );
  inv_1 U11060 ( .ip(n5284), .op(n9785) );
  not_ab_or_c_or_d U11061 ( .ip1(n6419), .ip2(n9766), .ip3(n9765), .ip4(n5484), 
        .op(i_ssi_U_sclkgen_N43) );
  xor2_1 U11062 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[5]), .ip2(n9768), .op(n9767) );
  inv_1 U11063 ( .ip(n5284), .op(n9788) );
  nor2_1 U11064 ( .ip1(n9767), .ip2(n9785), .op(i_ssi_U_sclkgen_N45) );
  inv_1 U11065 ( .ip(i_ssi_U_sclkgen_ssi_cnt[6]), .op(n9772) );
  inv_1 U11066 ( .ip(n9768), .op(n9769) );
  nand2_1 U11067 ( .ip1(n9769), .ip2(i_ssi_U_sclkgen_ssi_cnt[5]), .op(n9771)
         );
  not_ab_or_c_or_d U11068 ( .ip1(n9772), .ip2(n9771), .ip3(n9770), .ip4(n9788), 
        .op(i_ssi_U_sclkgen_N46) );
  xor2_1 U11069 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[8]), .ip2(n9774), .op(n9773) );
  nor2_1 U11070 ( .ip1(n9773), .ip2(n9785), .op(i_ssi_U_sclkgen_N48) );
  inv_1 U11071 ( .ip(i_ssi_U_sclkgen_ssi_cnt[9]), .op(n9778) );
  inv_1 U11072 ( .ip(n9774), .op(n9775) );
  nand2_1 U11073 ( .ip1(n9775), .ip2(i_ssi_U_sclkgen_ssi_cnt[8]), .op(n9777)
         );
  not_ab_or_c_or_d U11074 ( .ip1(n9778), .ip2(n9777), .ip3(n9776), .ip4(n9785), 
        .op(i_ssi_U_sclkgen_N49) );
  xor2_1 U11075 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[11]), .ip2(n9780), .op(n9779)
         );
  nor2_1 U11076 ( .ip1(n9779), .ip2(n5484), .op(i_ssi_U_sclkgen_N51) );
  inv_1 U11077 ( .ip(n9780), .op(n9781) );
  nand2_1 U11078 ( .ip1(n9781), .ip2(i_ssi_U_sclkgen_ssi_cnt[11]), .op(n9782)
         );
  not_ab_or_c_or_d U11079 ( .ip1(n9783), .ip2(n9782), .ip3(n9787), .ip4(n9788), 
        .op(i_ssi_U_sclkgen_N52) );
  xor2_1 U11080 ( .ip1(n9784), .ip2(n9787), .op(n9786) );
  nor2_1 U11081 ( .ip1(n9786), .ip2(n5484), .op(i_ssi_U_sclkgen_N53) );
  nand2_1 U11082 ( .ip1(n9787), .ip2(i_ssi_U_sclkgen_ssi_cnt[13]), .op(n9790)
         );
  not_ab_or_c_or_d U11083 ( .ip1(n9791), .ip2(n9790), .ip3(n9789), .ip4(n9788), 
        .op(i_ssi_U_sclkgen_N54) );
  inv_1 U11084 ( .ip(n10139), .op(n9792) );
  nand3_1 U11085 ( .ip1(n9792), .ip2(n11469), .ip3(n11468), .op(n9793) );
  mux2_1 U11086 ( .ip1(i_apb_pwdata_int[0]), .ip2(i_ssi_ser_0_), .s(n9793), 
        .op(n4627) );
  nand2_1 U11087 ( .ip1(n9811), .ip2(n11592), .op(n11097) );
  mux2_1 U11088 ( .ip1(i_apb_pwdata_int[9]), .ip2(n5272), .s(n11097), .op(
        n4589) );
  or2_1 U11089 ( .ip1(n9794), .ip2(n9795), .op(n9796) );
  nor2_1 U11090 ( .ip1(n5291), .ip2(n9796), .op(i_ssi_U_sclkgen_N75) );
  mux2_1 U11091 ( .ip1(i_apb_pwdata_int[8]), .ip2(i_ssi_tmod[0]), .s(n11097), 
        .op(n4588) );
  nor2_1 U11092 ( .ip1(n10111), .ip2(n5399), .op(n9798) );
  nor2_1 U11093 ( .ip1(n9798), .ip2(n9797), .op(n9799) );
  nor2_1 U11094 ( .ip1(i_ssi_U_mstfsm_tx_load_en_int), .ip2(n9799), .op(n9801)
         );
  nor4_1 U11095 ( .ip1(n5400), .ip2(i_ssi_tmod[0]), .ip3(n10429), .ip4(n5288), 
        .op(n9800) );
  nor2_1 U11096 ( .ip1(n9801), .ip2(n9800), .op(n4579) );
  inv_1 U11097 ( .ip(n9972), .op(n9804) );
  nand2_1 U11098 ( .ip1(n9802), .ip2(n9974), .op(n9803) );
  nand2_1 U11099 ( .ip1(n9804), .ip2(n9803), .op(n9805) );
  nand2_1 U11100 ( .ip1(n9805), .ip2(n5290), .op(n9806) );
  nand2_1 U11101 ( .ip1(n9806), .ip2(i_ssi_U_mstfsm_last_frame), .op(n9809) );
  nand3_1 U11102 ( .ip1(n9815), .ip2(n9807), .ip3(n5492), .op(n9808) );
  nand2_1 U11103 ( .ip1(n9809), .ip2(n9808), .op(n4422) );
  nand2_1 U11104 ( .ip1(n9811), .ip2(n11636), .op(n9903) );
  mux2_1 U11105 ( .ip1(i_apb_pwdata_int[12]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[12]), .s(n9903), .op(n4607) );
  nor2_1 U11106 ( .ip1(n10136), .ip2(n9810), .op(n11548) );
  nand2_1 U11107 ( .ip1(n9811), .ip2(n11548), .op(n10836) );
  mux2_1 U11108 ( .ip1(i_apb_pwdata_int[0]), .ip2(i_ssi_mwcr[0]), .s(n10836), 
        .op(n4630) );
  inv_1 U11109 ( .ip(i_ssi_U_mstfsm_bit_cnt[0]), .op(n9826) );
  nand2_1 U11110 ( .ip1(n9812), .ip2(i_ssi_U_mstfsm_c_state[2]), .op(n9813) );
  or2_1 U11111 ( .ip1(n10112), .ip2(n9813), .op(n9825) );
  nor2_1 U11112 ( .ip1(n9826), .ip2(n9813), .op(n9814) );
  and2_1 U11113 ( .ip1(n9814), .ip2(n9975), .op(n9832) );
  nand2_1 U11114 ( .ip1(n9815), .ip2(i_ssi_mwcr[0]), .op(n9816) );
  nor2_1 U11115 ( .ip1(n9816), .ip2(n9853), .op(n9820) );
  nor2_1 U11116 ( .ip1(n10114), .ip2(n9817), .op(n9818) );
  nor2_1 U11117 ( .ip1(n10112), .ip2(n9818), .op(n9819) );
  nor2_1 U11118 ( .ip1(n9820), .ip2(n9819), .op(n9824) );
  nand3_1 U11119 ( .ip1(n10699), .ip2(i_ssi_U_mstfsm_c_state[1]), .ip3(
        i_ssi_sclk_fe), .op(n9822) );
  nand2_1 U11120 ( .ip1(n9972), .ip2(i_ssi_sclk_re), .op(n9821) );
  and2_1 U11121 ( .ip1(n9822), .ip2(n9821), .op(n9823) );
  nand2_1 U11122 ( .ip1(n9824), .ip2(n9823), .op(n10271) );
  not_ab_or_c_or_d U11123 ( .ip1(n9826), .ip2(n9825), .ip3(n9832), .ip4(n10271), .op(n4199) );
  xor2_1 U11124 ( .ip1(n9827), .ip2(n9832), .op(n9828) );
  nor2_1 U11125 ( .ip1(n9828), .ip2(n10271), .op(n4198) );
  not_ab_or_c_or_d U11126 ( .ip1(i_apb_pwdata_int[1]), .ip2(
        i_apb_pwdata_int[0]), .ip3(i_apb_pwdata_int[2]), .ip4(
        i_apb_pwdata_int[3]), .op(n9829) );
  nor2_1 U11127 ( .ip1(n9829), .ip2(n11097), .op(n9845) );
  mux2_1 U11128 ( .ip1(n5351), .ip2(i_apb_pwdata_int[1]), .s(n9845), .op(n4582) );
  inv_1 U11129 ( .ip(n9845), .op(n9839) );
  nand2_1 U11130 ( .ip1(n9839), .ip2(n5353), .op(n9831) );
  inv_1 U11131 ( .ip(n11097), .op(n10962) );
  nand2_1 U11132 ( .ip1(n10962), .ip2(i_apb_pwdata_int[2]), .op(n9830) );
  nand2_1 U11133 ( .ip1(n9831), .ip2(n9830), .op(n4583) );
  nand2_1 U11134 ( .ip1(n9832), .ip2(i_ssi_U_mstfsm_bit_cnt[1]), .op(n9835) );
  xor2_1 U11135 ( .ip1(i_ssi_U_mstfsm_bit_cnt[2]), .ip2(n9835), .op(n9833) );
  nor2_1 U11136 ( .ip1(n9833), .ip2(n10271), .op(n4197) );
  inv_1 U11137 ( .ip(n9835), .op(n9834) );
  nand2_1 U11138 ( .ip1(n9834), .ip2(i_ssi_U_mstfsm_bit_cnt[2]), .op(n9837) );
  nand2_1 U11139 ( .ip1(i_ssi_U_mstfsm_bit_cnt[3]), .ip2(
        i_ssi_U_mstfsm_bit_cnt[2]), .op(n9836) );
  nor2_1 U11140 ( .ip1(n9836), .ip2(n9835), .op(n9842) );
  not_ab_or_c_or_d U11141 ( .ip1(n9838), .ip2(n9837), .ip3(n9842), .ip4(n10271), .op(n4196) );
  nand2_1 U11142 ( .ip1(n9839), .ip2(n5453), .op(n9841) );
  nand2_1 U11143 ( .ip1(n10962), .ip2(i_apb_pwdata_int[3]), .op(n9840) );
  nand2_1 U11144 ( .ip1(n9841), .ip2(n9840), .op(n4584) );
  inv_1 U11145 ( .ip(i_ssi_U_mstfsm_bit_cnt[4]), .op(n9843) );
  xor2_1 U11146 ( .ip1(n9843), .ip2(n9842), .op(n9844) );
  nor2_1 U11147 ( .ip1(n10271), .ip2(n9844), .op(n4195) );
  mux2_1 U11148 ( .ip1(n5343), .ip2(i_apb_pwdata_int[0]), .s(n9845), .op(n4581) );
  nor2_1 U11149 ( .ip1(n9846), .ip2(n5396), .op(n9850) );
  nand2_1 U11150 ( .ip1(n9850), .ip2(n10420), .op(n9852) );
  nand2_1 U11151 ( .ip1(n10114), .ip2(n9851), .op(n10422) );
  nand2_1 U11152 ( .ip1(n10418), .ip2(i_ssi_sclk_fe), .op(n9856) );
  inv_1 U11153 ( .ip(n9853), .op(n10110) );
  nand2_1 U11154 ( .ip1(n10110), .ip2(n5501), .op(n9855) );
  and2_1 U11155 ( .ip1(n9856), .ip2(n9855), .op(n9857) );
  nand2_1 U11156 ( .ip1(n10377), .ip2(i_ssi_U_mstfsm_spi0_control), .op(n9858)
         );
  nand2_1 U11157 ( .ip1(n9858), .ip2(n5492), .op(n4193) );
  inv_1 U11158 ( .ip(n9879), .op(n9876) );
  inv_1 U11159 ( .ip(n11836), .op(n9910) );
  nand2_1 U11160 ( .ip1(n5479), .ip2(n9910), .op(n9872) );
  inv_1 U11161 ( .ip(n9872), .op(n9859) );
  mux2_1 U11162 ( .ip1(n9876), .ip2(n9859), .s(i_ssi_U_mstfsm_frame_cnt[0]), 
        .op(n4176) );
  nand2_1 U11163 ( .ip1(n9859), .ip2(i_ssi_U_mstfsm_frame_cnt[1]), .op(n9862)
         );
  xor2_1 U11164 ( .ip1(i_ssi_U_mstfsm_frame_cnt[1]), .ip2(
        i_ssi_U_mstfsm_frame_cnt[0]), .op(n9860) );
  nand2_1 U11165 ( .ip1(n9876), .ip2(n9860), .op(n9861) );
  nand2_1 U11166 ( .ip1(n9862), .ip2(n9861), .op(n4177) );
  inv_1 U11167 ( .ip(n9875), .op(n9863) );
  nand2_1 U11168 ( .ip1(n9876), .ip2(n9863), .op(n9864) );
  nand2_1 U11169 ( .ip1(n9864), .ip2(n9872), .op(n9868) );
  nand2_1 U11170 ( .ip1(n9868), .ip2(i_ssi_U_mstfsm_frame_cnt[2]), .op(n9867)
         );
  or2_1 U11171 ( .ip1(n9865), .ip2(n9864), .op(n9866) );
  nand2_1 U11172 ( .ip1(n9867), .ip2(n9866), .op(n4178) );
  nand2_1 U11173 ( .ip1(n9868), .ip2(i_ssi_U_mstfsm_frame_cnt[3]), .op(n9871)
         );
  nand3_1 U11174 ( .ip1(n9876), .ip2(n9875), .ip3(n9869), .op(n9870) );
  nand2_1 U11175 ( .ip1(n9871), .ip2(n9870), .op(n4179) );
  nand2_1 U11176 ( .ip1(n9876), .ip2(n9874), .op(n9873) );
  nand2_1 U11177 ( .ip1(n9873), .ip2(n9872), .op(n9880) );
  nand2_1 U11178 ( .ip1(n9880), .ip2(i_ssi_U_mstfsm_frame_cnt[4]), .op(n9878)
         );
  nand4_1 U11179 ( .ip1(n9876), .ip2(i_ssi_U_mstfsm_frame_cnt[3]), .ip3(n9875), 
        .ip4(n9874), .op(n9877) );
  nand2_1 U11180 ( .ip1(n9878), .ip2(n9877), .op(n4180) );
  mux2_1 U11181 ( .ip1(n5378), .ip2(n9880), .s(i_ssi_U_mstfsm_frame_cnt[5]), 
        .op(n4181) );
  and2_1 U11182 ( .ip1(n5378), .ip2(i_ssi_U_mstfsm_frame_cnt[5]), .op(n9882)
         );
  nor2_1 U11183 ( .ip1(n9886), .ip2(n5479), .op(n9881) );
  or2_1 U11184 ( .ip1(n9881), .ip2(n9880), .op(n9884) );
  mux2_1 U11185 ( .ip1(n9882), .ip2(n9884), .s(i_ssi_U_mstfsm_frame_cnt[6]), 
        .op(n4182) );
  inv_1 U11186 ( .ip(n9883), .op(n9885) );
  mux2_1 U11187 ( .ip1(n9885), .ip2(n9884), .s(i_ssi_U_mstfsm_frame_cnt[7]), 
        .op(n4183) );
  nand3_1 U11188 ( .ip1(n5378), .ip2(n9886), .ip3(i_ssi_U_mstfsm_frame_cnt[7]), 
        .op(n9887) );
  not_ab_or_c_or_d U11189 ( .ip1(n9888), .ip2(n9887), .ip3(n11836), .ip4(n9889), .op(n4184) );
  inv_1 U11190 ( .ip(n9889), .op(n9891) );
  inv_1 U11191 ( .ip(n9890), .op(n9893) );
  not_ab_or_c_or_d U11192 ( .ip1(n9892), .ip2(n9891), .ip3(n11836), .ip4(n9893), .op(n4185) );
  nand2_1 U11193 ( .ip1(n9893), .ip2(i_ssi_U_mstfsm_frame_cnt[10]), .op(n9894)
         );
  not_ab_or_c_or_d U11194 ( .ip1(n5390), .ip2(n9894), .ip3(n9895), .ip4(n11836), .op(n4187) );
  mux2_1 U11195 ( .ip1(i_apb_pwdata_int[13]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[13]), .s(n9903), .op(n4606) );
  nand2_1 U11196 ( .ip1(n9895), .ip2(i_ssi_U_mstfsm_frame_cnt[12]), .op(n9896)
         );
  not_ab_or_c_or_d U11197 ( .ip1(n9897), .ip2(n9896), .ip3(n11836), .ip4(n9898), .op(n4189) );
  mux2_1 U11198 ( .ip1(i_apb_pwdata_int[14]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[14]), .s(n9903), .op(n4605) );
  mux2_1 U11199 ( .ip1(i_apb_pwdata_int[15]), .ip2(n5434), .s(n9903), .op(
        n4604) );
  nand2_1 U11200 ( .ip1(n9898), .ip2(i_ssi_U_mstfsm_frame_cnt[14]), .op(n9901)
         );
  inv_1 U11201 ( .ip(n9899), .op(n9900) );
  not_ab_or_c_or_d U11202 ( .ip1(n9902), .ip2(n9901), .ip3(n11836), .ip4(n9900), .op(n4191) );
  mux2_1 U11203 ( .ip1(i_apb_pwdata_int[2]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[2]), .s(n9903), .op(n4601) );
  mux2_1 U11204 ( .ip1(i_apb_pwdata_int[1]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[1]), .s(n9903), .op(n4602) );
  mux2_1 U11205 ( .ip1(i_apb_pwdata_int[0]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[0]), .s(n9903), .op(n4603) );
  mux2_1 U11206 ( .ip1(i_apb_pwdata_int[4]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[4]), .s(n9903), .op(n4599) );
  mux2_1 U11207 ( .ip1(i_apb_pwdata_int[10]), .ip2(
        i_ssi_U_regfile_ctrlr1_int[10]), .s(n9903), .op(n4609) );
  inv_1 U11208 ( .ip(n5714), .op(n9905) );
  nor2_1 U11209 ( .ip1(n9905), .ip2(n9904), .op(n9906) );
  mux2_1 U11210 ( .ip1(i_ssi_U_mstfsm_last_frame), .ip2(n9906), .s(n5272), 
        .op(n9909) );
  inv_1 U11211 ( .ip(n9907), .op(n9908) );
  nand2_1 U11212 ( .ip1(n9909), .ip2(n9908), .op(n9912) );
  nand2_1 U11213 ( .ip1(n9910), .ip2(i_ssi_U_mstfsm_abort_ir), .op(n9911) );
  nand2_1 U11214 ( .ip1(n9912), .ip2(n9911), .op(n4421) );
  xor2_1 U11215 ( .ip1(i_ssi_tx_pop), .ip2(n5283), .op(n4578) );
  nand2_1 U11216 ( .ip1(n9926), .ip2(i_ssi_tx_full), .op(n9916) );
  inv_1 U11217 ( .ip(i_ssi_U_fifo_unconnected_tx_wrd_count[2]), .op(n9934) );
  nand2_1 U11218 ( .ip1(i_ssi_U_fifo_unconnected_tx_wrd_count[0]), .ip2(
        i_ssi_U_fifo_unconnected_tx_wrd_count[1]), .op(n9929) );
  nor2_1 U11219 ( .ip1(n9934), .ip2(n9929), .op(n9914) );
  nand2_1 U11220 ( .ip1(n10758), .ip2(n9914), .op(n9915) );
  nand2_1 U11221 ( .ip1(n9916), .ip2(n9915), .op(n10787) );
  and2_1 U11222 ( .ip1(n10787), .ip2(n10759), .op(n11873) );
  nand2_1 U11223 ( .ip1(n9921), .ip2(i_ssi_U_fifo_unconnected_tx_wrd_count[0]), 
        .op(n9932) );
  inv_1 U11224 ( .ip(i_ssi_U_fifo_unconnected_tx_wrd_count[0]), .op(n9919) );
  nand2_1 U11225 ( .ip1(n9926), .ip2(n9919), .op(n9917) );
  nand2_1 U11226 ( .ip1(n9932), .ip2(n9917), .op(n9918) );
  inv_1 U11227 ( .ip(i_ssi_U_fifo_unconnected_tx_wrd_count[1]), .op(n9927) );
  nand2_1 U11228 ( .ip1(n9918), .ip2(n9927), .op(n9925) );
  nand2_1 U11229 ( .ip1(n9919), .ip2(i_ssi_U_fifo_unconnected_tx_wrd_count[1]), 
        .op(n9920) );
  nor2_1 U11230 ( .ip1(n9920), .ip2(n9926), .op(n9923) );
  nor2_1 U11231 ( .ip1(n9929), .ip2(n9921), .op(n9922) );
  nor2_1 U11232 ( .ip1(n9923), .ip2(n9922), .op(n9924) );
  nand2_1 U11233 ( .ip1(n9925), .ip2(n9924), .op(n10795) );
  nor2_1 U11234 ( .ip1(n10748), .ip2(n10795), .op(n11872) );
  inv_1 U11235 ( .ip(n9926), .op(n9928) );
  nand2_1 U11236 ( .ip1(n9928), .ip2(n9927), .op(n9930) );
  nand2_1 U11237 ( .ip1(n9930), .ip2(n9929), .op(n9931) );
  nand2_1 U11238 ( .ip1(n9932), .ip2(n9931), .op(n9933) );
  xnor2_1 U11239 ( .ip1(n9934), .ip2(n9933), .op(n10791) );
  inv_1 U11240 ( .ip(n10791), .op(n9935) );
  and2_1 U11241 ( .ip1(n9935), .ip2(n10759), .op(n11852) );
  or2_1 U11242 ( .ip1(n11873), .ip2(n11872), .op(n10790) );
  inv_1 U11243 ( .ip(n10790), .op(n9937) );
  nor2_1 U11244 ( .ip1(n11853), .ip2(n11852), .op(n9936) );
  nand2_1 U11245 ( .ip1(n9937), .ip2(n9936), .op(i_ssi_U_fifo_U_tx_fifo_N33)
         );
  nor2_1 U11246 ( .ip1(i_ssi_U_regfile_txflr[0]), .ip2(
        i_ssi_U_regfile_txflr[1]), .op(n9945) );
  nor2_1 U11247 ( .ip1(i_ssi_U_regfile_txflr[2]), .ip2(
        i_ssi_U_regfile_txflr[3]), .op(n9968) );
  nand2_1 U11248 ( .ip1(n9945), .ip2(n9968), .op(n9938) );
  nand3_1 U11249 ( .ip1(n9938), .ip2(i_ssi_tx_pop_sync), .ip3(n10802), .op(
        n9939) );
  nor2_1 U11250 ( .ip1(n9939), .ip2(n11854), .op(n9962) );
  inv_1 U11251 ( .ip(i_ssi_U_regfile_txflr[0]), .op(n9965) );
  nand2_1 U11252 ( .ip1(n9962), .ip2(n9965), .op(n9942) );
  nor3_1 U11253 ( .ip1(i_ssi_U_regfile_txflr[3]), .ip2(n5291), .ip3(
        i_ssi_tx_pop_sync), .op(n9940) );
  nand2_1 U11254 ( .ip1(n11854), .ip2(n9940), .op(n9948) );
  nand2_1 U11255 ( .ip1(n9942), .ip2(n9941), .op(n9944) );
  inv_1 U11256 ( .ip(n9948), .op(n9961) );
  nand2_1 U11257 ( .ip1(n9961), .ip2(n9965), .op(n9943) );
  nand2_1 U11258 ( .ip1(n9944), .ip2(n9943), .op(n9951) );
  and2_1 U11259 ( .ip1(n9962), .ip2(n9945), .op(n9950) );
  inv_1 U11260 ( .ip(i_ssi_U_regfile_txflr[1]), .op(n9946) );
  nand2_1 U11261 ( .ip1(n9946), .ip2(i_ssi_U_regfile_txflr[0]), .op(n9966) );
  nor2_1 U11262 ( .ip1(n9966), .ip2(n9948), .op(n9947) );
  ab_or_c_or_d U11263 ( .ip1(n9951), .ip2(i_ssi_U_regfile_txflr[1]), .ip3(
        n9950), .ip4(n9947), .op(n4446) );
  nand2_1 U11264 ( .ip1(i_ssi_U_regfile_txflr[0]), .ip2(
        i_ssi_U_regfile_txflr[1]), .op(n9949) );
  nor2_1 U11265 ( .ip1(n9949), .ip2(n9948), .op(n9958) );
  nor2_1 U11266 ( .ip1(n9958), .ip2(n9950), .op(n9953) );
  mux2_1 U11267 ( .ip1(n9961), .ip2(n9962), .s(i_ssi_U_regfile_txflr[1]), .op(
        n9952) );
  nor2_1 U11268 ( .ip1(n9952), .ip2(n9951), .op(n9956) );
  mux2_1 U11269 ( .ip1(n9953), .ip2(n9956), .s(i_ssi_U_regfile_txflr[2]), .op(
        n9954) );
  inv_1 U11270 ( .ip(n9954), .op(n4445) );
  nand2_1 U11271 ( .ip1(n9962), .ip2(i_ssi_U_regfile_txflr[2]), .op(n9955) );
  nand2_1 U11272 ( .ip1(n9956), .ip2(n9955), .op(n9957) );
  nand2_1 U11273 ( .ip1(n9957), .ip2(i_ssi_U_regfile_txflr[3]), .op(n9960) );
  nand2_1 U11274 ( .ip1(n9958), .ip2(i_ssi_U_regfile_txflr[2]), .op(n9959) );
  nand2_1 U11275 ( .ip1(n9960), .ip2(n9959), .op(n4448) );
  nor2_1 U11276 ( .ip1(n9965), .ip2(n5291), .op(n9964) );
  nor2_1 U11277 ( .ip1(n9962), .ip2(n9961), .op(n9963) );
  mux2_1 U11278 ( .ip1(n9965), .ip2(n9964), .s(n9963), .op(n4447) );
  inv_1 U11279 ( .ip(n11854), .op(n9969) );
  inv_1 U11280 ( .ip(n9966), .op(n9967) );
  nand4_1 U11281 ( .ip1(i_ssi_tx_pop_sync), .ip2(n9969), .ip3(n9968), .ip4(
        n9967), .op(n9970) );
  and3_1 U11282 ( .ip1(n9970), .ip2(i_ssi_U_fifo_U_tx_fifo_empty_n), .ip3(
        i_ssi_ser_0_), .op(i_ssi_U_regfile_N452) );
  nand2_1 U11283 ( .ip1(i_ssi_U_mstfsm_ss_in_n_sync), .ip2(n10987), .op(n9971)
         );
  nand2_1 U11284 ( .ip1(n10802), .ip2(n9971), .op(i_ssi_U_mstfsm_N220) );
  mux2_1 U11285 ( .ip1(i_apb_pwdata_int[12]), .ip2(i_ssi_cfs[0]), .s(n11097), 
        .op(n4592) );
  and2_1 U11286 ( .ip1(n9972), .ip2(i_ssi_sclk_fe), .op(n10433) );
  nor2_1 U11287 ( .ip1(i_ssi_U_mstfsm_ctrl_cnt[0]), .ip2(n10433), .op(n9979)
         );
  nand3_1 U11288 ( .ip1(n10699), .ip2(i_ssi_U_mstfsm_c_state[1]), .ip3(
        i_ssi_sclk_re), .op(n9977) );
  nand3_1 U11289 ( .ip1(n9975), .ip2(n9974), .ip3(n9973), .op(n9976) );
  nand2_1 U11290 ( .ip1(n9977), .ip2(n9976), .op(n9987) );
  nand2_1 U11291 ( .ip1(n10433), .ip2(i_ssi_U_mstfsm_ctrl_cnt[0]), .op(n9980)
         );
  inv_1 U11292 ( .ip(n9980), .op(n9978) );
  nor3_1 U11293 ( .ip1(n9979), .ip2(n9987), .ip3(n9978), .op(n4203) );
  mux2_1 U11294 ( .ip1(i_apb_pwdata_int[13]), .ip2(i_ssi_cfs[1]), .s(n11097), 
        .op(n4593) );
  inv_1 U11295 ( .ip(i_ssi_U_mstfsm_ctrl_cnt[1]), .op(n9981) );
  nor2_1 U11296 ( .ip1(n9981), .ip2(n9980), .op(n9982) );
  not_ab_or_c_or_d U11297 ( .ip1(n9981), .ip2(n9980), .ip3(n9987), .ip4(n9982), 
        .op(n4202) );
  mux2_1 U11298 ( .ip1(i_apb_pwdata_int[15]), .ip2(i_ssi_cfs[3]), .s(n11097), 
        .op(n4595) );
  nor2_1 U11299 ( .ip1(i_ssi_U_mstfsm_ctrl_cnt[2]), .ip2(n9982), .op(n9984) );
  nand2_1 U11300 ( .ip1(n9982), .ip2(i_ssi_U_mstfsm_ctrl_cnt[2]), .op(n9985)
         );
  inv_1 U11301 ( .ip(n9985), .op(n9983) );
  nor3_1 U11302 ( .ip1(n9984), .ip2(n9987), .ip3(n9983), .op(n4201) );
  xor2_1 U11303 ( .ip1(i_ssi_U_mstfsm_ctrl_cnt[3]), .ip2(n9985), .op(n9986) );
  nor2_1 U11304 ( .ip1(n9987), .ip2(n9986), .op(n4200) );
  mux2_1 U11305 ( .ip1(i_apb_pwdata_int[14]), .ip2(i_ssi_cfs[2]), .s(n11097), 
        .op(n4594) );
  mux2_1 U11306 ( .ip1(i_apb_pwdata_int[1]), .ip2(i_ssi_mwcr[1]), .s(n10836), 
        .op(n4629) );
  inv_1 U11307 ( .ip(n10981), .op(n10951) );
  nor3_1 U11308 ( .ip1(n9988), .ip2(n5291), .ip3(n10951), .op(
        i_ssi_U_mstfsm_N221) );
  inv_1 U11309 ( .ip(n9989), .op(n10978) );
  nand2_1 U11310 ( .ip1(n10978), .ip2(i_ssi_U_mstfsm_ss_in_n_sync), .op(n9990)
         );
  nand2_1 U11311 ( .ip1(n9990), .ip2(n10802), .op(i_ssi_U_mstfsm_N222) );
  and2_1 U11312 ( .ip1(n9991), .ip2(i_ssi_risr[5]), .op(n9992) );
  nor2_1 U11313 ( .ip1(n10015), .ip2(n9992), .op(n9993) );
  nor2_1 U11314 ( .ip1(n5291), .ip2(n9993), .op(n4240) );
  nand2_1 U11315 ( .ip1(i_ssi_imr[5]), .ip2(i_ssi_risr[5]), .op(
        i_ssi_ssi_mst_intr_n) );
  inv_1 U11316 ( .ip(i_ssi_U_dff_rx_mem[37]), .op(n9994) );
  nor2_1 U11317 ( .ip1(n11616), .ip2(n9994), .op(n10000) );
  nand2_1 U11318 ( .ip1(n11618), .ip2(i_ssi_U_dff_rx_mem[69]), .op(n9998) );
  nand2_1 U11319 ( .ip1(n11614), .ip2(i_ssi_U_dff_rx_mem[53]), .op(n9997) );
  nand2_1 U11320 ( .ip1(n11628), .ip2(i_ssi_U_dff_rx_mem[85]), .op(n9996) );
  nand2_1 U11321 ( .ip1(n11619), .ip2(i_ssi_U_dff_rx_mem[101]), .op(n9995) );
  nand4_1 U11322 ( .ip1(n9998), .ip2(n9997), .ip3(n9996), .ip4(n9995), .op(
        n9999) );
  not_ab_or_c_or_d U11323 ( .ip1(i_ssi_U_dff_rx_mem[117]), .ip2(n11627), .ip3(
        n10000), .ip4(n9999), .op(n10003) );
  nand2_1 U11324 ( .ip1(n11620), .ip2(i_ssi_U_dff_rx_mem[5]), .op(n10002) );
  nand2_1 U11325 ( .ip1(n11617), .ip2(i_ssi_U_dff_rx_mem[21]), .op(n10001) );
  nand3_1 U11326 ( .ip1(n10003), .ip2(n10002), .ip3(n10001), .op(n10004) );
  nand2_1 U11327 ( .ip1(n10004), .ip2(n11632), .op(n10013) );
  inv_1 U11328 ( .ip(i_ssi_imr[5]), .op(n10006) );
  nor2_1 U11329 ( .ip1(n10006), .ip2(n10005), .op(n10007) );
  not_ab_or_c_or_d U11330 ( .ip1(n11636), .ip2(n5419), .ip3(n11661), .ip4(
        n10007), .op(n10012) );
  nor2_1 U11331 ( .ip1(n11484), .ip2(n11603), .op(n11641) );
  inv_1 U11332 ( .ip(n11635), .op(n11591) );
  nor2_1 U11333 ( .ip1(n10008), .ip2(n11591), .op(n10010) );
  nand2_1 U11334 ( .ip1(n11482), .ip2(n11468), .op(n11634) );
  nor2_1 U11335 ( .ip1(i_ssi_ssi_mst_intr_n), .ip2(n11634), .op(n10009) );
  not_ab_or_c_or_d U11336 ( .ip1(i_ssi_risr[5]), .ip2(n11641), .ip3(n10010), 
        .ip4(n10009), .op(n10011) );
  nand3_1 U11337 ( .ip1(n10013), .ip2(n10012), .ip3(n10011), .op(n10014) );
  mux2_1 U11338 ( .ip1(i_ssi_prdata[5]), .ip2(n10014), .s(n6687), .op(n4232)
         );
  inv_1 U11339 ( .ip(n10015), .op(n10018) );
  nand2_1 U11340 ( .ip1(n11647), .ip2(n6687), .op(n10016) );
  nand2_1 U11341 ( .ip1(i_ssi_U_regfile_sr_6_), .ip2(n10016), .op(n10017) );
  nand2_1 U11342 ( .ip1(n10018), .ip2(n10017), .op(n4238) );
  nand2_1 U11343 ( .ip1(n11628), .ip2(i_ssi_U_dff_rx_mem[88]), .op(n10028) );
  inv_1 U11344 ( .ip(i_ssi_U_dff_rx_mem[40]), .op(n10019) );
  nor2_1 U11345 ( .ip1(n11616), .ip2(n10019), .op(n10025) );
  nand2_1 U11346 ( .ip1(n11619), .ip2(i_ssi_U_dff_rx_mem[104]), .op(n10023) );
  nand2_1 U11347 ( .ip1(n11614), .ip2(i_ssi_U_dff_rx_mem[56]), .op(n10022) );
  nand2_1 U11348 ( .ip1(n11617), .ip2(i_ssi_U_dff_rx_mem[24]), .op(n10021) );
  nand2_1 U11349 ( .ip1(n11618), .ip2(i_ssi_U_dff_rx_mem[72]), .op(n10020) );
  nand4_1 U11350 ( .ip1(n10023), .ip2(n10022), .ip3(n10021), .ip4(n10020), 
        .op(n10024) );
  not_ab_or_c_or_d U11351 ( .ip1(i_ssi_U_dff_rx_mem[8]), .ip2(n11620), .ip3(
        n10025), .ip4(n10024), .op(n10027) );
  nand2_1 U11352 ( .ip1(n11627), .ip2(i_ssi_U_dff_rx_mem[120]), .op(n10026) );
  nand3_1 U11353 ( .ip1(n10028), .ip2(n10027), .ip3(n10026), .op(n10034) );
  inv_1 U11354 ( .ip(i_ssi_tmod[0]), .op(n10427) );
  nor2_1 U11355 ( .ip1(n10427), .ip2(n11470), .op(n10031) );
  nor2_1 U11356 ( .ip1(n10029), .ip2(n11591), .op(n10030) );
  ab_or_c_or_d U11357 ( .ip1(n11636), .ip2(i_ssi_U_regfile_ctrlr1_int[8]), 
        .ip3(n10031), .ip4(n10030), .op(n10032) );
  mux2_1 U11358 ( .ip1(i_ssi_prdata[8]), .ip2(n10032), .s(n6687), .op(n10033)
         );
  ab_or_c_or_d U11359 ( .ip1(n6937), .ip2(n10034), .ip3(n10081), .ip4(n10033), 
        .op(n4229) );
  nand2_1 U11360 ( .ip1(n11617), .ip2(i_ssi_U_dff_rx_mem[25]), .op(n10044) );
  inv_1 U11361 ( .ip(i_ssi_U_dff_rx_mem[41]), .op(n10035) );
  nor2_1 U11362 ( .ip1(n11616), .ip2(n10035), .op(n10041) );
  nand2_1 U11363 ( .ip1(n11618), .ip2(i_ssi_U_dff_rx_mem[73]), .op(n10039) );
  nand2_1 U11364 ( .ip1(n11628), .ip2(i_ssi_U_dff_rx_mem[89]), .op(n10038) );
  nand2_1 U11365 ( .ip1(n11614), .ip2(i_ssi_U_dff_rx_mem[57]), .op(n10037) );
  nand2_1 U11366 ( .ip1(n11620), .ip2(i_ssi_U_dff_rx_mem[9]), .op(n10036) );
  nand4_1 U11367 ( .ip1(n10039), .ip2(n10038), .ip3(n10037), .ip4(n10036), 
        .op(n10040) );
  not_ab_or_c_or_d U11368 ( .ip1(i_ssi_U_dff_rx_mem[105]), .ip2(n11619), .ip3(
        n10041), .ip4(n10040), .op(n10043) );
  nand2_1 U11369 ( .ip1(n11627), .ip2(i_ssi_U_dff_rx_mem[121]), .op(n10042) );
  nand3_1 U11370 ( .ip1(n10044), .ip2(n10043), .ip3(n10042), .op(n10050) );
  nand2_1 U11371 ( .ip1(n11592), .ip2(n5272), .op(n10047) );
  nand2_1 U11372 ( .ip1(n11636), .ip2(n5383), .op(n10046) );
  nand2_1 U11373 ( .ip1(n11635), .ip2(i_ssi_baudr[9]), .op(n10045) );
  nand3_1 U11374 ( .ip1(n10047), .ip2(n10046), .ip3(n10045), .op(n10048) );
  mux2_1 U11375 ( .ip1(i_ssi_prdata[9]), .ip2(n10048), .s(n6687), .op(n10049)
         );
  ab_or_c_or_d U11376 ( .ip1(n6937), .ip2(n10050), .ip3(n10081), .ip4(n10049), 
        .op(n4228) );
  nand2_1 U11377 ( .ip1(n11618), .ip2(i_ssi_U_dff_rx_mem[76]), .op(n10060) );
  inv_1 U11378 ( .ip(i_ssi_U_dff_rx_mem[44]), .op(n10051) );
  nor2_1 U11379 ( .ip1(n11616), .ip2(n10051), .op(n10057) );
  nand2_1 U11380 ( .ip1(n11620), .ip2(i_ssi_U_dff_rx_mem[12]), .op(n10055) );
  nand2_1 U11381 ( .ip1(n11619), .ip2(i_ssi_U_dff_rx_mem[108]), .op(n10054) );
  nand2_1 U11382 ( .ip1(n11628), .ip2(i_ssi_U_dff_rx_mem[92]), .op(n10053) );
  nand2_1 U11383 ( .ip1(n11617), .ip2(i_ssi_U_dff_rx_mem[28]), .op(n10052) );
  nand4_1 U11384 ( .ip1(n10055), .ip2(n10054), .ip3(n10053), .ip4(n10052), 
        .op(n10056) );
  not_ab_or_c_or_d U11385 ( .ip1(i_ssi_U_dff_rx_mem[124]), .ip2(n11627), .ip3(
        n10057), .ip4(n10056), .op(n10059) );
  nand2_1 U11386 ( .ip1(n11614), .ip2(i_ssi_U_dff_rx_mem[60]), .op(n10058) );
  nand3_1 U11387 ( .ip1(n10060), .ip2(n10059), .ip3(n10058), .op(n10066) );
  nor2_1 U11388 ( .ip1(n10437), .ip2(n11470), .op(n10063) );
  inv_1 U11389 ( .ip(i_ssi_baudr[12]), .op(n10061) );
  nor2_1 U11390 ( .ip1(n10061), .ip2(n11591), .op(n10062) );
  ab_or_c_or_d U11391 ( .ip1(n11636), .ip2(i_ssi_U_regfile_ctrlr1_int[12]), 
        .ip3(n10063), .ip4(n10062), .op(n10064) );
  mux2_1 U11392 ( .ip1(i_ssi_prdata[12]), .ip2(n10064), .s(n6687), .op(n10065)
         );
  ab_or_c_or_d U11393 ( .ip1(n6937), .ip2(n10066), .ip3(n10081), .ip4(n10065), 
        .op(n4225) );
  nand2_1 U11394 ( .ip1(n11628), .ip2(i_ssi_U_dff_rx_mem[93]), .op(n10076) );
  inv_1 U11395 ( .ip(i_ssi_U_dff_rx_mem[45]), .op(n10067) );
  nor2_1 U11396 ( .ip1(n11616), .ip2(n10067), .op(n10073) );
  nand2_1 U11397 ( .ip1(n11617), .ip2(i_ssi_U_dff_rx_mem[29]), .op(n10071) );
  nand2_1 U11398 ( .ip1(n11614), .ip2(i_ssi_U_dff_rx_mem[61]), .op(n10070) );
  nand2_1 U11399 ( .ip1(n11619), .ip2(i_ssi_U_dff_rx_mem[109]), .op(n10069) );
  nand2_1 U11400 ( .ip1(n11620), .ip2(i_ssi_U_dff_rx_mem[13]), .op(n10068) );
  nand4_1 U11401 ( .ip1(n10071), .ip2(n10070), .ip3(n10069), .ip4(n10068), 
        .op(n10072) );
  not_ab_or_c_or_d U11402 ( .ip1(i_ssi_U_dff_rx_mem[77]), .ip2(n11618), .ip3(
        n10073), .ip4(n10072), .op(n10075) );
  nand2_1 U11403 ( .ip1(n11627), .ip2(i_ssi_U_dff_rx_mem[125]), .op(n10074) );
  nand3_1 U11404 ( .ip1(n10076), .ip2(n10075), .ip3(n10074), .op(n10082) );
  nor2_1 U11405 ( .ip1(n10438), .ip2(n11470), .op(n10078) );
  nor2_1 U11406 ( .ip1(n6389), .ip2(n11591), .op(n10077) );
  ab_or_c_or_d U11407 ( .ip1(n11636), .ip2(i_ssi_U_regfile_ctrlr1_int[13]), 
        .ip3(n10078), .ip4(n10077), .op(n10079) );
  mux2_1 U11408 ( .ip1(i_ssi_prdata[13]), .ip2(n10079), .s(n6687), .op(n10080)
         );
  ab_or_c_or_d U11409 ( .ip1(n6937), .ip2(n10082), .ip3(n10081), .ip4(n10080), 
        .op(n4224) );
  nand2_1 U11410 ( .ip1(n10084), .ip2(n10083), .op(n10086) );
  nand2_1 U11411 ( .ip1(n10086), .ip2(n10085), .op(n10088) );
  nand2_1 U11412 ( .ip1(n10088), .ip2(n10087), .op(n10090) );
  nand2_1 U11413 ( .ip1(n10090), .ip2(n10089), .op(n10109) );
  not_ab_or_c_or_d U11414 ( .ip1(n10094), .ip2(n10093), .ip3(n10092), .ip4(
        n10091), .op(n10107) );
  nor3_1 U11415 ( .ip1(n10097), .ip2(n10096), .ip3(n10095), .op(n10104) );
  not_ab_or_c_or_d U11416 ( .ip1(n10101), .ip2(n10100), .ip3(n10099), .ip4(
        n10098), .op(n10102) );
  or4_1 U11417 ( .ip1(n10105), .ip2(n10104), .ip3(n10103), .ip4(n10102), .op(
        n10106) );
  nor2_1 U11418 ( .ip1(n10107), .ip2(n10106), .op(n10108) );
  mux2_1 U11419 ( .ip1(n10109), .ip2(i_apb_hready_resp), .s(n10108), .op(n4817) );
  mux2_1 U11420 ( .ip1(i_apb_pwdata_int[11]), .ip2(i_ssi_ctrlr0[11]), .s(
        n11097), .op(n4591) );
  nand2_1 U11421 ( .ip1(n10110), .ip2(i_ssi_ctrlr0[11]), .op(n10116) );
  nand2_1 U11422 ( .ip1(n10112), .ip2(n10111), .op(n10113) );
  nand2_1 U11423 ( .ip1(n10114), .ip2(n10113), .op(n10115) );
  nand2_1 U11424 ( .ip1(n10116), .ip2(n10115), .op(n10121) );
  inv_1 U11425 ( .ip(i_ssi_U_mstfsm_spi0_control), .op(n10117) );
  nand2_1 U11426 ( .ip1(n10117), .ip2(n5272), .op(n10119) );
  not_ab_or_c_or_d U11427 ( .ip1(i_ssi_tmod[0]), .ip2(n10119), .ip3(n5291), 
        .ip4(n10118), .op(n10120) );
  and2_1 U11428 ( .ip1(n10121), .ip2(n10120), .op(n10122) );
  xor2_1 U11429 ( .ip1(i_ssi_rx_push), .ip2(n10122), .op(n4444) );
  nor2_1 U11430 ( .ip1(n10748), .ip2(n10123), .op(n11869) );
  and2_1 U11431 ( .ip1(n10124), .ip2(n10759), .op(n11870) );
  nor3_1 U11432 ( .ip1(n11871), .ip2(n11869), .ip3(n11850), .op(n10126) );
  inv_1 U11433 ( .ip(n11870), .op(n10125) );
  nand2_1 U11434 ( .ip1(n10126), .ip2(n10125), .op(i_ssi_U_fifo_U_rx_fifo_N33)
         );
  nor2_1 U11435 ( .ip1(n10127), .ip2(n10128), .op(n10132) );
  not_ab_or_c_or_d U11436 ( .ip1(n10128), .ip2(n10127), .ip3(n10132), .ip4(
        n10133), .op(n11849) );
  inv_1 U11437 ( .ip(n11849), .op(n10129) );
  nor2_1 U11438 ( .ip1(n10130), .ip2(n10129), .op(i_ssi_U_fifo_U_rx_fifo_N39)
         );
  inv_1 U11439 ( .ip(n10131), .op(n10135) );
  nor2_1 U11440 ( .ip1(i_ssi_rx_rd_addr[1]), .ip2(n10132), .op(n10134) );
  nor3_1 U11441 ( .ip1(n10135), .ip2(n10134), .ip3(n10133), .op(
        i_ssi_U_fifo_U_rx_fifo_N45) );
  inv_1 U11442 ( .ip(n10136), .op(n10137) );
  inv_1 U11443 ( .ip(n11463), .op(n10785) );
  nand2_1 U11444 ( .ip1(n10137), .ip2(n10785), .op(n11529) );
  inv_1 U11445 ( .ip(n11529), .op(n11546) );
  or3_1 U11446 ( .ip1(i_apb_pwdata_int[3]), .ip2(i_apb_pwdata_int[5]), .ip3(
        i_apb_pwdata_int[7]), .op(n10138) );
  nor4_1 U11447 ( .ip1(i_apb_pwdata_int[4]), .ip2(i_apb_pwdata_int[6]), .ip3(
        n10139), .ip4(n10138), .op(n10786) );
  nand2_1 U11448 ( .ip1(n11546), .ip2(n10786), .op(n10835) );
  mux2_1 U11449 ( .ip1(i_apb_pwdata_int[0]), .ip2(i_ssi_rxftlr[0]), .s(n10835), 
        .op(n4637) );
  mux2_1 U11450 ( .ip1(i_apb_pwdata_int[1]), .ip2(i_ssi_rxftlr[1]), .s(n10835), 
        .op(n4636) );
  inv_1 U11451 ( .ip(n10140), .op(n10141) );
  nor2_1 U11452 ( .ip1(i_i2c_slv_ack_det), .ip2(n10141), .op(n11315) );
  or2_1 U11453 ( .ip1(n10142), .ip2(n11315), .op(n10143) );
  and2_1 U11454 ( .ip1(i_i2c_U_DW_apb_i2c_sync_tx_empty_int_inv), .ip2(n10143), 
        .op(n11314) );
  nand2_1 U11455 ( .ip1(n10144), .ip2(n11057), .op(n11293) );
  and2_1 U11456 ( .ip1(n11293), .ip2(n10145), .op(n10146) );
  nor2_1 U11457 ( .ip1(n11314), .ip2(n10146), .op(n11240) );
  nand2_1 U11458 ( .ip1(n10147), .ip2(n11240), .op(
        i_i2c_U_DW_apb_i2c_toggle_tx_abrt) );
  nand2_1 U11459 ( .ip1(i_i2c_U_dff_tx_mem[49]), .ip2(n10178), .op(n10156) );
  and2_1 U11460 ( .ip1(n11214), .ip2(i_i2c_U_dff_tx_mem[4]), .op(n10153) );
  nand2_1 U11461 ( .ip1(n10180), .ip2(i_i2c_U_dff_tx_mem[31]), .op(n10151) );
  nand2_1 U11462 ( .ip1(n10179), .ip2(i_i2c_U_dff_tx_mem[22]), .op(n10150) );
  nand2_1 U11463 ( .ip1(n10190), .ip2(i_i2c_U_dff_tx_mem[40]), .op(n10149) );
  nand2_1 U11464 ( .ip1(n10182), .ip2(i_i2c_U_dff_tx_mem[67]), .op(n10148) );
  nand4_1 U11465 ( .ip1(n10151), .ip2(n10150), .ip3(n10149), .ip4(n10148), 
        .op(n10152) );
  not_ab_or_c_or_d U11466 ( .ip1(n10181), .ip2(i_i2c_U_dff_tx_mem[58]), .ip3(
        n10153), .ip4(n10152), .op(n10155) );
  nand2_1 U11467 ( .ip1(n10189), .ip2(i_i2c_U_dff_tx_mem[13]), .op(n10154) );
  nand3_1 U11468 ( .ip1(n10156), .ip2(n10155), .ip3(n10154), .op(n10157) );
  mux2_1 U11469 ( .ip1(i_i2c_tx_fifo_data_buf[4]), .ip2(n10157), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .op(n5218) );
  nand2_1 U11470 ( .ip1(i_i2c_U_dff_tx_mem[60]), .ip2(n10181), .op(n10166) );
  and2_1 U11471 ( .ip1(n11214), .ip2(i_i2c_U_dff_tx_mem[6]), .op(n10163) );
  nand2_1 U11472 ( .ip1(n10182), .ip2(i_i2c_U_dff_tx_mem[69]), .op(n10161) );
  nand2_1 U11473 ( .ip1(n10190), .ip2(i_i2c_U_dff_tx_mem[42]), .op(n10160) );
  nand2_1 U11474 ( .ip1(n10179), .ip2(i_i2c_U_dff_tx_mem[24]), .op(n10159) );
  nand2_1 U11475 ( .ip1(n10189), .ip2(i_i2c_U_dff_tx_mem[15]), .op(n10158) );
  nand4_1 U11476 ( .ip1(n10161), .ip2(n10160), .ip3(n10159), .ip4(n10158), 
        .op(n10162) );
  not_ab_or_c_or_d U11477 ( .ip1(n10178), .ip2(i_i2c_U_dff_tx_mem[51]), .ip3(
        n10163), .ip4(n10162), .op(n10165) );
  nand2_1 U11478 ( .ip1(n10180), .ip2(i_i2c_U_dff_tx_mem[33]), .op(n10164) );
  nand3_1 U11479 ( .ip1(n10166), .ip2(n10165), .ip3(n10164), .op(n10167) );
  mux2_1 U11480 ( .ip1(i_i2c_tx_fifo_data_buf[6]), .ip2(n10167), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .op(n5216) );
  nand2_1 U11481 ( .ip1(i_i2c_U_dff_tx_mem[59]), .ip2(n10181), .op(n10176) );
  and2_1 U11482 ( .ip1(n11214), .ip2(i_i2c_U_dff_tx_mem[5]), .op(n10173) );
  nand2_1 U11483 ( .ip1(n10190), .ip2(i_i2c_U_dff_tx_mem[41]), .op(n10171) );
  nand2_1 U11484 ( .ip1(n10179), .ip2(i_i2c_U_dff_tx_mem[23]), .op(n10170) );
  nand2_1 U11485 ( .ip1(n10180), .ip2(i_i2c_U_dff_tx_mem[32]), .op(n10169) );
  nand2_1 U11486 ( .ip1(n10189), .ip2(i_i2c_U_dff_tx_mem[14]), .op(n10168) );
  nand4_1 U11487 ( .ip1(n10171), .ip2(n10170), .ip3(n10169), .ip4(n10168), 
        .op(n10172) );
  not_ab_or_c_or_d U11488 ( .ip1(i_i2c_U_dff_tx_mem[68]), .ip2(n10182), .ip3(
        n10173), .ip4(n10172), .op(n10175) );
  nand2_1 U11489 ( .ip1(n10178), .ip2(i_i2c_U_dff_tx_mem[50]), .op(n10174) );
  nand3_1 U11490 ( .ip1(n10176), .ip2(n10175), .ip3(n10174), .op(n10177) );
  mux2_1 U11491 ( .ip1(i_i2c_tx_fifo_data_buf[5]), .ip2(n10177), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .op(n5217) );
  nand2_1 U11492 ( .ip1(n10178), .ip2(i_i2c_U_dff_tx_mem[48]), .op(n10193) );
  and2_1 U11493 ( .ip1(n11214), .ip2(i_i2c_U_dff_tx_mem[3]), .op(n10188) );
  nand2_1 U11494 ( .ip1(n10179), .ip2(i_i2c_U_dff_tx_mem[21]), .op(n10186) );
  nand2_1 U11495 ( .ip1(n10180), .ip2(i_i2c_U_dff_tx_mem[30]), .op(n10185) );
  nand2_1 U11496 ( .ip1(n10181), .ip2(i_i2c_U_dff_tx_mem[57]), .op(n10184) );
  nand2_1 U11497 ( .ip1(n10182), .ip2(i_i2c_U_dff_tx_mem[66]), .op(n10183) );
  nand4_1 U11498 ( .ip1(n10186), .ip2(n10185), .ip3(n10184), .ip4(n10183), 
        .op(n10187) );
  not_ab_or_c_or_d U11499 ( .ip1(n10189), .ip2(i_i2c_U_dff_tx_mem[12]), .ip3(
        n10188), .ip4(n10187), .op(n10192) );
  nand2_1 U11500 ( .ip1(n10190), .ip2(i_i2c_U_dff_tx_mem[39]), .op(n10191) );
  nand3_1 U11501 ( .ip1(n10193), .ip2(n10192), .ip3(n10191), .op(n10194) );
  mux2_1 U11502 ( .ip1(i_i2c_tx_fifo_data_buf[3]), .ip2(n10194), .s(
        i_i2c_U_DW_apb_i2c_tx_shift_N90), .op(n5219) );
  not_ab_or_c_or_d U11503 ( .ip1(n11216), .ip2(n10195), .ip3(n11215), .ip4(
        n11026), .op(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N38) );
  inv_1 U11504 ( .ip(n10199), .op(n10197) );
  nand2_1 U11505 ( .ip1(n10197), .ip2(i_ssi_U_fifo_U_tx_fifo_wr_addr_at_max), 
        .op(n10196) );
  nand2_1 U11506 ( .ip1(n10196), .ip2(n10759), .op(n10205) );
  not_ab_or_c_or_d U11507 ( .ip1(n10220), .ip2(n10203), .ip3(n10205), .ip4(
        n5608), .op(i_ssi_U_fifo_U_tx_fifo_N43) );
  nor2_1 U11508 ( .ip1(n10198), .ip2(n10197), .op(n10200) );
  nor2_1 U11509 ( .ip1(n10200), .ip2(n10226), .op(n10201) );
  nor2_1 U11510 ( .ip1(n10201), .ip2(n10205), .op(n11848) );
  nand2_1 U11511 ( .ip1(i_ssi_tx_wr_addr[1]), .ip2(i_ssi_tx_wr_addr[2]), .op(
        n10224) );
  inv_1 U11512 ( .ip(n11848), .op(n10202) );
  nor2_1 U11513 ( .ip1(n10224), .ip2(n10202), .op(i_ssi_U_fifo_U_tx_fifo_N40)
         );
  inv_1 U11514 ( .ip(n10228), .op(n10206) );
  inv_1 U11515 ( .ip(i_ssi_tx_wr_addr[1]), .op(n10221) );
  inv_1 U11516 ( .ip(n10203), .op(n10204) );
  not_ab_or_c_or_d U11517 ( .ip1(n10206), .ip2(n10221), .ip3(n10205), .ip4(
        n10204), .op(i_ssi_U_fifo_U_tx_fifo_N42) );
  mux2_1 U11518 ( .ip1(i_ssi_U_dff_tx_mem[66]), .ip2(i_apb_pwdata_int[2]), .s(
        n10354), .op(n4510) );
  nand2_1 U11519 ( .ip1(i_ssi_tx_rd_addr[0]), .ip2(i_ssi_tx_rd_addr[1]), .op(
        n10244) );
  nor2_1 U11520 ( .ip1(n5588), .ip2(n10244), .op(n10213) );
  inv_1 U11521 ( .ip(i_ssi_U_fifo_U_tx_fifo_rd_addr_at_max), .op(n10208) );
  nand2_1 U11522 ( .ip1(n10208), .ip2(i_ssi_tx_rd_addr[0]), .op(n10207) );
  nor2_1 U11523 ( .ip1(n10207), .ip2(n5588), .op(n10210) );
  inv_1 U11524 ( .ip(i_ssi_tx_rd_addr[1]), .op(n10239) );
  nor2_1 U11525 ( .ip1(n10208), .ip2(n5588), .op(n10215) );
  nor2_1 U11526 ( .ip1(n10239), .ip2(n10215), .op(n10209) );
  nor2_1 U11527 ( .ip1(n10210), .ip2(n10209), .op(n10211) );
  nor2_1 U11528 ( .ip1(n10213), .ip2(n10211), .op(n10212) );
  and2_1 U11529 ( .ip1(n10759), .ip2(n10212), .op(i_ssi_U_fifo_U_tx_fifo_N45)
         );
  inv_1 U11530 ( .ip(i_ssi_tx_rd_addr[2]), .op(n10243) );
  xor2_1 U11531 ( .ip1(n10243), .ip2(n10213), .op(n10214) );
  nor3_1 U11532 ( .ip1(n10215), .ip2(n10214), .ip3(n10748), .op(
        i_ssi_U_fifo_U_tx_fifo_N46) );
  nor2_1 U11533 ( .ip1(i_ssi_tx_rd_addr[0]), .ip2(
        i_ssi_U_fifo_U_tx_fifo_rd_addr_at_max), .op(n10217) );
  mux2_1 U11534 ( .ip1(n10217), .ip2(i_ssi_tx_rd_addr[0]), .s(n5588), .op(
        n10218) );
  and2_1 U11535 ( .ip1(n10759), .ip2(n10218), .op(n11847) );
  nand2_1 U11536 ( .ip1(i_ssi_tx_rd_addr[1]), .ip2(i_ssi_tx_rd_addr[2]), .op(
        n10241) );
  inv_1 U11537 ( .ip(n11847), .op(n10219) );
  nor2_1 U11538 ( .ip1(n10241), .ip2(n10219), .op(i_ssi_U_fifo_U_tx_fifo_N39)
         );
  nor2_1 U11539 ( .ip1(i_ssi_tx_wr_addr[2]), .ip2(i_ssi_tx_wr_addr[1]), .op(
        n10227) );
  mux2_1 U11540 ( .ip1(i_apb_pwdata_int[2]), .ip2(i_ssi_U_dff_tx_mem[114]), 
        .s(n5254), .op(n4462) );
  mux2_1 U11541 ( .ip1(i_ssi_U_dff_tx_mem[2]), .ip2(i_apb_pwdata_int[2]), .s(
        n5608), .op(n4574) );
  nor2_1 U11542 ( .ip1(i_ssi_tx_wr_addr[1]), .ip2(n10220), .op(n10223) );
  mux2_1 U11543 ( .ip1(i_apb_pwdata_int[2]), .ip2(i_ssi_U_dff_tx_mem[34]), .s(
        n10365), .op(n4542) );
  nor2_1 U11544 ( .ip1(i_ssi_tx_wr_addr[2]), .ip2(n10221), .op(n10222) );
  mux2_1 U11545 ( .ip1(i_apb_pwdata_int[2]), .ip2(i_ssi_U_dff_tx_mem[82]), .s(
        n5255), .op(n4494) );
  mux2_1 U11546 ( .ip1(i_apb_pwdata_int[2]), .ip2(i_ssi_U_dff_tx_mem[50]), .s(
        n5253), .op(n4526) );
  inv_1 U11547 ( .ip(n10224), .op(n10225) );
  mux2_1 U11548 ( .ip1(i_apb_pwdata_int[2]), .ip2(i_ssi_U_dff_tx_mem[18]), .s(
        n5256), .op(n4558) );
  mux2_1 U11549 ( .ip1(i_apb_pwdata_int[2]), .ip2(i_ssi_U_dff_tx_mem[98]), .s(
        n5286), .op(n4478) );
  mux2_1 U11550 ( .ip1(i_ssi_U_dff_tx_mem[64]), .ip2(i_apb_pwdata_int[0]), .s(
        n10354), .op(n4512) );
  mux2_1 U11551 ( .ip1(i_apb_pwdata_int[0]), .ip2(i_ssi_U_dff_tx_mem[112]), 
        .s(n5254), .op(n4464) );
  mux2_1 U11552 ( .ip1(i_ssi_U_dff_tx_mem[0]), .ip2(i_apb_pwdata_int[0]), .s(
        n5608), .op(n4576) );
  mux2_1 U11553 ( .ip1(i_apb_pwdata_int[0]), .ip2(i_ssi_U_dff_tx_mem[32]), .s(
        n10365), .op(n4544) );
  mux2_1 U11554 ( .ip1(i_apb_pwdata_int[0]), .ip2(i_ssi_U_dff_tx_mem[80]), .s(
        n5255), .op(n4496) );
  mux2_1 U11555 ( .ip1(i_apb_pwdata_int[0]), .ip2(i_ssi_U_dff_tx_mem[48]), .s(
        n5253), .op(n4528) );
  mux2_1 U11556 ( .ip1(i_apb_pwdata_int[0]), .ip2(i_ssi_U_dff_tx_mem[16]), .s(
        n5256), .op(n4560) );
  mux2_1 U11557 ( .ip1(i_apb_pwdata_int[0]), .ip2(i_ssi_U_dff_tx_mem[96]), .s(
        n5286), .op(n4480) );
  mux2_1 U11558 ( .ip1(i_apb_pwdata_int[1]), .ip2(i_ssi_U_dff_tx_mem[113]), 
        .s(n5254), .op(n4463) );
  mux2_1 U11559 ( .ip1(i_apb_pwdata_int[1]), .ip2(i_ssi_U_dff_tx_mem[33]), .s(
        n10365), .op(n4543) );
  mux2_1 U11560 ( .ip1(i_apb_pwdata_int[1]), .ip2(i_ssi_U_dff_tx_mem[81]), .s(
        n5255), .op(n4495) );
  mux2_1 U11561 ( .ip1(i_apb_pwdata_int[1]), .ip2(i_ssi_U_dff_tx_mem[49]), .s(
        n5253), .op(n4527) );
  mux2_1 U11562 ( .ip1(i_apb_pwdata_int[1]), .ip2(i_ssi_U_dff_tx_mem[17]), .s(
        n5256), .op(n4559) );
  mux2_1 U11563 ( .ip1(i_apb_pwdata_int[1]), .ip2(i_ssi_U_dff_tx_mem[97]), .s(
        n5286), .op(n4479) );
  mux2_1 U11564 ( .ip1(i_ssi_U_dff_tx_mem[67]), .ip2(i_apb_pwdata_int[3]), .s(
        n10354), .op(n4509) );
  mux2_1 U11565 ( .ip1(i_apb_pwdata_int[3]), .ip2(i_ssi_U_dff_tx_mem[115]), 
        .s(n5254), .op(n4461) );
  mux2_1 U11566 ( .ip1(i_apb_pwdata_int[3]), .ip2(i_ssi_U_dff_tx_mem[35]), .s(
        n10365), .op(n4541) );
  mux2_1 U11567 ( .ip1(i_apb_pwdata_int[3]), .ip2(i_ssi_U_dff_tx_mem[83]), .s(
        n5255), .op(n4493) );
  mux2_1 U11568 ( .ip1(i_apb_pwdata_int[3]), .ip2(i_ssi_U_dff_tx_mem[51]), .s(
        n5253), .op(n4525) );
  mux2_1 U11569 ( .ip1(i_apb_pwdata_int[3]), .ip2(i_ssi_U_dff_tx_mem[19]), .s(
        n5256), .op(n4557) );
  mux2_1 U11570 ( .ip1(i_apb_pwdata_int[3]), .ip2(i_ssi_U_dff_tx_mem[99]), .s(
        n5286), .op(n4477) );
  nand2_1 U11571 ( .ip1(n10230), .ip2(i_ssi_sclk_re), .op(n10232) );
  nor2_1 U11572 ( .ip1(n10232), .ip2(n10231), .op(i_ssi_load_start_bit) );
  nand2_1 U11573 ( .ip1(n10400), .ip2(i_ssi_U_dff_tx_mem[82]), .op(n10238) );
  and3_1 U11574 ( .ip1(n10239), .ip2(i_ssi_tx_rd_addr[0]), .ip3(n10243), .op(
        n10401) );
  nand2_1 U11575 ( .ip1(n10401), .ip2(i_ssi_U_dff_tx_mem[98]), .op(n10237) );
  inv_1 U11576 ( .ip(i_ssi_tx_rd_addr[0]), .op(n10233) );
  nand2_1 U11577 ( .ip1(n10402), .ip2(i_ssi_U_dff_tx_mem[50]), .op(n10236) );
  nand2_1 U11578 ( .ip1(n10389), .ip2(i_ssi_U_dff_tx_mem[34]), .op(n10235) );
  and2_1 U11579 ( .ip1(n10240), .ip2(n10239), .op(n10407) );
  nand2_1 U11580 ( .ip1(n10407), .ip2(i_ssi_U_dff_tx_mem[114]), .op(n10248) );
  nor2_1 U11581 ( .ip1(i_ssi_tx_rd_addr[0]), .ip2(n10241), .op(n10408) );
  inv_1 U11582 ( .ip(n10408), .op(n10242) );
  inv_1 U11583 ( .ip(n10242), .op(n10370) );
  nand2_1 U11584 ( .ip1(n10370), .ip2(i_ssi_U_dff_tx_mem[18]), .op(n10247) );
  nand2_1 U11585 ( .ip1(n5609), .ip2(i_ssi_U_dff_tx_mem[2]), .op(n10246) );
  nand2_1 U11586 ( .ip1(n5252), .ip2(i_ssi_U_dff_tx_mem[66]), .op(n10245) );
  or2_1 U11587 ( .ip1(n10250), .ip2(n10249), .op(n10652) );
  mux2_1 U11588 ( .ip1(n10652), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[2]), 
        .s(n10377), .op(n4418) );
  and2_1 U11589 ( .ip1(n10370), .ip2(i_ssi_U_dff_tx_mem[17]), .op(n10254) );
  nand2_1 U11590 ( .ip1(n5609), .ip2(i_ssi_U_dff_tx_mem[1]), .op(n10252) );
  nand2_1 U11591 ( .ip1(n5252), .ip2(i_ssi_U_dff_tx_mem[65]), .op(n10251) );
  nand2_1 U11592 ( .ip1(n10252), .ip2(n10251), .op(n10253) );
  not_ab_or_c_or_d U11593 ( .ip1(n10407), .ip2(i_ssi_U_dff_tx_mem[113]), .ip3(
        n10254), .ip4(n10253), .op(n10260) );
  and2_1 U11594 ( .ip1(n10401), .ip2(i_ssi_U_dff_tx_mem[97]), .op(n10258) );
  nand2_1 U11595 ( .ip1(n10402), .ip2(i_ssi_U_dff_tx_mem[49]), .op(n10256) );
  nand2_1 U11596 ( .ip1(n10389), .ip2(i_ssi_U_dff_tx_mem[33]), .op(n10255) );
  nand2_1 U11597 ( .ip1(n10256), .ip2(n10255), .op(n10257) );
  not_ab_or_c_or_d U11598 ( .ip1(n10400), .ip2(i_ssi_U_dff_tx_mem[81]), .ip3(
        n10258), .ip4(n10257), .op(n10259) );
  nand2_1 U11599 ( .ip1(n10260), .ip2(n10259), .op(n10650) );
  mux2_1 U11600 ( .ip1(n10650), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[1]), 
        .s(n10377), .op(n4419) );
  and2_1 U11601 ( .ip1(n10370), .ip2(i_ssi_U_dff_tx_mem[16]), .op(n10264) );
  nand2_1 U11602 ( .ip1(n5609), .ip2(i_ssi_U_dff_tx_mem[0]), .op(n10262) );
  nand2_1 U11603 ( .ip1(n5252), .ip2(i_ssi_U_dff_tx_mem[64]), .op(n10261) );
  nand2_1 U11604 ( .ip1(n10262), .ip2(n10261), .op(n10263) );
  not_ab_or_c_or_d U11605 ( .ip1(n10407), .ip2(i_ssi_U_dff_tx_mem[112]), .ip3(
        n10264), .ip4(n10263), .op(n10270) );
  and2_1 U11606 ( .ip1(n10401), .ip2(i_ssi_U_dff_tx_mem[96]), .op(n10268) );
  nand2_1 U11607 ( .ip1(n10402), .ip2(i_ssi_U_dff_tx_mem[48]), .op(n10266) );
  nand2_1 U11608 ( .ip1(n10389), .ip2(i_ssi_U_dff_tx_mem[32]), .op(n10265) );
  nand2_1 U11609 ( .ip1(n10266), .ip2(n10265), .op(n10267) );
  not_ab_or_c_or_d U11610 ( .ip1(n10400), .ip2(i_ssi_U_dff_tx_mem[80]), .ip3(
        n10268), .ip4(n10267), .op(n10269) );
  nand2_1 U11611 ( .ip1(n10270), .ip2(n10269), .op(n10653) );
  inv_2 U11612 ( .ip(n10415), .op(n10377) );
  mux2_1 U11613 ( .ip1(n10653), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[0]), 
        .s(n10377), .op(n4420) );
  inv_1 U11614 ( .ip(n10271), .op(n10272) );
  nand2_1 U11615 ( .ip1(n10272), .ip2(i_ssi_U_mstfsm_spi1_control), .op(n10273) );
  nand2_1 U11616 ( .ip1(n10273), .ip2(n5492), .op(n4194) );
  mux2_1 U11617 ( .ip1(i_ssi_U_dff_tx_mem[79]), .ip2(i_apb_pwdata_int[15]), 
        .s(n10354), .op(n4497) );
  mux2_1 U11618 ( .ip1(i_apb_pwdata_int[15]), .ip2(i_ssi_U_dff_tx_mem[127]), 
        .s(n5254), .op(n4449) );
  mux2_1 U11619 ( .ip1(i_ssi_U_dff_tx_mem[15]), .ip2(i_apb_pwdata_int[15]), 
        .s(n5608), .op(n4561) );
  mux2_1 U11620 ( .ip1(i_apb_pwdata_int[15]), .ip2(i_ssi_U_dff_tx_mem[47]), 
        .s(n10365), .op(n4529) );
  mux2_1 U11621 ( .ip1(i_apb_pwdata_int[15]), .ip2(i_ssi_U_dff_tx_mem[95]), 
        .s(n5255), .op(n4481) );
  mux2_1 U11622 ( .ip1(i_apb_pwdata_int[15]), .ip2(i_ssi_U_dff_tx_mem[63]), 
        .s(n5253), .op(n4513) );
  mux2_1 U11623 ( .ip1(i_apb_pwdata_int[15]), .ip2(i_ssi_U_dff_tx_mem[31]), 
        .s(n5256), .op(n4545) );
  mux2_1 U11624 ( .ip1(i_apb_pwdata_int[15]), .ip2(i_ssi_U_dff_tx_mem[111]), 
        .s(n5286), .op(n4465) );
  nand2_1 U11625 ( .ip1(n10400), .ip2(i_ssi_U_dff_tx_mem[95]), .op(n10277) );
  nand2_1 U11626 ( .ip1(n10401), .ip2(i_ssi_U_dff_tx_mem[111]), .op(n10276) );
  nand2_1 U11627 ( .ip1(n10402), .ip2(i_ssi_U_dff_tx_mem[63]), .op(n10275) );
  nand2_1 U11628 ( .ip1(n10389), .ip2(i_ssi_U_dff_tx_mem[47]), .op(n10274) );
  nand2_1 U11629 ( .ip1(n10407), .ip2(i_ssi_U_dff_tx_mem[127]), .op(n10281) );
  nand2_1 U11630 ( .ip1(n10370), .ip2(i_ssi_U_dff_tx_mem[31]), .op(n10280) );
  nand2_1 U11631 ( .ip1(n5609), .ip2(i_ssi_U_dff_tx_mem[15]), .op(n10279) );
  nand2_1 U11632 ( .ip1(n5252), .ip2(i_ssi_U_dff_tx_mem[79]), .op(n10278) );
  or2_1 U11633 ( .ip1(n10283), .ip2(n10282), .op(n10617) );
  mux2_1 U11634 ( .ip1(n10617), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[15]), 
        .s(n10377), .op(n4405) );
  mux2_1 U11635 ( .ip1(i_ssi_U_dff_tx_mem[78]), .ip2(i_apb_pwdata_int[14]), 
        .s(n10354), .op(n4498) );
  mux2_1 U11636 ( .ip1(i_apb_pwdata_int[14]), .ip2(i_ssi_U_dff_tx_mem[126]), 
        .s(n5254), .op(n4450) );
  mux2_1 U11637 ( .ip1(i_ssi_U_dff_tx_mem[14]), .ip2(i_apb_pwdata_int[14]), 
        .s(n5608), .op(n4562) );
  mux2_1 U11638 ( .ip1(i_apb_pwdata_int[14]), .ip2(i_ssi_U_dff_tx_mem[46]), 
        .s(n10365), .op(n4530) );
  mux2_1 U11639 ( .ip1(i_apb_pwdata_int[14]), .ip2(i_ssi_U_dff_tx_mem[94]), 
        .s(n5255), .op(n4482) );
  mux2_1 U11640 ( .ip1(i_apb_pwdata_int[14]), .ip2(i_ssi_U_dff_tx_mem[62]), 
        .s(n5253), .op(n4514) );
  mux2_1 U11641 ( .ip1(i_apb_pwdata_int[14]), .ip2(i_ssi_U_dff_tx_mem[30]), 
        .s(n5256), .op(n4546) );
  mux2_1 U11642 ( .ip1(i_apb_pwdata_int[14]), .ip2(i_ssi_U_dff_tx_mem[110]), 
        .s(n5286), .op(n4466) );
  nand2_1 U11643 ( .ip1(n10400), .ip2(i_ssi_U_dff_tx_mem[94]), .op(n10287) );
  nand2_1 U11644 ( .ip1(n10401), .ip2(i_ssi_U_dff_tx_mem[110]), .op(n10286) );
  nand2_1 U11645 ( .ip1(n10402), .ip2(i_ssi_U_dff_tx_mem[62]), .op(n10285) );
  nand2_1 U11646 ( .ip1(n10389), .ip2(i_ssi_U_dff_tx_mem[46]), .op(n10284) );
  nand2_1 U11647 ( .ip1(n10407), .ip2(i_ssi_U_dff_tx_mem[126]), .op(n10291) );
  nand2_1 U11648 ( .ip1(n10370), .ip2(i_ssi_U_dff_tx_mem[30]), .op(n10290) );
  nand2_1 U11649 ( .ip1(n5609), .ip2(i_ssi_U_dff_tx_mem[14]), .op(n10289) );
  nand2_1 U11650 ( .ip1(n5252), .ip2(i_ssi_U_dff_tx_mem[78]), .op(n10288) );
  or2_1 U11651 ( .ip1(n10293), .ip2(n10292), .op(n10614) );
  mux2_1 U11652 ( .ip1(n10614), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[14]), 
        .s(n10377), .op(n4406) );
  mux2_1 U11653 ( .ip1(i_apb_pwdata_int[13]), .ip2(i_ssi_U_dff_tx_mem[125]), 
        .s(n5254), .op(n4451) );
  mux2_1 U11654 ( .ip1(i_apb_pwdata_int[13]), .ip2(i_ssi_U_dff_tx_mem[45]), 
        .s(n10365), .op(n4531) );
  mux2_1 U11655 ( .ip1(i_apb_pwdata_int[13]), .ip2(i_ssi_U_dff_tx_mem[93]), 
        .s(n5255), .op(n4483) );
  mux2_1 U11656 ( .ip1(i_apb_pwdata_int[13]), .ip2(i_ssi_U_dff_tx_mem[61]), 
        .s(n5253), .op(n4515) );
  mux2_1 U11657 ( .ip1(i_apb_pwdata_int[13]), .ip2(i_ssi_U_dff_tx_mem[29]), 
        .s(n5256), .op(n4547) );
  mux2_1 U11658 ( .ip1(i_apb_pwdata_int[13]), .ip2(i_ssi_U_dff_tx_mem[109]), 
        .s(n5286), .op(n4467) );
  nand2_1 U11659 ( .ip1(n10400), .ip2(i_ssi_U_dff_tx_mem[93]), .op(n10297) );
  nand2_1 U11660 ( .ip1(n10401), .ip2(i_ssi_U_dff_tx_mem[109]), .op(n10296) );
  nand2_1 U11661 ( .ip1(n10402), .ip2(i_ssi_U_dff_tx_mem[61]), .op(n10295) );
  nand2_1 U11662 ( .ip1(n10389), .ip2(i_ssi_U_dff_tx_mem[45]), .op(n10294) );
  nand2_1 U11663 ( .ip1(n10407), .ip2(i_ssi_U_dff_tx_mem[125]), .op(n10301) );
  nand2_1 U11664 ( .ip1(n10408), .ip2(i_ssi_U_dff_tx_mem[29]), .op(n10300) );
  nand2_1 U11665 ( .ip1(n5609), .ip2(i_ssi_U_dff_tx_mem[13]), .op(n10299) );
  nand2_1 U11666 ( .ip1(n5252), .ip2(i_ssi_U_dff_tx_mem[77]), .op(n10298) );
  or2_1 U11667 ( .ip1(n10303), .ip2(n10302), .op(n10622) );
  mux2_1 U11668 ( .ip1(n10622), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[13]), 
        .s(n10377), .op(n4407) );
  mux2_1 U11669 ( .ip1(i_ssi_U_dff_tx_mem[76]), .ip2(i_apb_pwdata_int[12]), 
        .s(n10354), .op(n4500) );
  mux2_1 U11670 ( .ip1(i_apb_pwdata_int[12]), .ip2(i_ssi_U_dff_tx_mem[124]), 
        .s(n5254), .op(n4452) );
  mux2_1 U11671 ( .ip1(i_ssi_U_dff_tx_mem[12]), .ip2(i_apb_pwdata_int[12]), 
        .s(n5608), .op(n4564) );
  mux2_1 U11672 ( .ip1(i_apb_pwdata_int[12]), .ip2(i_ssi_U_dff_tx_mem[44]), 
        .s(n10365), .op(n4532) );
  mux2_1 U11673 ( .ip1(i_apb_pwdata_int[12]), .ip2(i_ssi_U_dff_tx_mem[92]), 
        .s(n5255), .op(n4484) );
  mux2_1 U11674 ( .ip1(i_apb_pwdata_int[12]), .ip2(i_ssi_U_dff_tx_mem[60]), 
        .s(n5253), .op(n4516) );
  mux2_1 U11675 ( .ip1(i_apb_pwdata_int[12]), .ip2(i_ssi_U_dff_tx_mem[28]), 
        .s(n5256), .op(n4548) );
  mux2_1 U11676 ( .ip1(i_apb_pwdata_int[12]), .ip2(i_ssi_U_dff_tx_mem[108]), 
        .s(n5286), .op(n4468) );
  nand2_1 U11677 ( .ip1(n10400), .ip2(i_ssi_U_dff_tx_mem[92]), .op(n10307) );
  nand2_1 U11678 ( .ip1(n10401), .ip2(i_ssi_U_dff_tx_mem[108]), .op(n10306) );
  nand2_1 U11679 ( .ip1(n10402), .ip2(i_ssi_U_dff_tx_mem[60]), .op(n10305) );
  nand2_1 U11680 ( .ip1(n10389), .ip2(i_ssi_U_dff_tx_mem[44]), .op(n10304) );
  nand2_1 U11681 ( .ip1(n10407), .ip2(i_ssi_U_dff_tx_mem[124]), .op(n10311) );
  nand2_1 U11682 ( .ip1(n10370), .ip2(i_ssi_U_dff_tx_mem[28]), .op(n10310) );
  nand2_1 U11683 ( .ip1(n5609), .ip2(i_ssi_U_dff_tx_mem[12]), .op(n10309) );
  nand2_1 U11684 ( .ip1(n5252), .ip2(i_ssi_U_dff_tx_mem[76]), .op(n10308) );
  or2_1 U11685 ( .ip1(n10313), .ip2(n10312), .op(n10616) );
  mux2_1 U11686 ( .ip1(n10616), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[12]), 
        .s(n10377), .op(n4408) );
  mux2_1 U11687 ( .ip1(i_ssi_U_dff_tx_mem[75]), .ip2(i_apb_pwdata_int[11]), 
        .s(n10354), .op(n4501) );
  mux2_1 U11688 ( .ip1(i_apb_pwdata_int[11]), .ip2(i_ssi_U_dff_tx_mem[123]), 
        .s(n5254), .op(n4453) );
  mux2_1 U11689 ( .ip1(i_ssi_U_dff_tx_mem[11]), .ip2(i_apb_pwdata_int[11]), 
        .s(n5608), .op(n4565) );
  mux2_1 U11690 ( .ip1(i_apb_pwdata_int[11]), .ip2(i_ssi_U_dff_tx_mem[43]), 
        .s(n10365), .op(n4533) );
  mux2_1 U11691 ( .ip1(i_apb_pwdata_int[11]), .ip2(i_ssi_U_dff_tx_mem[91]), 
        .s(n5255), .op(n4485) );
  mux2_1 U11692 ( .ip1(i_apb_pwdata_int[11]), .ip2(i_ssi_U_dff_tx_mem[59]), 
        .s(n5253), .op(n4517) );
  mux2_1 U11693 ( .ip1(i_apb_pwdata_int[11]), .ip2(i_ssi_U_dff_tx_mem[27]), 
        .s(n5256), .op(n4549) );
  mux2_1 U11694 ( .ip1(i_apb_pwdata_int[11]), .ip2(i_ssi_U_dff_tx_mem[107]), 
        .s(n5286), .op(n4469) );
  nand2_1 U11695 ( .ip1(n10400), .ip2(i_ssi_U_dff_tx_mem[91]), .op(n10317) );
  nand2_1 U11696 ( .ip1(n10401), .ip2(i_ssi_U_dff_tx_mem[107]), .op(n10316) );
  nand2_1 U11697 ( .ip1(n10402), .ip2(i_ssi_U_dff_tx_mem[59]), .op(n10315) );
  nand2_1 U11698 ( .ip1(n10389), .ip2(i_ssi_U_dff_tx_mem[43]), .op(n10314) );
  nand2_1 U11699 ( .ip1(n10407), .ip2(i_ssi_U_dff_tx_mem[123]), .op(n10321) );
  nand2_1 U11700 ( .ip1(n10370), .ip2(i_ssi_U_dff_tx_mem[27]), .op(n10320) );
  nand2_1 U11701 ( .ip1(n5609), .ip2(i_ssi_U_dff_tx_mem[11]), .op(n10319) );
  nand2_1 U11702 ( .ip1(n5252), .ip2(i_ssi_U_dff_tx_mem[75]), .op(n10318) );
  or2_1 U11703 ( .ip1(n10323), .ip2(n10322), .op(n10659) );
  mux2_1 U11704 ( .ip1(n10659), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[11]), 
        .s(n10377), .op(n4409) );
  mux2_1 U11705 ( .ip1(i_apb_pwdata_int[10]), .ip2(i_ssi_U_dff_tx_mem[122]), 
        .s(n5254), .op(n4454) );
  mux2_1 U11706 ( .ip1(i_apb_pwdata_int[10]), .ip2(i_ssi_U_dff_tx_mem[42]), 
        .s(n10365), .op(n4534) );
  mux2_1 U11707 ( .ip1(i_apb_pwdata_int[10]), .ip2(i_ssi_U_dff_tx_mem[90]), 
        .s(n5255), .op(n4486) );
  mux2_1 U11708 ( .ip1(i_apb_pwdata_int[10]), .ip2(i_ssi_U_dff_tx_mem[58]), 
        .s(n5253), .op(n4518) );
  mux2_1 U11709 ( .ip1(i_apb_pwdata_int[10]), .ip2(i_ssi_U_dff_tx_mem[26]), 
        .s(n5256), .op(n4550) );
  mux2_1 U11710 ( .ip1(i_apb_pwdata_int[10]), .ip2(i_ssi_U_dff_tx_mem[106]), 
        .s(n5286), .op(n4470) );
  nand2_1 U11711 ( .ip1(n10400), .ip2(i_ssi_U_dff_tx_mem[90]), .op(n10327) );
  nand2_1 U11712 ( .ip1(n10401), .ip2(i_ssi_U_dff_tx_mem[106]), .op(n10326) );
  nand2_1 U11713 ( .ip1(n10402), .ip2(i_ssi_U_dff_tx_mem[58]), .op(n10325) );
  nand2_1 U11714 ( .ip1(n10389), .ip2(i_ssi_U_dff_tx_mem[42]), .op(n10324) );
  nand2_1 U11715 ( .ip1(n10407), .ip2(i_ssi_U_dff_tx_mem[122]), .op(n10331) );
  nand2_1 U11716 ( .ip1(n10408), .ip2(i_ssi_U_dff_tx_mem[26]), .op(n10330) );
  nand2_1 U11717 ( .ip1(n5609), .ip2(i_ssi_U_dff_tx_mem[10]), .op(n10329) );
  nand2_1 U11718 ( .ip1(n5252), .ip2(i_ssi_U_dff_tx_mem[74]), .op(n10328) );
  or2_1 U11719 ( .ip1(n10333), .ip2(n10332), .op(n10661) );
  mux2_1 U11720 ( .ip1(n10661), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[10]), 
        .s(n10377), .op(n4410) );
  mux2_1 U11721 ( .ip1(i_ssi_U_dff_tx_mem[73]), .ip2(i_apb_pwdata_int[9]), .s(
        n10354), .op(n4503) );
  mux2_1 U11722 ( .ip1(i_apb_pwdata_int[9]), .ip2(i_ssi_U_dff_tx_mem[121]), 
        .s(n5254), .op(n4455) );
  mux2_1 U11723 ( .ip1(i_ssi_U_dff_tx_mem[9]), .ip2(i_apb_pwdata_int[9]), .s(
        n5608), .op(n4567) );
  mux2_1 U11724 ( .ip1(i_apb_pwdata_int[9]), .ip2(i_ssi_U_dff_tx_mem[41]), .s(
        n10365), .op(n4535) );
  mux2_1 U11725 ( .ip1(i_apb_pwdata_int[9]), .ip2(i_ssi_U_dff_tx_mem[89]), .s(
        n5255), .op(n4487) );
  mux2_1 U11726 ( .ip1(i_apb_pwdata_int[9]), .ip2(i_ssi_U_dff_tx_mem[57]), .s(
        n5253), .op(n4519) );
  mux2_1 U11727 ( .ip1(i_apb_pwdata_int[9]), .ip2(i_ssi_U_dff_tx_mem[25]), .s(
        n5256), .op(n4551) );
  mux2_1 U11728 ( .ip1(i_apb_pwdata_int[9]), .ip2(i_ssi_U_dff_tx_mem[105]), 
        .s(n5286), .op(n4471) );
  nand2_1 U11729 ( .ip1(n10400), .ip2(i_ssi_U_dff_tx_mem[89]), .op(n10337) );
  nand2_1 U11730 ( .ip1(n10401), .ip2(i_ssi_U_dff_tx_mem[105]), .op(n10336) );
  nand2_1 U11731 ( .ip1(n10402), .ip2(i_ssi_U_dff_tx_mem[57]), .op(n10335) );
  nand2_1 U11732 ( .ip1(n10389), .ip2(i_ssi_U_dff_tx_mem[41]), .op(n10334) );
  nand2_1 U11733 ( .ip1(n10407), .ip2(i_ssi_U_dff_tx_mem[121]), .op(n10341) );
  nand2_1 U11734 ( .ip1(n10370), .ip2(i_ssi_U_dff_tx_mem[25]), .op(n10340) );
  nand2_1 U11735 ( .ip1(n5609), .ip2(i_ssi_U_dff_tx_mem[9]), .op(n10339) );
  nand2_1 U11736 ( .ip1(n5252), .ip2(i_ssi_U_dff_tx_mem[73]), .op(n10338) );
  or2_1 U11737 ( .ip1(n10343), .ip2(n10342), .op(n10658) );
  mux2_1 U11738 ( .ip1(n10658), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[9]), 
        .s(n10377), .op(n4411) );
  mux2_1 U11739 ( .ip1(i_ssi_U_dff_tx_mem[72]), .ip2(i_apb_pwdata_int[8]), .s(
        n10354), .op(n4504) );
  mux2_1 U11740 ( .ip1(i_apb_pwdata_int[8]), .ip2(i_ssi_U_dff_tx_mem[120]), 
        .s(n5254), .op(n4456) );
  mux2_1 U11741 ( .ip1(i_ssi_U_dff_tx_mem[8]), .ip2(i_apb_pwdata_int[8]), .s(
        n5608), .op(n4568) );
  mux2_1 U11742 ( .ip1(i_apb_pwdata_int[8]), .ip2(i_ssi_U_dff_tx_mem[40]), .s(
        n10365), .op(n4536) );
  mux2_1 U11743 ( .ip1(i_apb_pwdata_int[8]), .ip2(i_ssi_U_dff_tx_mem[88]), .s(
        n5255), .op(n4488) );
  mux2_1 U11744 ( .ip1(i_apb_pwdata_int[8]), .ip2(i_ssi_U_dff_tx_mem[56]), .s(
        n5253), .op(n4520) );
  mux2_1 U11745 ( .ip1(i_apb_pwdata_int[8]), .ip2(i_ssi_U_dff_tx_mem[24]), .s(
        n5256), .op(n4552) );
  mux2_1 U11746 ( .ip1(i_apb_pwdata_int[8]), .ip2(i_ssi_U_dff_tx_mem[104]), 
        .s(n5286), .op(n4472) );
  nand2_1 U11747 ( .ip1(n10400), .ip2(i_ssi_U_dff_tx_mem[88]), .op(n10347) );
  nand2_1 U11748 ( .ip1(n10401), .ip2(i_ssi_U_dff_tx_mem[104]), .op(n10346) );
  nand2_1 U11749 ( .ip1(n10402), .ip2(i_ssi_U_dff_tx_mem[56]), .op(n10345) );
  nand2_1 U11750 ( .ip1(n10389), .ip2(i_ssi_U_dff_tx_mem[40]), .op(n10344) );
  nand2_1 U11751 ( .ip1(n10407), .ip2(i_ssi_U_dff_tx_mem[120]), .op(n10351) );
  nand2_1 U11752 ( .ip1(n10370), .ip2(i_ssi_U_dff_tx_mem[24]), .op(n10350) );
  nand2_1 U11753 ( .ip1(n5609), .ip2(i_ssi_U_dff_tx_mem[8]), .op(n10349) );
  nand2_1 U11754 ( .ip1(n5252), .ip2(i_ssi_U_dff_tx_mem[72]), .op(n10348) );
  or2_1 U11755 ( .ip1(n10353), .ip2(n10352), .op(n10662) );
  mux2_1 U11756 ( .ip1(n10662), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[8]), 
        .s(n10377), .op(n4412) );
  mux2_1 U11757 ( .ip1(i_ssi_U_dff_tx_mem[71]), .ip2(i_apb_pwdata_int[7]), .s(
        n10354), .op(n4505) );
  mux2_1 U11758 ( .ip1(i_apb_pwdata_int[7]), .ip2(i_ssi_U_dff_tx_mem[119]), 
        .s(n5254), .op(n4457) );
  mux2_1 U11759 ( .ip1(i_ssi_U_dff_tx_mem[7]), .ip2(i_apb_pwdata_int[7]), .s(
        n5608), .op(n4569) );
  mux2_1 U11760 ( .ip1(i_apb_pwdata_int[7]), .ip2(i_ssi_U_dff_tx_mem[39]), .s(
        n10365), .op(n4537) );
  mux2_1 U11761 ( .ip1(i_apb_pwdata_int[7]), .ip2(i_ssi_U_dff_tx_mem[87]), .s(
        n5255), .op(n4489) );
  mux2_1 U11762 ( .ip1(i_apb_pwdata_int[7]), .ip2(i_ssi_U_dff_tx_mem[55]), .s(
        n5253), .op(n4521) );
  mux2_1 U11763 ( .ip1(i_apb_pwdata_int[7]), .ip2(i_ssi_U_dff_tx_mem[23]), .s(
        n5256), .op(n4553) );
  mux2_1 U11764 ( .ip1(i_apb_pwdata_int[7]), .ip2(i_ssi_U_dff_tx_mem[103]), 
        .s(n5286), .op(n4473) );
  nand2_1 U11765 ( .ip1(n10400), .ip2(i_ssi_U_dff_tx_mem[87]), .op(n10358) );
  nand2_1 U11766 ( .ip1(n10401), .ip2(i_ssi_U_dff_tx_mem[103]), .op(n10357) );
  nand2_1 U11767 ( .ip1(n10402), .ip2(i_ssi_U_dff_tx_mem[55]), .op(n10356) );
  nand2_1 U11768 ( .ip1(n10389), .ip2(i_ssi_U_dff_tx_mem[39]), .op(n10355) );
  nand2_1 U11769 ( .ip1(n10407), .ip2(i_ssi_U_dff_tx_mem[119]), .op(n10362) );
  nand2_1 U11770 ( .ip1(n10408), .ip2(i_ssi_U_dff_tx_mem[23]), .op(n10361) );
  nand2_1 U11771 ( .ip1(n5609), .ip2(i_ssi_U_dff_tx_mem[7]), .op(n10360) );
  nand2_1 U11772 ( .ip1(n5252), .ip2(i_ssi_U_dff_tx_mem[71]), .op(n10359) );
  or2_1 U11773 ( .ip1(n10364), .ip2(n10363), .op(n10682) );
  mux2_1 U11774 ( .ip1(n10682), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[7]), 
        .s(n10377), .op(n4413) );
  mux2_1 U11775 ( .ip1(i_apb_pwdata_int[6]), .ip2(i_ssi_U_dff_tx_mem[118]), 
        .s(n5254), .op(n4458) );
  mux2_1 U11776 ( .ip1(i_apb_pwdata_int[6]), .ip2(i_ssi_U_dff_tx_mem[38]), .s(
        n10365), .op(n4538) );
  mux2_1 U11777 ( .ip1(i_apb_pwdata_int[6]), .ip2(i_ssi_U_dff_tx_mem[86]), .s(
        n5255), .op(n4490) );
  mux2_1 U11778 ( .ip1(i_apb_pwdata_int[6]), .ip2(i_ssi_U_dff_tx_mem[54]), .s(
        n5253), .op(n4522) );
  mux2_1 U11779 ( .ip1(i_apb_pwdata_int[6]), .ip2(i_ssi_U_dff_tx_mem[22]), .s(
        n5256), .op(n4554) );
  mux2_1 U11780 ( .ip1(i_apb_pwdata_int[6]), .ip2(i_ssi_U_dff_tx_mem[102]), 
        .s(n5286), .op(n4474) );
  nand2_1 U11781 ( .ip1(n10400), .ip2(i_ssi_U_dff_tx_mem[86]), .op(n10369) );
  nand2_1 U11782 ( .ip1(n10401), .ip2(i_ssi_U_dff_tx_mem[102]), .op(n10368) );
  nand2_1 U11783 ( .ip1(n10402), .ip2(i_ssi_U_dff_tx_mem[54]), .op(n10367) );
  nand2_1 U11784 ( .ip1(n10389), .ip2(i_ssi_U_dff_tx_mem[38]), .op(n10366) );
  nand2_1 U11785 ( .ip1(n10407), .ip2(i_ssi_U_dff_tx_mem[118]), .op(n10374) );
  nand2_1 U11786 ( .ip1(n10370), .ip2(i_ssi_U_dff_tx_mem[22]), .op(n10373) );
  nand2_1 U11787 ( .ip1(n5609), .ip2(i_ssi_U_dff_tx_mem[6]), .op(n10372) );
  nand2_1 U11788 ( .ip1(n5252), .ip2(i_ssi_U_dff_tx_mem[70]), .op(n10371) );
  or2_1 U11789 ( .ip1(n10376), .ip2(n10375), .op(n10688) );
  mux2_1 U11790 ( .ip1(n10688), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[6]), 
        .s(n10377), .op(n4414) );
  mux2_1 U11791 ( .ip1(i_ssi_U_dff_tx_mem[69]), .ip2(i_apb_pwdata_int[5]), .s(
        n10354), .op(n4507) );
  mux2_1 U11792 ( .ip1(i_apb_pwdata_int[5]), .ip2(i_ssi_U_dff_tx_mem[117]), 
        .s(n5254), .op(n4459) );
  mux2_1 U11793 ( .ip1(i_ssi_U_dff_tx_mem[5]), .ip2(i_apb_pwdata_int[5]), .s(
        n5608), .op(n4571) );
  mux2_1 U11794 ( .ip1(i_apb_pwdata_int[5]), .ip2(i_ssi_U_dff_tx_mem[37]), .s(
        n10365), .op(n4539) );
  mux2_1 U11795 ( .ip1(i_apb_pwdata_int[5]), .ip2(i_ssi_U_dff_tx_mem[85]), .s(
        n5255), .op(n4491) );
  mux2_1 U11796 ( .ip1(i_apb_pwdata_int[5]), .ip2(i_ssi_U_dff_tx_mem[53]), .s(
        n5253), .op(n4523) );
  mux2_1 U11797 ( .ip1(i_apb_pwdata_int[5]), .ip2(i_ssi_U_dff_tx_mem[21]), .s(
        n5256), .op(n4555) );
  mux2_1 U11798 ( .ip1(i_apb_pwdata_int[5]), .ip2(i_ssi_U_dff_tx_mem[101]), 
        .s(n5286), .op(n4475) );
  nand2_1 U11799 ( .ip1(n10400), .ip2(i_ssi_U_dff_tx_mem[85]), .op(n10381) );
  nand2_1 U11800 ( .ip1(n10401), .ip2(i_ssi_U_dff_tx_mem[101]), .op(n10380) );
  nand2_1 U11801 ( .ip1(n10402), .ip2(i_ssi_U_dff_tx_mem[53]), .op(n10379) );
  nand2_1 U11802 ( .ip1(n10389), .ip2(i_ssi_U_dff_tx_mem[37]), .op(n10378) );
  nand2_1 U11803 ( .ip1(n10407), .ip2(i_ssi_U_dff_tx_mem[117]), .op(n10385) );
  nand2_1 U11804 ( .ip1(n10408), .ip2(i_ssi_U_dff_tx_mem[21]), .op(n10384) );
  nand2_1 U11805 ( .ip1(n5609), .ip2(i_ssi_U_dff_tx_mem[5]), .op(n10383) );
  nand2_1 U11806 ( .ip1(n5252), .ip2(i_ssi_U_dff_tx_mem[69]), .op(n10382) );
  nor2_1 U11807 ( .ip1(n10387), .ip2(n10386), .op(n10679) );
  inv_1 U11808 ( .ip(n10679), .op(n10388) );
  mux2_1 U11809 ( .ip1(n10388), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[5]), 
        .s(n10377), .op(n4415) );
  mux2_1 U11810 ( .ip1(i_apb_pwdata_int[4]), .ip2(i_ssi_U_dff_tx_mem[116]), 
        .s(n5254), .op(n4460) );
  mux2_1 U11811 ( .ip1(i_apb_pwdata_int[4]), .ip2(i_ssi_U_dff_tx_mem[36]), .s(
        n10365), .op(n4540) );
  mux2_1 U11812 ( .ip1(i_apb_pwdata_int[4]), .ip2(i_ssi_U_dff_tx_mem[84]), .s(
        n5255), .op(n4492) );
  mux2_1 U11813 ( .ip1(i_apb_pwdata_int[4]), .ip2(i_ssi_U_dff_tx_mem[52]), .s(
        n5253), .op(n4524) );
  mux2_1 U11814 ( .ip1(i_apb_pwdata_int[4]), .ip2(i_ssi_U_dff_tx_mem[20]), .s(
        n5256), .op(n4556) );
  mux2_1 U11815 ( .ip1(i_apb_pwdata_int[4]), .ip2(i_ssi_U_dff_tx_mem[100]), 
        .s(n5286), .op(n4476) );
  nand2_1 U11816 ( .ip1(n10400), .ip2(i_ssi_U_dff_tx_mem[84]), .op(n10393) );
  nand2_1 U11817 ( .ip1(n10401), .ip2(i_ssi_U_dff_tx_mem[100]), .op(n10392) );
  nand2_1 U11818 ( .ip1(n10402), .ip2(i_ssi_U_dff_tx_mem[52]), .op(n10391) );
  nand2_1 U11819 ( .ip1(n10389), .ip2(i_ssi_U_dff_tx_mem[36]), .op(n10390) );
  nand2_1 U11820 ( .ip1(n10407), .ip2(i_ssi_U_dff_tx_mem[116]), .op(n10397) );
  nand2_1 U11821 ( .ip1(n10408), .ip2(i_ssi_U_dff_tx_mem[20]), .op(n10396) );
  nand2_1 U11822 ( .ip1(n5609), .ip2(i_ssi_U_dff_tx_mem[4]), .op(n10395) );
  nand2_1 U11823 ( .ip1(n5252), .ip2(i_ssi_U_dff_tx_mem[68]), .op(n10394) );
  or2_1 U11824 ( .ip1(n10399), .ip2(n10398), .op(n10680) );
  mux2_1 U11825 ( .ip1(n10680), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[4]), 
        .s(n10377), .op(n4416) );
  nand2_1 U11826 ( .ip1(n10400), .ip2(i_ssi_U_dff_tx_mem[83]), .op(n10406) );
  nand2_1 U11827 ( .ip1(n10401), .ip2(i_ssi_U_dff_tx_mem[99]), .op(n10405) );
  nand2_1 U11828 ( .ip1(n10402), .ip2(i_ssi_U_dff_tx_mem[51]), .op(n10404) );
  nand2_1 U11829 ( .ip1(n10389), .ip2(i_ssi_U_dff_tx_mem[35]), .op(n10403) );
  nand2_1 U11830 ( .ip1(n10407), .ip2(i_ssi_U_dff_tx_mem[115]), .op(n10412) );
  nand2_1 U11831 ( .ip1(n10408), .ip2(i_ssi_U_dff_tx_mem[19]), .op(n10411) );
  nand2_1 U11832 ( .ip1(n5609), .ip2(i_ssi_U_dff_tx_mem[3]), .op(n10410) );
  nand2_1 U11833 ( .ip1(n5252), .ip2(i_ssi_U_dff_tx_mem[67]), .op(n10409) );
  or2_1 U11834 ( .ip1(n10414), .ip2(n10413), .op(n10651) );
  mux2_1 U11835 ( .ip1(n10651), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[3]), 
        .s(n10377), .op(n4417) );
  nand2_1 U11836 ( .ip1(n5283), .ip2(n10651), .op(n10436) );
  not_ab_or_c_or_d U11837 ( .ip1(n10422), .ip2(n5288), .ip3(
        i_ssi_U_mstfsm_tx_load_en_int), .ip4(n10421), .op(n10423) );
  inv_1 U11838 ( .ip(n10589), .op(n10425) );
  inv_1 U11839 ( .ip(n10425), .op(n10453) );
  nand2_1 U11840 ( .ip1(n5271), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[3]), 
        .op(n10435) );
  nor2_1 U11841 ( .ip1(i_ssi_U_mstfsm_spi0_control), .ip2(
        i_ssi_U_mstfsm_spi1_control), .op(n10426) );
  nor2_1 U11842 ( .ip1(n10427), .ip2(n10426), .op(n10428) );
  nor2_1 U11843 ( .ip1(n10429), .ip2(n10428), .op(n10431) );
  nor2_1 U11844 ( .ip1(n10431), .ip2(n10430), .op(n10432) );
  nor2_1 U11845 ( .ip1(n10433), .ip2(n10432), .op(n10568) );
  inv_1 U11846 ( .ip(n10568), .op(n10577) );
  nand2_1 U11847 ( .ip1(n10577), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[2]), .op(n10434) );
  nand4_1 U11848 ( .ip1(n10436), .ip2(n10416), .ip3(n10435), .ip4(n10434), 
        .op(n10448) );
  inv_1 U11849 ( .ip(i_ssi_dfs[0]), .op(n11471) );
  nor2_1 U11850 ( .ip1(n5342), .ip2(n5341), .op(n10439) );
  nand2_1 U11851 ( .ip1(n10488), .ip2(n10683), .op(n10529) );
  inv_1 U11852 ( .ip(n10529), .op(n10446) );
  inv_1 U11853 ( .ip(n5327), .op(n10860) );
  nor2_1 U11854 ( .ip1(n5416), .ip2(n5514), .op(n10444) );
  nand2_1 U11855 ( .ip1(n10444), .ip2(n5373), .op(n10445) );
  mux2_1 U11856 ( .ip1(n10448), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[3]), .s(n10447), .op(n4400) );
  nand2_1 U11857 ( .ip1(n5283), .ip2(n10680), .op(n10451) );
  nand2_1 U11858 ( .ip1(n5271), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[4]), 
        .op(n10450) );
  nand2_1 U11859 ( .ip1(n10577), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[3]), .op(n10449) );
  nand4_1 U11860 ( .ip1(n10451), .ip2(n10416), .ip3(n10450), .ip4(n10449), 
        .op(n10452) );
  mux2_1 U11861 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[4]), .ip2(
        n10452), .s(n10469), .op(n4399) );
  or2_1 U11862 ( .ip1(n10679), .ip2(n10440), .op(n10456) );
  nand2_1 U11863 ( .ip1(n5271), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[5]), 
        .op(n10455) );
  nand2_1 U11864 ( .ip1(n10577), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[4]), .op(n10454) );
  nand4_1 U11865 ( .ip1(n10456), .ip2(n10416), .ip3(n10455), .ip4(n10454), 
        .op(n10463) );
  inv_1 U11866 ( .ip(n10488), .op(n10567) );
  nor3_1 U11867 ( .ip1(n5357), .ip2(n10681), .ip3(n10567), .op(n10461) );
  nand2_1 U11868 ( .ip1(n5357), .ip2(n10457), .op(n10460) );
  nand2_1 U11869 ( .ip1(n10577), .ip2(n5324), .op(n10458) );
  nor2_1 U11870 ( .ip1(n10516), .ip2(n10461), .op(n10462) );
  mux2_1 U11871 ( .ip1(n10463), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[5]), .s(n10462), .op(n4398) );
  nand2_1 U11872 ( .ip1(n5283), .ip2(n10688), .op(n10466) );
  nand2_1 U11873 ( .ip1(n5271), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[6]), 
        .op(n10465) );
  nand2_1 U11874 ( .ip1(n10577), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[5]), .op(n10464) );
  nand4_1 U11875 ( .ip1(n10466), .ip2(n10416), .ip3(n10465), .ip4(n10464), 
        .op(n10472) );
  nor2_1 U11876 ( .ip1(n10540), .ip2(n5324), .op(n10468) );
  nand2_1 U11877 ( .ip1(n10530), .ip2(n10468), .op(n10470) );
  nand2_1 U11878 ( .ip1(n10470), .ip2(n10469), .op(n10471) );
  mux2_1 U11879 ( .ip1(n10472), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[6]), .s(n10471), .op(n4397) );
  nand2_1 U11880 ( .ip1(n5283), .ip2(n10682), .op(n10475) );
  nand2_1 U11881 ( .ip1(n5271), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[7]), 
        .op(n10474) );
  nand2_1 U11882 ( .ip1(n10577), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[6]), .op(n10473) );
  nand4_1 U11883 ( .ip1(n10475), .ip2(n10416), .ip3(n10474), .ip4(n10473), 
        .op(n10478) );
  nor2_1 U11884 ( .ip1(n5357), .ip2(n10529), .op(n10476) );
  nor2_1 U11885 ( .ip1(n10516), .ip2(n10476), .op(n10477) );
  mux2_1 U11886 ( .ip1(n10478), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[7]), .s(n10477), .op(n4396) );
  nand2_1 U11887 ( .ip1(n5283), .ip2(n10662), .op(n10482) );
  nand2_1 U11888 ( .ip1(n5271), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[8]), 
        .op(n10481) );
  nand2_1 U11889 ( .ip1(n10577), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[7]), .op(n10480) );
  nand4_1 U11890 ( .ip1(n10482), .ip2(n10416), .ip3(n10481), .ip4(n10480), 
        .op(n10483) );
  nand2_1 U11891 ( .ip1(n5283), .ip2(n10658), .op(n10486) );
  nand2_1 U11892 ( .ip1(n5271), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[9]), 
        .op(n10485) );
  nand2_1 U11893 ( .ip1(n10577), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[8]), .op(n10484) );
  nand4_1 U11894 ( .ip1(n10486), .ip2(n10485), .ip3(n10416), .ip4(n10484), 
        .op(n10490) );
  inv_1 U11895 ( .ip(n10502), .op(n10487) );
  nand3_1 U11896 ( .ip1(n10551), .ip2(n5324), .ip3(n5486), .op(n10489) );
  nand2_1 U11897 ( .ip1(n5283), .ip2(n10661), .op(n10493) );
  nand2_1 U11898 ( .ip1(n5271), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[10]), 
        .op(n10492) );
  nand2_1 U11899 ( .ip1(n10577), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[9]), .op(n10491) );
  nand4_1 U11900 ( .ip1(n10493), .ip2(n10416), .ip3(n10492), .ip4(n10491), 
        .op(n10495) );
  mux2_1 U11901 ( .ip1(n10495), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[10]), .s(n10494), .op(n4393)
         );
  nand2_1 U11902 ( .ip1(n5283), .ip2(n10659), .op(n10498) );
  nand2_1 U11903 ( .ip1(n5271), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[11]), 
        .op(n10497) );
  nand2_1 U11904 ( .ip1(n10577), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[10]), .op(n10496) );
  nand4_1 U11905 ( .ip1(n10498), .ip2(n10416), .ip3(n10497), .ip4(n10496), 
        .op(n10507) );
  nor2_1 U11906 ( .ip1(n5438), .ip2(n10529), .op(n10505) );
  nand2_1 U11907 ( .ip1(n5357), .ip2(n10577), .op(n10499) );
  nor2_1 U11908 ( .ip1(n10499), .ip2(n5373), .op(n10500) );
  nand2_1 U11909 ( .ip1(n10500), .ip2(n10502), .op(n10504) );
  nand2_1 U11910 ( .ip1(n10501), .ip2(n10502), .op(n10503) );
  mux2_1 U11911 ( .ip1(n10507), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[11]), .s(n10506), .op(n4392)
         );
  nand2_1 U11912 ( .ip1(n5283), .ip2(n10616), .op(n10510) );
  nand2_1 U11913 ( .ip1(n5271), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[12]), 
        .op(n10509) );
  nand2_1 U11914 ( .ip1(n10577), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[11]), .op(n10508) );
  nand4_1 U11915 ( .ip1(n10510), .ip2(n10416), .ip3(n10509), .ip4(n10508), 
        .op(n10511) );
  mux2_1 U11916 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[12]), .ip2(
        n10511), .s(n5437), .op(n4391) );
  nand2_1 U11917 ( .ip1(n5283), .ip2(n10622), .op(n10514) );
  nand2_1 U11918 ( .ip1(n5271), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[13]), 
        .op(n10513) );
  nand2_1 U11919 ( .ip1(n10577), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[12]), .op(n10512) );
  nand4_1 U11920 ( .ip1(n10514), .ip2(n10416), .ip3(n10513), .ip4(n10512), 
        .op(n10519) );
  nand2_1 U11921 ( .ip1(n5281), .ip2(n5373), .op(n10515) );
  nand2_1 U11922 ( .ip1(n10530), .ip2(n10515), .op(n10517) );
  nand2_1 U11923 ( .ip1(n10516), .ip2(n10517), .op(n10518) );
  mux2_1 U11924 ( .ip1(n10519), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[13]), .s(n10518), .op(n4390)
         );
  nand2_1 U11925 ( .ip1(n5283), .ip2(n10614), .op(n10522) );
  nand2_1 U11926 ( .ip1(n5271), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[14]), 
        .op(n10521) );
  nand2_1 U11927 ( .ip1(n10577), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[13]), .op(n10520) );
  nand4_1 U11928 ( .ip1(n10522), .ip2(n10416), .ip3(n10521), .ip4(n10520), 
        .op(n10525) );
  nand2_1 U11929 ( .ip1(n10530), .ip2(n5423), .op(n10523) );
  nand2_1 U11930 ( .ip1(n10523), .ip2(n5436), .op(n10524) );
  mux2_1 U11931 ( .ip1(n10525), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[14]), .s(n10524), .op(n4404)
         );
  nand2_1 U11932 ( .ip1(n5283), .ip2(n10617), .op(n10528) );
  nand2_1 U11933 ( .ip1(n5271), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[15]), 
        .op(n10527) );
  nand2_1 U11934 ( .ip1(n10577), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[14]), .op(n10526) );
  nand4_1 U11935 ( .ip1(n10528), .ip2(n10416), .ip3(n10527), .ip4(n10526), 
        .op(n10533) );
  inv_1 U11936 ( .ip(n5362), .op(n10629) );
  nor2_1 U11937 ( .ip1(n10629), .ip2(n10529), .op(n10532) );
  nor2_1 U11938 ( .ip1(n10567), .ip2(n10530), .op(n10531) );
  nand2_1 U11939 ( .ip1(n10415), .ip2(n10653), .op(n10537) );
  inv_1 U11940 ( .ip(i_ssi_U_shift_U_tx_shifter_tx_buffer[0]), .op(n10534) );
  nor2_1 U11941 ( .ip1(n10534), .ip2(n5358), .op(n10535) );
  nor2_1 U11942 ( .ip1(i_ssi_load_start_bit), .ip2(n10535), .op(n10536) );
  nand2_1 U11943 ( .ip1(n10537), .ip2(n10536), .op(n10552) );
  not_ab_or_c_or_d U11944 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[0]), 
        .ip2(n10567), .ip3(n10577), .ip4(n10552), .op(n10566) );
  nand2_1 U11945 ( .ip1(n10672), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[8]), .op(n10598) );
  nand3_1 U11946 ( .ip1(n10598), .ip2(n10600), .ip3(n10599), .op(n10564) );
  inv_1 U11947 ( .ip(n5347), .op(n10615) );
  inv_1 U11948 ( .ip(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[6]), .op(n10541)
         );
  inv_2 U11949 ( .ip(n10648), .op(n10633) );
  nand2_2 U11950 ( .ip1(n10542), .ip2(n10543), .op(n10544) );
  nor2_1 U11951 ( .ip1(n10587), .ip2(n10615), .op(n10563) );
  nand2_1 U11952 ( .ip1(n5279), .ip2(n5359), .op(n10561) );
  not_ab_or_c_or_d U11953 ( .ip1(n10553), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[15]), .ip3(n5478), .ip4(n10552), .op(n10560) );
  nand2_1 U11954 ( .ip1(n10672), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[11]), .op(n10557) );
  nand2_1 U11955 ( .ip1(n10633), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[3]), .op(n10556) );
  nand2_1 U11956 ( .ip1(n10678), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[7]), .op(n10555) );
  nand2_1 U11957 ( .ip1(n5362), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[15]), .op(n10554) );
  nand4_1 U11958 ( .ip1(n10557), .ip2(n10556), .ip3(n10555), .ip4(n10554), 
        .op(n10558) );
  nand2_1 U11959 ( .ip1(n10660), .ip2(n10558), .op(n10559) );
  nand3_1 U11960 ( .ip1(n10561), .ip2(n10560), .ip3(n10559), .op(n10562) );
  not_ab_or_c_or_d U11961 ( .ip1(n10681), .ip2(n10564), .ip3(n10562), .ip4(
        n10563), .op(n10565) );
  nor2_1 U11962 ( .ip1(n10566), .ip2(n10565), .op(n4403) );
  nand2_1 U11963 ( .ip1(n10567), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[1]), .op(n10573) );
  inv_1 U11964 ( .ip(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[0]), .op(n10569)
         );
  nor2_1 U11965 ( .ip1(n10569), .ip2(n10568), .op(n10570) );
  not_ab_or_c_or_d U11966 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_buffer[1]), 
        .ip2(n5271), .ip3(i_ssi_load_start_bit), .ip4(n10570), .op(n10572) );
  nand2_1 U11967 ( .ip1(n5283), .ip2(n10650), .op(n10571) );
  nand3_1 U11968 ( .ip1(n10573), .ip2(n10572), .ip3(n10571), .op(n4402) );
  nand2_1 U11969 ( .ip1(n5283), .ip2(n10652), .op(n10576) );
  nand2_1 U11970 ( .ip1(n5271), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[2]), 
        .op(n10575) );
  nand2_1 U11971 ( .ip1(n10577), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[1]), .op(n10574) );
  nand4_1 U11972 ( .ip1(n10576), .ip2(n10416), .ip3(n10575), .ip4(n10574), 
        .op(n10582) );
  nand2_1 U11973 ( .ip1(n5279), .ip2(n5393), .op(n10578) );
  nand2_1 U11974 ( .ip1(n10578), .ip2(n10577), .op(n10580) );
  nand2_1 U11975 ( .ip1(n10580), .ip2(n10579), .op(n10581) );
  mux2_1 U11976 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[2]), .ip2(
        n10582), .s(n10581), .op(n4401) );
  inv_1 U11977 ( .ip(i_ssi_U_shift_U_tx_shifter_load_start_bit_ir), .op(n10583) );
  nand2_1 U11978 ( .ip1(n5358), .ip2(n10583), .op(n10584) );
  inv_1 U11979 ( .ip(n10584), .op(n10585) );
  nand2_1 U11980 ( .ip1(n10591), .ip2(n10585), .op(n10639) );
  nor2_1 U11981 ( .ip1(n10639), .ip2(n10615), .op(n10608) );
  inv_1 U11982 ( .ip(n10639), .op(n10586) );
  nand2_1 U11983 ( .ip1(n10683), .ip2(n10586), .op(n10588) );
  nor2_1 U11984 ( .ip1(n5322), .ip2(
        i_ssi_U_shift_U_tx_shifter_load_start_bit_ir), .op(n10673) );
  inv_1 U11985 ( .ip(n10673), .op(n10630) );
  nor2_1 U11986 ( .ip1(n10630), .ip2(n5514), .op(n10596) );
  inv_1 U11987 ( .ip(i_ssi_txd), .op(n10592) );
  nor4_1 U11988 ( .ip1(i_ssi_U_shift_U_tx_shifter_load_start_bit_ir), .ip2(
        n10592), .ip3(n10591), .ip4(n10415), .op(n10594) );
  and2_1 U11989 ( .ip1(i_ssi_U_shift_U_tx_shifter_tx_shift_reg[15]), .ip2(
        i_ssi_U_shift_U_tx_shifter_load_start_bit_ir), .op(n10593) );
  not_ab_or_c_or_d U11990 ( .ip1(n10596), .ip2(n10595), .ip3(n10594), .ip4(
        n10593), .op(n10604) );
  nand2_1 U11991 ( .ip1(n5393), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[0]), .op(n10597) );
  nand4_1 U11992 ( .ip1(n10600), .ip2(n10598), .ip3(n10599), .ip4(n10597), 
        .op(n10602) );
  nor2_1 U11993 ( .ip1(n10639), .ip2(n5397), .op(n10601) );
  nand2_1 U11994 ( .ip1(n10601), .ip2(n10602), .op(n10603) );
  nand2_1 U11995 ( .ip1(n10604), .ip2(n10603), .op(n10605) );
  not_ab_or_c_or_d U11996 ( .ip1(n10608), .ip2(n10607), .ip3(n10605), .ip4(
        n10606), .op(n10698) );
  nor2_1 U11997 ( .ip1(n10630), .ip2(n5337), .op(n10647) );
  nand2_1 U11998 ( .ip1(n5279), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[5]), 
        .op(n10613) );
  nand2_1 U11999 ( .ip1(n10660), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[7]), 
        .op(n10612) );
  nand2_1 U12000 ( .ip1(n5347), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[6]), 
        .op(n10611) );
  nand2_1 U12001 ( .ip1(n10681), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[4]), 
        .op(n10610) );
  nand4_1 U12002 ( .ip1(n10613), .ip2(n10612), .ip3(n10611), .ip4(n10610), 
        .op(n10646) );
  nand2_1 U12003 ( .ip1(n5374), .ip2(n10677), .op(n10624) );
  nand2_1 U12004 ( .ip1(n10681), .ip2(n10616), .op(n10619) );
  nand2_1 U12005 ( .ip1(n5422), .ip2(n10617), .op(n10618) );
  nand2_1 U12006 ( .ip1(n10619), .ip2(n10618), .op(n10620) );
  not_ab_or_c_or_d U12007 ( .ip1(n5279), .ip2(n10622), .ip3(n10621), .ip4(
        n10620), .op(n10623) );
  nor2_1 U12008 ( .ip1(n10624), .ip2(n10623), .op(n10645) );
  nand2_1 U12009 ( .ip1(n5279), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[13]), 
        .op(n10628) );
  nand2_1 U12010 ( .ip1(n10681), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[12]), .op(n10625) );
  nor2_1 U12011 ( .ip1(n10630), .ip2(n10629), .op(n10631) );
  nand2_1 U12012 ( .ip1(n10631), .ip2(n10632), .op(n10643) );
  nand2_1 U12013 ( .ip1(n10672), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[7]), .op(n10637) );
  nand2_1 U12014 ( .ip1(n10633), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[14]), .op(n10636) );
  nand2_1 U12015 ( .ip1(n10678), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[3]), .op(n10635) );
  nand2_1 U12016 ( .ip1(n5362), .ip2(
        i_ssi_U_shift_U_tx_shifter_tx_shift_reg[11]), .op(n10634) );
  nand4_1 U12017 ( .ip1(n10637), .ip2(n10636), .ip3(n10635), .ip4(n10634), 
        .op(n10641) );
  nor2_1 U12018 ( .ip1(n10639), .ip2(n5373), .op(n10640) );
  nand2_1 U12019 ( .ip1(n10640), .ip2(n10641), .op(n10642) );
  nand2_1 U12020 ( .ip1(n10643), .ip2(n10642), .op(n10644) );
  not_ab_or_c_or_d U12021 ( .ip1(n10647), .ip2(n10646), .ip3(n10644), .ip4(
        n10645), .op(n10697) );
  inv_1 U12022 ( .ip(n10677), .op(n10649) );
  nor2_1 U12023 ( .ip1(n10649), .ip2(n5514), .op(n10695) );
  nand2_1 U12024 ( .ip1(n5279), .ip2(n10650), .op(n10657) );
  nand2_1 U12025 ( .ip1(n10660), .ip2(n10651), .op(n10656) );
  nand2_1 U12026 ( .ip1(n5347), .ip2(n10652), .op(n10655) );
  nand2_1 U12027 ( .ip1(n10681), .ip2(n10653), .op(n10654) );
  nand4_1 U12028 ( .ip1(n10657), .ip2(n10656), .ip3(n10655), .ip4(n10654), 
        .op(n10694) );
  nand2_1 U12029 ( .ip1(n5279), .ip2(n10658), .op(n10666) );
  nand2_1 U12030 ( .ip1(n5422), .ip2(n10659), .op(n10665) );
  nand3_1 U12031 ( .ip1(n10672), .ip2(n10677), .ip3(n10667), .op(n10676) );
  nand2_1 U12032 ( .ip1(n5279), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[9]), 
        .op(n10671) );
  nand2_1 U12033 ( .ip1(n10683), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[11]), .op(n10670) );
  nand2_1 U12034 ( .ip1(n10689), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[10]), .op(n10669) );
  nand2_1 U12035 ( .ip1(n10681), .ip2(i_ssi_U_shift_U_tx_shifter_tx_buffer[8]), 
        .op(n10668) );
  nand4_1 U12036 ( .ip1(n10669), .ip2(n10671), .ip3(n10670), .ip4(n10668), 
        .op(n10674) );
  nand2_1 U12037 ( .ip1(n10676), .ip2(n10675), .op(n10693) );
  nand2_1 U12038 ( .ip1(n10678), .ip2(n10677), .op(n10691) );
  nor2_1 U12039 ( .ip1(n10679), .ip2(n5397), .op(n10687) );
  nand2_1 U12040 ( .ip1(n10681), .ip2(n10680), .op(n10685) );
  nand2_1 U12041 ( .ip1(n10684), .ip2(n10685), .op(n10686) );
  not_ab_or_c_or_d U12042 ( .ip1(n5347), .ip2(n10688), .ip3(n10687), .ip4(
        n10686), .op(n10690) );
  nor2_1 U12043 ( .ip1(n10691), .ip2(n10690), .op(n10692) );
  not_ab_or_c_or_d U12044 ( .ip1(n10695), .ip2(n10694), .ip3(n10693), .ip4(
        n10692), .op(n10696) );
  nand3_1 U12045 ( .ip1(n10696), .ip2(n10698), .ip3(n10697), .op(n4388) );
  mux2_1 U12046 ( .ip1(i_ssi_rxd), .ip2(i_ssi_txd), .s(i_ssi_ctrlr0[11]), .op(
        n10706) );
  inv_1 U12047 ( .ip(n10699), .op(n10700) );
  nand2_1 U12048 ( .ip1(n10701), .ip2(n10700), .op(n10702) );
  nand2_1 U12049 ( .ip1(n10702), .ip2(i_ssi_sclk_re), .op(n10704) );
  nand2_1 U12050 ( .ip1(n10704), .ip2(n10703), .op(n10705) );
  mux2_1 U12051 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[0]), .ip2(
        n10706), .s(n10865), .op(n4387) );
  mux2_1 U12052 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[1]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[0]), .s(n10865), .op(n4386) );
  mux2_1 U12053 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[2]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[1]), .s(n10865), .op(n4385) );
  mux2_1 U12054 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[3]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[2]), .s(n10865), .op(n4384) );
  mux2_1 U12055 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[4]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[3]), .s(n10865), .op(n4383) );
  mux2_1 U12056 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[5]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[4]), .s(n10865), .op(n4382) );
  mux2_1 U12057 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[6]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[5]), .s(n10865), .op(n4381) );
  nor2_1 U12058 ( .ip1(n5351), .ip2(n5453), .op(n10707) );
  nor2_1 U12059 ( .ip1(n10707), .ip2(n10843), .op(n10708) );
  nand2_1 U12060 ( .ip1(n10122), .ip2(n10708), .op(n10858) );
  inv_1 U12061 ( .ip(n10858), .op(n10709) );
  nand2_1 U12062 ( .ip1(n10709), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[6]), .op(n10711) );
  nand2_1 U12063 ( .ip1(n10868), .ip2(i_ssi_rx_push_data[6]), .op(n10710) );
  nand2_1 U12064 ( .ip1(n10711), .ip2(n10710), .op(n4432) );
  inv_1 U12065 ( .ip(i_ssi_rx_full), .op(n10851) );
  nor2_1 U12066 ( .ip1(n10851), .ip2(n6937), .op(n10712) );
  nand2_1 U12067 ( .ip1(n10720), .ip2(i_ssi_U_fifo_U_rx_fifo_wr_addr_at_max), 
        .op(n10714) );
  nand2_1 U12068 ( .ip1(n10714), .ip2(n10759), .op(n10724) );
  inv_1 U12069 ( .ip(n10724), .op(n10719) );
  inv_1 U12070 ( .ip(n10720), .op(n10715) );
  nand2_1 U12071 ( .ip1(n10715), .ip2(i_ssi_rx_wr_addr[0]), .op(n10717) );
  inv_1 U12072 ( .ip(i_ssi_rx_wr_addr[0]), .op(n10716) );
  nand2_1 U12073 ( .ip1(n10720), .ip2(n10716), .op(n10783) );
  nand2_1 U12074 ( .ip1(n10717), .ip2(n10783), .op(n10718) );
  and2_1 U12075 ( .ip1(n10719), .ip2(n10718), .op(n11846) );
  inv_1 U12076 ( .ip(i_ssi_rx_wr_addr[1]), .op(n10780) );
  nand2_1 U12077 ( .ip1(n10720), .ip2(i_ssi_rx_wr_addr[0]), .op(n10781) );
  nor2_1 U12078 ( .ip1(n10780), .ip2(n10781), .op(n10776) );
  not_ab_or_c_or_d U12079 ( .ip1(n10780), .ip2(n10781), .ip3(n10724), .ip4(
        n10776), .op(i_ssi_U_fifo_U_rx_fifo_N42) );
  and2_1 U12080 ( .ip1(i_ssi_rx_wr_addr[1]), .ip2(i_ssi_rx_wr_addr[2]), .op(
        n10774) );
  and2_1 U12081 ( .ip1(n11846), .ip2(n10774), .op(i_ssi_U_fifo_U_rx_fifo_N40)
         );
  inv_1 U12082 ( .ip(i_ssi_rx_wr_addr[2]), .op(n10779) );
  nor2_1 U12083 ( .ip1(n10779), .ip2(n10776), .op(n10722) );
  nor2_1 U12084 ( .ip1(n10722), .ip2(n10721), .op(n10723) );
  nor2_1 U12085 ( .ip1(n10724), .ip2(n10723), .op(i_ssi_U_fifo_U_rx_fifo_N43)
         );
  mux2_1 U12086 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[7]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[6]), .s(n10865), .op(n4380) );
  mux2_1 U12087 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[8]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[7]), .s(n10865), .op(n4379) );
  nand2_1 U12088 ( .ip1(n10122), .ip2(n5453), .op(n10742) );
  inv_1 U12089 ( .ip(n10742), .op(n10733) );
  nand2_1 U12090 ( .ip1(n10733), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[8]), .op(n10726) );
  nand2_1 U12091 ( .ip1(n10868), .ip2(i_ssi_rx_push_data[8]), .op(n10725) );
  nand2_1 U12092 ( .ip1(n10726), .ip2(n10725), .op(n4430) );
  mux2_1 U12093 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[9]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[8]), .s(n10865), .op(n4378) );
  inv_1 U12094 ( .ip(i_ssi_rx_push_data[9]), .op(n10727) );
  nor2_1 U12095 ( .ip1(n10727), .ip2(n10122), .op(n10731) );
  nand2_1 U12096 ( .ip1(n11471), .ip2(n10737), .op(n10831) );
  inv_1 U12097 ( .ip(n10831), .op(n10729) );
  inv_1 U12098 ( .ip(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[9]), .op(n10728)
         );
  not_ab_or_c_or_d U12099 ( .ip1(n10729), .ip2(n10743), .ip3(n10728), .ip4(
        n10742), .op(n10730) );
  or2_1 U12100 ( .ip1(n10731), .ip2(n10730), .op(n4429) );
  mux2_1 U12101 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[10]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[9]), .s(n10865), .op(n4377) );
  nand2_1 U12102 ( .ip1(n10737), .ip2(n10743), .op(n10732) );
  nand3_1 U12103 ( .ip1(n10733), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[10]), .ip3(n10732), .op(n10735) );
  nand2_1 U12104 ( .ip1(n10868), .ip2(i_ssi_rx_push_data[10]), .op(n10734) );
  nand2_1 U12105 ( .ip1(n10735), .ip2(n10734), .op(n4428) );
  mux2_1 U12106 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[11]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[10]), .s(n10865), .op(n4376)
         );
  inv_1 U12107 ( .ip(i_ssi_rx_push_data[11]), .op(n10736) );
  nor2_1 U12108 ( .ip1(n10736), .ip2(n10122), .op(n10741) );
  nor2_1 U12109 ( .ip1(n10737), .ip2(n11471), .op(n10866) );
  inv_1 U12110 ( .ip(n10866), .op(n10739) );
  inv_1 U12111 ( .ip(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[11]), .op(n10738)
         );
  not_ab_or_c_or_d U12112 ( .ip1(n10743), .ip2(n10739), .ip3(n10738), .ip4(
        n10742), .op(n10740) );
  or2_1 U12113 ( .ip1(n10741), .ip2(n10740), .op(n4427) );
  mux2_1 U12114 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[12]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[11]), .s(n10865), .op(n4375)
         );
  nor2_1 U12115 ( .ip1(n10743), .ip2(n10742), .op(n10867) );
  nand2_1 U12116 ( .ip1(n10867), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[12]), .op(n10745) );
  nand2_1 U12117 ( .ip1(n10868), .ip2(i_ssi_rx_push_data[12]), .op(n10744) );
  nand2_1 U12118 ( .ip1(n10745), .ip2(n10744), .op(n4426) );
  mux2_1 U12119 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[13]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[12]), .s(n10865), .op(n4374)
         );
  nand3_1 U12120 ( .ip1(n10867), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[13]), .ip3(n10831), .op(n10747) );
  nand2_1 U12121 ( .ip1(n10868), .ip2(i_ssi_rx_push_data[13]), .op(n10746) );
  nand2_1 U12122 ( .ip1(n10747), .ip2(n10746), .op(n4425) );
  mux2_1 U12123 ( .ip1(i_ssi_imr[2]), .ip2(i_apb_pwdata_int[2]), .s(n10846), 
        .op(n4641) );
  nand2_1 U12124 ( .ip1(n11837), .ip2(i_ssi_rx_full), .op(n10750) );
  not_ab_or_c_or_d U12125 ( .ip1(n6688), .ip2(n10750), .ip3(n10749), .ip4(
        n10748), .op(i_ssi_U_fifo_U_rx_fifo_N38) );
  inv_1 U12126 ( .ip(i_ssi_U_fifo_rx_error_ir), .op(n10751) );
  inv_1 U12127 ( .ip(i_ssi_U_fifo_rx_pop_dly), .op(n10767) );
  nor3_1 U12128 ( .ip1(i_ssi_U_fifo_U_rx_fifo_empty_n), .ip2(n10751), .ip3(
        n10767), .op(n10756) );
  inv_1 U12129 ( .ip(i_ssi_risr[2]), .op(n10754) );
  nor4_1 U12130 ( .ip1(i_ssi_reg_addr[2]), .ip2(i_ssi_reg_addr[0]), .ip3(
        n10752), .ip4(n11663), .op(n10753) );
  nor2_1 U12131 ( .ip1(n10754), .ip2(n10753), .op(n10755) );
  nor2_1 U12132 ( .ip1(n10756), .ip2(n10755), .op(n10757) );
  nor2_1 U12133 ( .ip1(n5291), .ip2(n10757), .op(n4442) );
  nand2_1 U12134 ( .ip1(i_ssi_risr[2]), .ip2(i_ssi_imr[2]), .op(
        i_ssi_ssi_rxu_intr_n) );
  mux2_1 U12135 ( .ip1(i_ssi_imr[1]), .ip2(i_apb_pwdata_int[1]), .s(n10846), 
        .op(n4642) );
  and3_1 U12136 ( .ip1(n10759), .ip2(n10758), .ip3(i_ssi_tx_full), .op(
        i_ssi_U_fifo_U_tx_fifo_N38) );
  nand2_1 U12137 ( .ip1(n11482), .ip2(n10785), .op(n11456) );
  nand2_1 U12138 ( .ip1(n11456), .ip2(n10760), .op(n10761) );
  nand2_1 U12139 ( .ip1(n6687), .ip2(n10761), .op(n10762) );
  nand2_1 U12140 ( .ip1(n10762), .ip2(i_ssi_risr[1]), .op(n10765) );
  inv_1 U12141 ( .ip(i_ssi_U_fifo_tx_pop_sync_dly), .op(n10763) );
  nand3_1 U12142 ( .ip1(n10763), .ip2(i_ssi_U_fifo_tx_error_ir), .ip3(
        i_ssi_U_fifo_tx_push_dly), .op(n10764) );
  nand2_1 U12143 ( .ip1(n10765), .ip2(n10764), .op(n10766) );
  and2_1 U12144 ( .ip1(n10766), .ip2(n10802), .op(n4577) );
  and2_1 U12145 ( .ip1(i_ssi_imr[1]), .ip2(i_ssi_risr[1]), .op(n11460) );
  inv_1 U12146 ( .ip(n11460), .op(i_ssi_ssi_txo_intr_n) );
  mux2_1 U12147 ( .ip1(i_ssi_imr[3]), .ip2(i_apb_pwdata_int[3]), .s(n10846), 
        .op(n4640) );
  and3_1 U12148 ( .ip1(n10767), .ip2(i_ssi_U_fifo_rx_error_ir), .ip3(
        i_ssi_U_fifo_rx_push_sync_dly), .op(n10772) );
  inv_1 U12149 ( .ip(i_ssi_risr[3]), .op(n11605) );
  nor2_1 U12150 ( .ip1(n11463), .ip2(n11484), .op(n10768) );
  nor2_1 U12151 ( .ip1(n10768), .ip2(n11467), .op(n10769) );
  nor2_1 U12152 ( .ip1(n10769), .ip2(n11663), .op(n10770) );
  nor2_1 U12153 ( .ip1(n11605), .ip2(n10770), .op(n10771) );
  nor2_1 U12154 ( .ip1(n10772), .ip2(n10771), .op(n10773) );
  nor2_1 U12155 ( .ip1(n5291), .ip2(n10773), .op(n4443) );
  nand2_1 U12156 ( .ip1(i_ssi_imr[3]), .ip2(i_ssi_risr[3]), .op(
        i_ssi_ssi_rxo_intr_n) );
  mux2_1 U12157 ( .ip1(i_ssi_rx_push_data[0]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[0]), .s(n10122), .op(n4371) );
  inv_1 U12158 ( .ip(n10774), .op(n10775) );
  or2_1 U12159 ( .ip1(n10775), .ip2(n10783), .op(n11452) );
  mux2_1 U12160 ( .ip1(i_ssi_rx_push_data[0]), .ip2(i_ssi_U_dff_rx_mem[16]), 
        .s(n11452), .op(n4369) );
  nand2_1 U12161 ( .ip1(n10780), .ip2(i_ssi_rx_wr_addr[2]), .op(n10784) );
  mux2_1 U12162 ( .ip1(i_ssi_U_dff_rx_mem[32]), .ip2(i_ssi_rx_push_data[0]), 
        .s(n5610), .op(n4368) );
  mux2_1 U12163 ( .ip1(i_ssi_U_dff_rx_mem[0]), .ip2(i_ssi_rx_push_data[0]), 
        .s(n10777), .op(n4370) );
  nand2_1 U12164 ( .ip1(n10779), .ip2(i_ssi_rx_wr_addr[1]), .op(n10778) );
  or2_1 U12165 ( .ip1(n10778), .ip2(n10783), .op(n11454) );
  mux2_1 U12166 ( .ip1(i_ssi_rx_push_data[0]), .ip2(i_ssi_U_dff_rx_mem[80]), 
        .s(n11454), .op(n4365) );
  nand2_1 U12167 ( .ip1(n10780), .ip2(n10779), .op(n10782) );
  or2_1 U12168 ( .ip1(n10782), .ip2(n10783), .op(n11455) );
  mux2_1 U12169 ( .ip1(i_ssi_rx_push_data[0]), .ip2(i_ssi_U_dff_rx_mem[112]), 
        .s(n11455), .op(n4363) );
  mux2_1 U12170 ( .ip1(i_ssi_U_dff_rx_mem[96]), .ip2(i_ssi_rx_push_data[0]), 
        .s(n5611), .op(n4364) );
  or2_1 U12171 ( .ip1(n10784), .ip2(n10783), .op(n11453) );
  mux2_1 U12172 ( .ip1(i_ssi_rx_push_data[0]), .ip2(i_ssi_U_dff_rx_mem[48]), 
        .s(n11453), .op(n4367) );
  mux2_1 U12173 ( .ip1(i_ssi_U_dff_rx_mem[64]), .ip2(i_ssi_rx_push_data[0]), 
        .s(n10721), .op(n4366) );
  mux2_1 U12174 ( .ip1(i_ssi_imr[0]), .ip2(i_apb_pwdata_int[0]), .s(n10846), 
        .op(n4643) );
  nand2_1 U12175 ( .ip1(n11469), .ip2(n10785), .op(n11527) );
  inv_1 U12176 ( .ip(n11527), .op(n11547) );
  nand2_1 U12177 ( .ip1(n11547), .ip2(n10786), .op(n11451) );
  mux2_1 U12178 ( .ip1(i_apb_pwdata_int[1]), .ip2(i_ssi_txftlr[1]), .s(n11451), 
        .op(n4633) );
  mux2_1 U12179 ( .ip1(i_apb_pwdata_int[0]), .ip2(i_ssi_txftlr[0]), .s(n11451), 
        .op(n4634) );
  nor2_1 U12180 ( .ip1(i_ssi_txftlr[1]), .ip2(i_ssi_txftlr[2]), .op(n10788) );
  or2_1 U12181 ( .ip1(n10788), .ip2(n10787), .op(n10789) );
  nand2_1 U12182 ( .ip1(n10790), .ip2(n10789), .op(n10800) );
  nand2_1 U12183 ( .ip1(n10791), .ip2(i_ssi_txftlr[2]), .op(n10794) );
  nand2_1 U12184 ( .ip1(n10795), .ip2(i_ssi_txftlr[1]), .op(n10793) );
  inv_1 U12185 ( .ip(i_ssi_txftlr[0]), .op(n10792) );
  nand4_1 U12186 ( .ip1(n10794), .ip2(n11853), .ip3(n10793), .ip4(n10792), 
        .op(n10799) );
  or2_1 U12187 ( .ip1(i_ssi_txftlr[1]), .ip2(n10795), .op(n10796) );
  nand2_1 U12188 ( .ip1(n10796), .ip2(i_ssi_txftlr[2]), .op(n10797) );
  nand2_1 U12189 ( .ip1(n10797), .ip2(n11852), .op(n10798) );
  nand3_1 U12190 ( .ip1(n10800), .ip2(n10799), .ip3(n10798), .op(
        i_ssi_U_fifo_U_tx_fifo_N34) );
  inv_1 U12191 ( .ip(i_ssi_U_fifo_U_tx_fifo_almost_empty_n), .op(n10801) );
  nand2_1 U12192 ( .ip1(i_ssi_imr[0]), .ip2(i_ssi_risr[0]), .op(
        i_ssi_ssi_txe_intr_n) );
  nor2_1 U12193 ( .ip1(i_ssi_U_regfile_rxflr[3]), .ip2(n5291), .op(n10804) );
  nand2_1 U12194 ( .ip1(n11837), .ip2(n10804), .op(n10805) );
  nor2_1 U12195 ( .ip1(n10805), .ip2(n6937), .op(n10828) );
  nor2_1 U12196 ( .ip1(n5291), .ip2(n10828), .op(n10809) );
  nor2_1 U12197 ( .ip1(i_ssi_U_regfile_rxflr[3]), .ip2(
        i_ssi_U_regfile_rxflr[2]), .op(n10806) );
  nor2_1 U12198 ( .ip1(i_ssi_U_regfile_rxflr[0]), .ip2(
        i_ssi_U_regfile_rxflr[1]), .op(n10812) );
  not_ab_or_c_or_d U12199 ( .ip1(n10806), .ip2(n10812), .ip3(n5291), .ip4(
        n11837), .op(n10807) );
  and2_1 U12200 ( .ip1(n6937), .ip2(n10807), .op(n10827) );
  inv_1 U12201 ( .ip(i_ssi_U_regfile_rxflr[0]), .op(n11486) );
  nand2_1 U12202 ( .ip1(n10827), .ip2(n11486), .op(n10808) );
  nand2_1 U12203 ( .ip1(n10809), .ip2(n10808), .op(n10811) );
  nand2_1 U12204 ( .ip1(n10828), .ip2(n11486), .op(n10810) );
  nand2_1 U12205 ( .ip1(n10811), .ip2(n10810), .op(n10817) );
  and2_1 U12206 ( .ip1(n10827), .ip2(n10812), .op(n10816) );
  inv_1 U12207 ( .ip(i_ssi_U_regfile_rxflr[1]), .op(n10813) );
  and3_1 U12208 ( .ip1(n10828), .ip2(i_ssi_U_regfile_rxflr[0]), .ip3(n10813), 
        .op(n10814) );
  ab_or_c_or_d U12209 ( .ip1(n10817), .ip2(i_ssi_U_regfile_rxflr[1]), .ip3(
        n10816), .ip4(n10814), .op(n4439) );
  and2_1 U12210 ( .ip1(i_ssi_U_regfile_rxflr[1]), .ip2(
        i_ssi_U_regfile_rxflr[0]), .op(n10815) );
  and2_1 U12211 ( .ip1(n10828), .ip2(n10815), .op(n10824) );
  nor2_1 U12212 ( .ip1(n10824), .ip2(n10816), .op(n10819) );
  mux2_1 U12213 ( .ip1(n10828), .ip2(n10827), .s(i_ssi_U_regfile_rxflr[1]), 
        .op(n10818) );
  nor2_1 U12214 ( .ip1(n10818), .ip2(n10817), .op(n10822) );
  mux2_1 U12215 ( .ip1(n10819), .ip2(n10822), .s(i_ssi_U_regfile_rxflr[2]), 
        .op(n10820) );
  inv_1 U12216 ( .ip(n10820), .op(n4438) );
  nand2_1 U12217 ( .ip1(n10827), .ip2(i_ssi_U_regfile_rxflr[2]), .op(n10821)
         );
  nand2_1 U12218 ( .ip1(n10822), .ip2(n10821), .op(n10823) );
  nand2_1 U12219 ( .ip1(n10823), .ip2(i_ssi_U_regfile_rxflr[3]), .op(n10826)
         );
  nand2_1 U12220 ( .ip1(n10824), .ip2(i_ssi_U_regfile_rxflr[2]), .op(n10825)
         );
  nand2_1 U12221 ( .ip1(n10826), .ip2(n10825), .op(n4441) );
  nor2_1 U12222 ( .ip1(n11486), .ip2(n5291), .op(n10830) );
  nor2_1 U12223 ( .ip1(n10828), .ip2(n10827), .op(n10829) );
  mux2_1 U12224 ( .ip1(n11486), .ip2(n10830), .s(n10829), .op(n4440) );
  inv_1 U12225 ( .ip(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[1]), .op(n10833)
         );
  inv_1 U12226 ( .ip(n10843), .op(n10852) );
  nor2_1 U12227 ( .ip1(n10831), .ip2(n10852), .op(n10832) );
  nor2_1 U12228 ( .ip1(n10833), .ip2(n10832), .op(n10834) );
  mux2_1 U12229 ( .ip1(i_ssi_rx_push_data[1]), .ip2(n10834), .s(n10122), .op(
        n4437) );
  mux2_1 U12230 ( .ip1(i_ssi_U_dff_rx_mem[65]), .ip2(i_ssi_rx_push_data[1]), 
        .s(n10721), .op(n4358) );
  mux2_1 U12231 ( .ip1(i_ssi_U_dff_rx_mem[33]), .ip2(i_ssi_rx_push_data[1]), 
        .s(n5610), .op(n4360) );
  mux2_1 U12232 ( .ip1(i_ssi_U_dff_rx_mem[1]), .ip2(i_ssi_rx_push_data[1]), 
        .s(n10777), .op(n4362) );
  mux2_1 U12233 ( .ip1(i_ssi_rx_push_data[1]), .ip2(i_ssi_U_dff_rx_mem[113]), 
        .s(n11455), .op(n4355) );
  mux2_1 U12234 ( .ip1(i_ssi_rx_push_data[1]), .ip2(i_ssi_U_dff_rx_mem[81]), 
        .s(n11454), .op(n4357) );
  mux2_1 U12235 ( .ip1(i_ssi_rx_push_data[1]), .ip2(i_ssi_U_dff_rx_mem[17]), 
        .s(n11452), .op(n4361) );
  mux2_1 U12236 ( .ip1(i_ssi_rx_push_data[1]), .ip2(i_ssi_U_dff_rx_mem[49]), 
        .s(n11453), .op(n4359) );
  mux2_1 U12237 ( .ip1(i_ssi_U_dff_rx_mem[97]), .ip2(i_ssi_rx_push_data[1]), 
        .s(n5611), .op(n4356) );
  mux2_1 U12238 ( .ip1(i_apb_pwdata_int[2]), .ip2(i_ssi_rxftlr[2]), .s(n10835), 
        .op(n4635) );
  mux2_1 U12239 ( .ip1(i_apb_pwdata_int[2]), .ip2(i_ssi_mwcr[2]), .s(n10836), 
        .op(n4628) );
  inv_1 U12240 ( .ip(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[2]), .op(n10838)
         );
  nor2_1 U12241 ( .ip1(n5351), .ip2(n10852), .op(n10837) );
  nor2_1 U12242 ( .ip1(n10838), .ip2(n10837), .op(n10839) );
  mux2_1 U12243 ( .ip1(i_ssi_rx_push_data[2]), .ip2(n10839), .s(n10122), .op(
        n4436) );
  mux2_1 U12244 ( .ip1(i_ssi_U_dff_rx_mem[2]), .ip2(i_ssi_rx_push_data[2]), 
        .s(n10777), .op(n4354) );
  mux2_1 U12245 ( .ip1(i_ssi_U_dff_rx_mem[34]), .ip2(i_ssi_rx_push_data[2]), 
        .s(n5610), .op(n4352) );
  mux2_1 U12246 ( .ip1(i_ssi_U_dff_rx_mem[66]), .ip2(i_ssi_rx_push_data[2]), 
        .s(n10721), .op(n4350) );
  mux2_1 U12247 ( .ip1(i_ssi_rx_push_data[2]), .ip2(i_ssi_U_dff_rx_mem[50]), 
        .s(n11453), .op(n4351) );
  mux2_1 U12248 ( .ip1(i_ssi_rx_push_data[2]), .ip2(i_ssi_U_dff_rx_mem[114]), 
        .s(n11455), .op(n4347) );
  mux2_1 U12249 ( .ip1(i_ssi_U_dff_rx_mem[98]), .ip2(i_ssi_rx_push_data[2]), 
        .s(n5611), .op(n4348) );
  mux2_1 U12250 ( .ip1(i_ssi_rx_push_data[2]), .ip2(i_ssi_U_dff_rx_mem[18]), 
        .s(n11452), .op(n4353) );
  mux2_1 U12251 ( .ip1(i_ssi_rx_push_data[2]), .ip2(i_ssi_U_dff_rx_mem[82]), 
        .s(n11454), .op(n4349) );
  inv_1 U12252 ( .ip(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[3]), .op(n10841)
         );
  nor2_1 U12253 ( .ip1(n10852), .ip2(n10866), .op(n10840) );
  nor2_1 U12254 ( .ip1(n10841), .ip2(n10840), .op(n10842) );
  mux2_1 U12255 ( .ip1(i_ssi_rx_push_data[3]), .ip2(n10842), .s(n10122), .op(
        n4435) );
  mux2_1 U12256 ( .ip1(i_ssi_U_dff_rx_mem[35]), .ip2(i_ssi_rx_push_data[3]), 
        .s(n5610), .op(n4344) );
  mux2_1 U12257 ( .ip1(i_ssi_U_dff_rx_mem[67]), .ip2(i_ssi_rx_push_data[3]), 
        .s(n10721), .op(n4342) );
  mux2_1 U12258 ( .ip1(i_ssi_U_dff_rx_mem[99]), .ip2(i_ssi_rx_push_data[3]), 
        .s(n5611), .op(n4340) );
  mux2_1 U12259 ( .ip1(i_ssi_rx_push_data[3]), .ip2(i_ssi_U_dff_rx_mem[51]), 
        .s(n11453), .op(n4343) );
  mux2_1 U12260 ( .ip1(i_ssi_U_dff_rx_mem[3]), .ip2(i_ssi_rx_push_data[3]), 
        .s(n10777), .op(n4346) );
  mux2_1 U12261 ( .ip1(i_ssi_rx_push_data[3]), .ip2(i_ssi_U_dff_rx_mem[19]), 
        .s(n11452), .op(n4345) );
  mux2_1 U12262 ( .ip1(i_ssi_rx_push_data[3]), .ip2(i_ssi_U_dff_rx_mem[83]), 
        .s(n11454), .op(n4341) );
  mux2_1 U12263 ( .ip1(i_ssi_rx_push_data[3]), .ip2(i_ssi_U_dff_rx_mem[115]), 
        .s(n11455), .op(n4339) );
  inv_1 U12264 ( .ip(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[4]), .op(n10844)
         );
  nor2_1 U12265 ( .ip1(n10844), .ip2(n10843), .op(n10845) );
  mux2_1 U12266 ( .ip1(i_ssi_rx_push_data[4]), .ip2(n10845), .s(n10122), .op(
        n4434) );
  mux2_1 U12267 ( .ip1(i_ssi_rx_push_data[4]), .ip2(i_ssi_U_dff_rx_mem[52]), 
        .s(n11453), .op(n4335) );
  mux2_1 U12268 ( .ip1(i_ssi_U_dff_rx_mem[36]), .ip2(i_ssi_rx_push_data[4]), 
        .s(n5610), .op(n4336) );
  mux2_1 U12269 ( .ip1(i_ssi_rx_push_data[4]), .ip2(i_ssi_U_dff_rx_mem[20]), 
        .s(n11452), .op(n4337) );
  mux2_1 U12270 ( .ip1(i_ssi_U_dff_rx_mem[68]), .ip2(i_ssi_rx_push_data[4]), 
        .s(n10721), .op(n4334) );
  mux2_1 U12271 ( .ip1(i_ssi_U_dff_rx_mem[100]), .ip2(i_ssi_rx_push_data[4]), 
        .s(n5611), .op(n4332) );
  mux2_1 U12272 ( .ip1(i_ssi_U_dff_rx_mem[4]), .ip2(i_ssi_rx_push_data[4]), 
        .s(n10777), .op(n4338) );
  mux2_1 U12273 ( .ip1(i_ssi_rx_push_data[4]), .ip2(i_ssi_U_dff_rx_mem[116]), 
        .s(n11455), .op(n4331) );
  mux2_1 U12274 ( .ip1(i_ssi_rx_push_data[4]), .ip2(i_ssi_U_dff_rx_mem[84]), 
        .s(n11454), .op(n4333) );
  mux2_1 U12275 ( .ip1(i_ssi_imr[4]), .ip2(i_apb_pwdata_int[4]), .s(n10846), 
        .op(n4639) );
  nor2_1 U12276 ( .ip1(n10848), .ip2(n10847), .op(n10850) );
  nor2_1 U12277 ( .ip1(i_ssi_U_fifo_switch_almost_full), .ip2(n10850), .op(
        n10849) );
  not_ab_or_c_or_d U12278 ( .ip1(n10851), .ip2(n10850), .ip3(n5291), .ip4(
        n10849), .op(i_ssi_U_intctl_N33) );
  nand2_1 U12279 ( .ip1(i_ssi_imr[4]), .ip2(i_ssi_risr[4]), .op(
        i_ssi_ssi_rxf_intr_n) );
  nand3_1 U12280 ( .ip1(n10122), .ip2(n5343), .ip3(n10852), .op(n10853) );
  nand2_1 U12281 ( .ip1(n10853), .ip2(n10858), .op(n10854) );
  nand2_1 U12282 ( .ip1(n10854), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[5]), .op(n10856) );
  nand2_1 U12283 ( .ip1(n10868), .ip2(i_ssi_rx_push_data[5]), .op(n10855) );
  nand2_1 U12284 ( .ip1(n10856), .ip2(n10855), .op(n4433) );
  mux2_1 U12285 ( .ip1(i_ssi_rx_push_data[5]), .ip2(i_ssi_U_dff_rx_mem[21]), 
        .s(n11452), .op(n4329) );
  mux2_1 U12286 ( .ip1(i_ssi_U_dff_rx_mem[37]), .ip2(i_ssi_rx_push_data[5]), 
        .s(n5610), .op(n4328) );
  mux2_1 U12287 ( .ip1(i_ssi_U_dff_rx_mem[69]), .ip2(i_ssi_rx_push_data[5]), 
        .s(n10721), .op(n4326) );
  mux2_1 U12288 ( .ip1(i_ssi_rx_push_data[5]), .ip2(i_ssi_U_dff_rx_mem[53]), 
        .s(n11453), .op(n4327) );
  mux2_1 U12289 ( .ip1(i_ssi_rx_push_data[5]), .ip2(i_ssi_U_dff_rx_mem[85]), 
        .s(n11454), .op(n4325) );
  mux2_1 U12290 ( .ip1(i_ssi_U_dff_rx_mem[101]), .ip2(i_ssi_rx_push_data[5]), 
        .s(n5611), .op(n4324) );
  mux2_1 U12291 ( .ip1(i_ssi_rx_push_data[5]), .ip2(i_ssi_U_dff_rx_mem[117]), 
        .s(n11455), .op(n4323) );
  mux2_1 U12292 ( .ip1(i_ssi_U_dff_rx_mem[5]), .ip2(i_ssi_rx_push_data[5]), 
        .s(n10777), .op(n4330) );
  inv_1 U12293 ( .ip(i_ssi_rx_push_data[7]), .op(n10857) );
  nor2_1 U12294 ( .ip1(n10857), .ip2(n10122), .op(n10862) );
  inv_1 U12295 ( .ip(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[7]), .op(n10859)
         );
  not_ab_or_c_or_d U12296 ( .ip1(n10860), .ip2(n11471), .ip3(n10859), .ip4(
        n10858), .op(n10861) );
  or2_1 U12297 ( .ip1(n10862), .ip2(n10861), .op(n4431) );
  mux2_1 U12298 ( .ip1(i_ssi_rx_push_data[7]), .ip2(i_ssi_U_dff_rx_mem[87]), 
        .s(n11454), .op(n4309) );
  mux2_1 U12299 ( .ip1(i_ssi_U_dff_rx_mem[39]), .ip2(i_ssi_rx_push_data[7]), 
        .s(n5610), .op(n4312) );
  mux2_1 U12300 ( .ip1(i_ssi_rx_push_data[7]), .ip2(i_ssi_U_dff_rx_mem[23]), 
        .s(n11452), .op(n4313) );
  mux2_1 U12301 ( .ip1(i_ssi_U_dff_rx_mem[7]), .ip2(i_ssi_rx_push_data[7]), 
        .s(n10777), .op(n4314) );
  mux2_1 U12302 ( .ip1(i_ssi_rx_push_data[7]), .ip2(i_ssi_U_dff_rx_mem[55]), 
        .s(n11453), .op(n4311) );
  mux2_1 U12303 ( .ip1(i_ssi_U_dff_rx_mem[71]), .ip2(i_ssi_rx_push_data[7]), 
        .s(n10721), .op(n4310) );
  mux2_1 U12304 ( .ip1(i_ssi_rx_push_data[7]), .ip2(i_ssi_U_dff_rx_mem[119]), 
        .s(n11455), .op(n4307) );
  mux2_1 U12305 ( .ip1(i_ssi_U_dff_rx_mem[103]), .ip2(i_ssi_rx_push_data[7]), 
        .s(n5611), .op(n4308) );
  mux2_1 U12306 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[14]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[13]), .s(n10865), .op(n4373)
         );
  nand3_1 U12307 ( .ip1(n10867), .ip2(n5351), .ip3(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[14]), .op(n10864) );
  nand2_1 U12308 ( .ip1(n10868), .ip2(i_ssi_rx_push_data[14]), .op(n10863) );
  nand2_1 U12309 ( .ip1(n10864), .ip2(n10863), .op(n4424) );
  mux2_1 U12310 ( .ip1(i_ssi_rx_push_data[14]), .ip2(i_ssi_U_dff_rx_mem[62]), 
        .s(n11453), .op(n4255) );
  mux2_1 U12311 ( .ip1(i_ssi_U_dff_rx_mem[46]), .ip2(i_ssi_rx_push_data[14]), 
        .s(n5610), .op(n4256) );
  mux2_1 U12312 ( .ip1(i_ssi_rx_push_data[14]), .ip2(i_ssi_U_dff_rx_mem[94]), 
        .s(n11454), .op(n4253) );
  mux2_1 U12313 ( .ip1(i_ssi_rx_push_data[14]), .ip2(i_ssi_U_dff_rx_mem[30]), 
        .s(n11452), .op(n4257) );
  mux2_1 U12314 ( .ip1(i_ssi_U_dff_rx_mem[110]), .ip2(i_ssi_rx_push_data[14]), 
        .s(n5611), .op(n4252) );
  mux2_1 U12315 ( .ip1(i_ssi_U_dff_rx_mem[14]), .ip2(i_ssi_rx_push_data[14]), 
        .s(n10777), .op(n4258) );
  mux2_1 U12316 ( .ip1(i_ssi_U_dff_rx_mem[78]), .ip2(i_ssi_rx_push_data[14]), 
        .s(n10721), .op(n4254) );
  mux2_1 U12317 ( .ip1(i_ssi_rx_push_data[14]), .ip2(i_ssi_U_dff_rx_mem[126]), 
        .s(n11455), .op(n4251) );
  mux2_1 U12318 ( .ip1(i_ssi_U_shift_U_rx_shifter_rx_shift_reg[15]), .ip2(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[14]), .s(n10865), .op(n4372)
         );
  nand3_1 U12319 ( .ip1(n10867), .ip2(n10866), .ip3(
        i_ssi_U_shift_U_rx_shifter_rx_shift_reg[15]), .op(n10870) );
  nand2_1 U12320 ( .ip1(n10868), .ip2(i_ssi_rx_push_data[15]), .op(n10869) );
  nand2_1 U12321 ( .ip1(n10870), .ip2(n10869), .op(n4423) );
  mux2_1 U12322 ( .ip1(i_ssi_rx_push_data[15]), .ip2(i_ssi_U_dff_rx_mem[31]), 
        .s(n11452), .op(n4249) );
  mux2_1 U12323 ( .ip1(i_ssi_U_dff_rx_mem[47]), .ip2(i_ssi_rx_push_data[15]), 
        .s(n5610), .op(n4248) );
  mux2_1 U12324 ( .ip1(i_ssi_rx_push_data[15]), .ip2(i_ssi_U_dff_rx_mem[95]), 
        .s(n11454), .op(n4245) );
  mux2_1 U12325 ( .ip1(i_ssi_rx_push_data[15]), .ip2(i_ssi_U_dff_rx_mem[127]), 
        .s(n11455), .op(n4243) );
  mux2_1 U12326 ( .ip1(i_ssi_U_dff_rx_mem[111]), .ip2(i_ssi_rx_push_data[15]), 
        .s(n5611), .op(n4244) );
  mux2_1 U12327 ( .ip1(i_ssi_rx_push_data[15]), .ip2(i_ssi_U_dff_rx_mem[63]), 
        .s(n11453), .op(n4247) );
  mux2_1 U12328 ( .ip1(i_ssi_U_dff_rx_mem[15]), .ip2(i_ssi_rx_push_data[15]), 
        .s(n10777), .op(n4250) );
  mux2_1 U12329 ( .ip1(i_ssi_U_dff_rx_mem[79]), .ip2(i_ssi_rx_push_data[15]), 
        .s(n10721), .op(n4246) );
  inv_1 U12330 ( .ip(n11296), .op(n10872) );
  nand2_1 U12331 ( .ip1(n10872), .ip2(n10871), .op(n10874) );
  nand2_1 U12332 ( .ip1(n11126), .ip2(i_i2c_mst_rxbyte_rdy), .op(n10873) );
  nand2_1 U12333 ( .ip1(n10874), .ip2(n10873), .op(
        i_i2c_U_DW_apb_i2c_rx_shift_N30) );
  nor2_1 U12334 ( .ip1(n10876), .ip2(n10875), .op(n10877) );
  mux2_1 U12335 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[0]), .ip2(
        n11833), .s(n10877), .op(n4929) );
  nor2_1 U12336 ( .ip1(n10881), .ip2(n10878), .op(n10885) );
  nand2_1 U12337 ( .ip1(n10885), .ip2(i_i2c_mst_rx_bit_count[2]), .op(n10879)
         );
  mux2_1 U12338 ( .ip1(n11833), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[1]), .s(n10879), .op(
        n4928) );
  nand2_1 U12339 ( .ip1(n10888), .ip2(i_i2c_mst_rx_bit_count[2]), .op(n10880)
         );
  mux2_1 U12340 ( .ip1(n11833), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[2]), .s(n10880), .op(
        n4927) );
  nand3_1 U12341 ( .ip1(n10882), .ip2(i_i2c_mst_rx_bit_count[2]), .ip3(n10881), 
        .op(n10883) );
  mux2_1 U12342 ( .ip1(n11833), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[3]), .s(n10883), .op(
        n4926) );
  mux2_1 U12343 ( .ip1(n11833), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[4]), .s(n10884), .op(
        n4925) );
  nand2_1 U12344 ( .ip1(n10885), .ip2(n10887), .op(n10886) );
  mux2_1 U12345 ( .ip1(n11833), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[5]), .s(n10886), .op(
        n4924) );
  nand2_1 U12346 ( .ip1(n10888), .ip2(n10887), .op(n10889) );
  mux2_1 U12347 ( .ip1(n11833), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[6]), .s(n10889), .op(
        n4923) );
  nand2_1 U12348 ( .ip1(n10890), .ip2(n11038), .op(n10891) );
  mux2_1 U12349 ( .ip1(n11833), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[7]), .s(n10891), .op(
        n4922) );
  inv_1 U12350 ( .ip(n10919), .op(n11066) );
  nor2_1 U12351 ( .ip1(n11066), .ip2(n10947), .op(n10950) );
  nand2_1 U12352 ( .ip1(n10938), .ip2(i_i2c_ic_tar[7]), .op(n10894) );
  nand2_1 U12353 ( .ip1(n10941), .ip2(i_i2c_tx_fifo_data_buf[7]), .op(n10893)
         );
  nand2_1 U12354 ( .ip1(n10942), .ip2(i_i2c_ic_tar[6]), .op(n10892) );
  nand3_1 U12355 ( .ip1(n10894), .ip2(n10893), .ip3(n10892), .op(n10895) );
  mux2_1 U12356 ( .ip1(n10895), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[7]), .s(n10947), .op(n10896)
         );
  or2_1 U12357 ( .ip1(n10950), .ip2(n10896), .op(n5033) );
  inv_1 U12358 ( .ip(i_i2c_ic_tar[5]), .op(n10934) );
  nor2_1 U12359 ( .ip1(n10934), .ip2(n10917), .op(n10899) );
  nor2_1 U12360 ( .ip1(n10897), .ip2(n11068), .op(n10898) );
  not_ab_or_c_or_d U12361 ( .ip1(n10942), .ip2(i_i2c_ic_tar[4]), .ip3(n10899), 
        .ip4(n10898), .op(n10900) );
  nor2_1 U12362 ( .ip1(n10900), .ip2(n10947), .op(n10901) );
  ab_or_c_or_d U12363 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[5]), 
        .ip2(n10947), .ip3(n10901), .ip4(n10950), .op(n5035) );
  nand2_1 U12364 ( .ip1(n10938), .ip2(i_i2c_ic_tar[3]), .op(n10906) );
  nand2_1 U12365 ( .ip1(n10942), .ip2(i_i2c_ic_tar[2]), .op(n10904) );
  nand2_1 U12366 ( .ip1(n10902), .ip2(i_i2c_tx_fifo_data_buf[3]), .op(n10903)
         );
  nand4_1 U12367 ( .ip1(n10906), .ip2(n10905), .ip3(n10904), .ip4(n10903), 
        .op(n10907) );
  mux2_1 U12368 ( .ip1(n10907), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[3]), .s(n10947), .op(n5037)
         );
  inv_1 U12369 ( .ip(i_i2c_ic_tar[1]), .op(n10908) );
  nor2_1 U12370 ( .ip1(n10908), .ip2(n10917), .op(n10913) );
  nand2_1 U12371 ( .ip1(n10941), .ip2(i_i2c_tx_fifo_data_buf[1]), .op(n10911)
         );
  nand2_1 U12372 ( .ip1(n10919), .ip2(i_i2c_ic_tar[8]), .op(n10910) );
  nand2_1 U12373 ( .ip1(n10926), .ip2(i_i2c_ic_hs_maddr[1]), .op(n10909) );
  nand3_1 U12374 ( .ip1(n10911), .ip2(n10910), .ip3(n10909), .op(n10912) );
  not_ab_or_c_or_d U12375 ( .ip1(n10942), .ip2(i_i2c_ic_tar[0]), .ip3(n10913), 
        .ip4(n10912), .op(n10915) );
  mux2_1 U12376 ( .ip1(n10915), .ip2(n10914), .s(n10947), .op(n10916) );
  inv_1 U12377 ( .ip(n10916), .op(n5039) );
  inv_1 U12378 ( .ip(i_i2c_ic_tar[2]), .op(n10918) );
  nor2_1 U12379 ( .ip1(n10918), .ip2(n10917), .op(n10924) );
  nand2_1 U12380 ( .ip1(n10941), .ip2(i_i2c_tx_fifo_data_buf[2]), .op(n10922)
         );
  nand2_1 U12381 ( .ip1(n10919), .ip2(i_i2c_ic_tar[9]), .op(n10921) );
  nand2_1 U12382 ( .ip1(n10926), .ip2(i_i2c_ic_hs_maddr[2]), .op(n10920) );
  nand3_1 U12383 ( .ip1(n10922), .ip2(n10921), .ip3(n10920), .op(n10923) );
  ab_or_c_or_d U12384 ( .ip1(i_i2c_ic_tar[1]), .ip2(n10942), .ip3(n10924), 
        .ip4(n10923), .op(n10925) );
  mux2_1 U12385 ( .ip1(n10925), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[2]), .s(n10947), .op(n5038)
         );
  nand2_1 U12386 ( .ip1(n10941), .ip2(i_i2c_tx_fifo_data_buf[0]), .op(n10928)
         );
  nand2_1 U12387 ( .ip1(n10926), .ip2(i_i2c_ic_hs_maddr[0]), .op(n10927) );
  nand2_1 U12388 ( .ip1(n10928), .ip2(n10927), .op(n10929) );
  not_ab_or_c_or_d U12389 ( .ip1(i_i2c_ic_tar[0]), .ip2(n10938), .ip3(n10930), 
        .ip4(n10929), .op(n10931) );
  nand2_1 U12390 ( .ip1(n10932), .ip2(n10931), .op(n10933) );
  mux2_1 U12391 ( .ip1(n10933), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[0]), .s(n10947), .op(n5040)
         );
  nor2_1 U12392 ( .ip1(n10934), .ip2(n11071), .op(n10937) );
  inv_1 U12393 ( .ip(i_i2c_tx_fifo_data_buf[6]), .op(n10935) );
  nor2_1 U12394 ( .ip1(n10935), .ip2(n11068), .op(n10936) );
  not_ab_or_c_or_d U12395 ( .ip1(i_i2c_ic_tar[6]), .ip2(n10938), .ip3(n10937), 
        .ip4(n10936), .op(n10939) );
  nor2_1 U12396 ( .ip1(n10939), .ip2(n10947), .op(n10940) );
  ab_or_c_or_d U12397 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[6]), 
        .ip2(n10947), .ip3(n10940), .ip4(n10950), .op(n5034) );
  nand2_1 U12398 ( .ip1(n10941), .ip2(i_i2c_tx_fifo_data_buf[4]), .op(n10946)
         );
  nand2_1 U12399 ( .ip1(n10942), .ip2(i_i2c_ic_tar[3]), .op(n10945) );
  nand2_1 U12400 ( .ip1(n10943), .ip2(i_i2c_ic_tar[4]), .op(n10944) );
  nand3_1 U12401 ( .ip1(n10946), .ip2(n10945), .ip3(n10944), .op(n10948) );
  mux2_1 U12402 ( .ip1(n10948), .ip2(
        i_i2c_U_DW_apb_i2c_tx_shift_tx_shift_buf[4]), .s(n10947), .op(n10949)
         );
  or2_1 U12403 ( .ip1(n10950), .ip2(n10949), .op(n5036) );
  and2_1 U12404 ( .ip1(n5291), .ip2(i_ssi_fsm_sleep), .op(i_ssi_U_regfile_N451) );
  nor2_1 U12405 ( .ip1(n10978), .ip2(n10951), .op(n10955) );
  inv_1 U12406 ( .ip(n5247), .op(n10954) );
  inv_1 U12407 ( .ip(i_ssi_ser_0_), .op(n10953) );
  not_ab_or_c_or_d U12408 ( .ip1(n10955), .ip2(n10954), .ip3(n10953), .ip4(
        n10952), .op(n11838) );
  mux2_1 U12409 ( .ip1(i_apb_pwdata_int[7]), .ip2(
        i_ssi_U_regfile_ctrlr0_ir_int_7), .s(n11097), .op(n4587) );
  inv_1 U12410 ( .ip(i_apb_pwdata_int[5]), .op(n10961) );
  nand2_1 U12411 ( .ip1(n10962), .ip2(n10961), .op(n10956) );
  nand2_1 U12412 ( .ip1(n10956), .ip2(i_ssi_U_regfile_ctrlr0_ir_int[5]), .op(
        n10958) );
  nand3_1 U12413 ( .ip1(n10962), .ip2(i_apb_pwdata_int[5]), .ip3(n10959), .op(
        n10957) );
  nand2_1 U12414 ( .ip1(n10958), .ip2(n10957), .op(n4586) );
  nand2_1 U12415 ( .ip1(n10962), .ip2(n10959), .op(n10960) );
  nand2_1 U12416 ( .ip1(n10960), .ip2(i_ssi_U_regfile_ctrlr0_ir_int[4]), .op(
        n10964) );
  nand3_1 U12417 ( .ip1(n10962), .ip2(i_apb_pwdata_int[4]), .ip3(n10961), .op(
        n10963) );
  nand2_1 U12418 ( .ip1(n10964), .ip2(n10963), .op(n4585) );
  nor2_1 U12419 ( .ip1(i_ssi_U_regfile_ctrlr0_ir_int[5]), .ip2(
        i_ssi_U_regfile_ctrlr0_ir_int[4]), .op(n10965) );
  nand2_1 U12420 ( .ip1(n10965), .ip2(i_ssi_U_regfile_ctrlr0_ir_int_7), .op(
        n5235) );
  inv_1 U12421 ( .ip(i_ssi_sclk_active), .op(n10986) );
  nand2_1 U12422 ( .ip1(n10966), .ip2(n5247), .op(n10975) );
  nor4_1 U12423 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[2]), .ip2(
        i_ssi_U_sclkgen_ssi_cnt[1]), .ip3(i_ssi_U_sclkgen_ssi_cnt[5]), .ip4(
        i_ssi_U_sclkgen_ssi_cnt[8]), .op(n10969) );
  nor4_2 U12424 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[9]), .ip2(
        i_ssi_U_sclkgen_ssi_cnt[6]), .ip3(i_ssi_U_sclkgen_ssi_cnt[15]), .ip4(
        i_ssi_U_sclkgen_ssi_cnt[3]), .op(n10968) );
  nor4_1 U12425 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[11]), .ip2(
        i_ssi_U_sclkgen_ssi_cnt[13]), .ip3(i_ssi_U_sclkgen_ssi_cnt[4]), .ip4(
        i_ssi_U_sclkgen_ssi_cnt[0]), .op(n10967) );
  and4_1 U12426 ( .ip1(n10970), .ip2(n10969), .ip3(n10968), .ip4(n10967), .op(
        n10971) );
  not_ab_or_c_or_d U12427 ( .ip1(n10973), .ip2(n10972), .ip3(n10971), .ip4(
        n5291), .op(n10974) );
  nand2_1 U12428 ( .ip1(n10975), .ip2(n10974), .op(n10991) );
  nor2_1 U12429 ( .ip1(n10987), .ip2(n10981), .op(n10976) );
  nor2_1 U12430 ( .ip1(n10991), .ip2(n10976), .op(n10984) );
  nand2_1 U12431 ( .ip1(n10978), .ip2(n5492), .op(n10979) );
  nand2_1 U12432 ( .ip1(n10982), .ip2(n10990), .op(n10983) );
  nand2_1 U12433 ( .ip1(n10984), .ip2(n10983), .op(n10985) );
  nand2_1 U12434 ( .ip1(n10986), .ip2(n10985), .op(n11016) );
  nand2_1 U12435 ( .ip1(n10988), .ip2(n10987), .op(n10989) );
  nand2_1 U12436 ( .ip1(n10990), .ip2(n10989), .op(n11014) );
  inv_1 U12437 ( .ip(n10991), .op(n11013) );
  xor2_1 U12438 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[7]), .ip2(i_ssi_baudr[8]), .op(
        n10995) );
  xor2_1 U12439 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[4]), .ip2(i_ssi_baudr[5]), .op(
        n10994) );
  xor2_1 U12440 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[10]), .ip2(i_ssi_baudr[11]), 
        .op(n10993) );
  xor2_1 U12441 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[12]), .ip2(i_ssi_baudr[13]), 
        .op(n10992) );
  xor2_1 U12442 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[2]), .ip2(i_ssi_baudr[3]), .op(
        n10999) );
  xor2_1 U12443 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[13]), .ip2(i_ssi_baudr[14]), 
        .op(n10998) );
  xor2_1 U12444 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[11]), .ip2(i_ssi_baudr[12]), 
        .op(n10997) );
  xor2_1 U12445 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[5]), .ip2(i_ssi_baudr[6]), .op(
        n11003) );
  xor2_1 U12446 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[6]), .ip2(i_ssi_baudr[7]), .op(
        n11002) );
  xor2_1 U12447 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[3]), .ip2(i_ssi_baudr[4]), .op(
        n11001) );
  xor2_1 U12448 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[14]), .ip2(i_ssi_baudr[15]), 
        .op(n11000) );
  xor2_1 U12449 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[1]), .ip2(i_ssi_baudr[2]), .op(
        n11006) );
  xor2_1 U12450 ( .ip1(i_ssi_U_sclkgen_ssi_cnt[8]), .ip2(i_ssi_baudr[9]), .op(
        n11005) );
  nor3_1 U12451 ( .ip1(n11006), .ip2(n11005), .ip3(n11004), .op(n11007) );
  nand4_1 U12452 ( .ip1(n11010), .ip2(n11009), .ip3(n11008), .ip4(n11007), 
        .op(n11011) );
  mux2_1 U12453 ( .ip1(i_ssi_sclk_active), .ip2(i_ssi_sclk_out), .s(n11011), 
        .op(n11012) );
  nand3_1 U12454 ( .ip1(n11014), .ip2(n11013), .ip3(n11012), .op(n11015) );
  nand2_1 U12455 ( .ip1(n11016), .ip2(n11015), .op(n4242) );
  nor3_1 U12456 ( .ip1(n11018), .ip2(n11017), .ip3(n11052), .op(
        i_i2c_U_DW_apb_i2c_toggle_N33) );
  nand3_1 U12457 ( .ip1(n11019), .ip2(i_i2c_slv_debug_cstate[0]), .ip3(
        i_i2c_slv_debug_cstate[2]), .op(n11020) );
  nand3_1 U12458 ( .ip1(n11068), .ip2(n11021), .ip3(n11020), .op(
        i_i2c_U_DW_apb_i2c_toggle_N31) );
  inv_1 U12459 ( .ip(n11022), .op(n11024) );
  nand3_1 U12460 ( .ip1(n11024), .ip2(n11244), .ip3(n11023), .op(
        i_i2c_U_DW_apb_i2c_toggle_N32) );
  inv_1 U12461 ( .ip(i_i2c_ic_tx_tl[1]), .op(n11140) );
  nand2_1 U12462 ( .ip1(n11029), .ip2(n11140), .op(n11025) );
  nand2_1 U12463 ( .ip1(n11025), .ip2(i_i2c_ic_tx_tl[2]), .op(n11028) );
  nor3_1 U12464 ( .ip1(i_i2c_ic_tx_tl[2]), .ip2(n11026), .ip3(n11025), .op(
        n11027) );
  not_ab_or_c_or_d U12465 ( .ip1(n11866), .ip2(n11028), .ip3(n11027), .ip4(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N37), .op(n11034) );
  nor2_1 U12466 ( .ip1(n11029), .ip2(n11140), .op(n11030) );
  not_ab_or_c_or_d U12467 ( .ip1(i_i2c_ic_tx_tl[2]), .ip2(n11031), .ip3(n11030), .ip4(i_i2c_ic_tx_tl[0]), .op(n11032) );
  nand2_1 U12468 ( .ip1(n11032), .ip2(n11867), .op(n11033) );
  nand2_1 U12469 ( .ip1(n11034), .ip2(n11033), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N34) );
  nor2_1 U12470 ( .ip1(n11055), .ip2(n11035), .op(n11036) );
  xor2_1 U12471 ( .ip1(i_i2c_tx_abrt_source[5]), .ip2(n11036), .op(n4933) );
  or2_1 U12472 ( .ip1(i_i2c_split_start_en), .ip2(i_i2c_re_start_en), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_N207) );
  nand2_1 U12473 ( .ip1(n11038), .ip2(n11037), .op(n11039) );
  and2_1 U12474 ( .ip1(n11039), .ip2(i_i2c_rx_current_src_en), .op(n11043) );
  nor4_1 U12475 ( .ip1(i_i2c_mst_rx_bit_count[3]), .ip2(n11041), .ip3(n11040), 
        .ip4(n11045), .op(n11042) );
  nor2_1 U12476 ( .ip1(n11043), .ip2(n11042), .op(n11044) );
  nor2_1 U12477 ( .ip1(n11044), .ip2(n11052), .op(n5063) );
  nor4_1 U12478 ( .ip1(i_i2c_U_DW_apb_i2c_tx_shift_tx_bit_count[3]), .ip2(
        n11046), .ip3(n11045), .ip4(n11048), .op(n11051) );
  nand2_1 U12479 ( .ip1(n11048), .ip2(n11047), .op(n11049) );
  and2_1 U12480 ( .ip1(n11049), .ip2(i_i2c_tx_current_src_en), .op(n11050) );
  nor2_1 U12481 ( .ip1(n11051), .ip2(n11050), .op(n11053) );
  nor2_1 U12482 ( .ip1(n11053), .ip2(n11052), .op(n5062) );
  or2_1 U12483 ( .ip1(i_i2c_rx_current_src_en), .ip2(i_i2c_tx_current_src_en), 
        .op(i_i2c_U_DW_apb_i2c_toggle_N29) );
  xor2_1 U12484 ( .ip1(i_i2c_tx_abrt_source[16]), .ip2(n11054), .op(n5198) );
  nand2_1 U12485 ( .ip1(n11056), .ip2(n11055), .op(n11058) );
  nand2_1 U12486 ( .ip1(n11058), .ip2(n11057), .op(n11059) );
  nand2_1 U12487 ( .ip1(n11059), .ip2(n11096), .op(n11060) );
  xnor2_1 U12488 ( .ip1(i_i2c_tx_abrt_source[14]), .ip2(n11060), .op(n5213) );
  xor2_1 U12489 ( .ip1(i_i2c_tx_abrt_source[10]), .ip2(n11061), .op(n5202) );
  nor2_1 U12490 ( .ip1(n11062), .ip2(n11070), .op(n11063) );
  xor2_1 U12491 ( .ip1(i_i2c_tx_abrt_source[4]), .ip2(n11063), .op(n5179) );
  nor2_1 U12492 ( .ip1(n11064), .ip2(n11070), .op(n11065) );
  xor2_1 U12493 ( .ip1(i_i2c_tx_abrt_source[2]), .ip2(n11065), .op(n5181) );
  nor2_1 U12494 ( .ip1(n11066), .ip2(n11070), .op(n11067) );
  xor2_1 U12495 ( .ip1(i_i2c_tx_abrt_source[1]), .ip2(n11067), .op(n5185) );
  nor2_1 U12496 ( .ip1(n11068), .ip2(n11070), .op(n11069) );
  xor2_1 U12497 ( .ip1(i_i2c_tx_abrt_source[3]), .ip2(n11069), .op(n5186) );
  nor2_1 U12498 ( .ip1(n11071), .ip2(n11070), .op(n11072) );
  xor2_1 U12499 ( .ip1(i_i2c_tx_abrt_source[0]), .ip2(n11072), .op(n5187) );
  nor2_1 U12500 ( .ip1(n11074), .ip2(n11073), .op(n11075) );
  xor2_1 U12501 ( .ip1(i_i2c_tx_abrt_source[7]), .ip2(n11075), .op(n5180) );
  xor2_1 U12502 ( .ip1(i_i2c_tx_abrt_source[6]), .ip2(n11076), .op(n5182) );
  nor3_1 U12503 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_10bit_slv_sync_inv), .ip2(
        n11078), .ip3(n11077), .op(n11081) );
  nor2_1 U12504 ( .ip1(n11288), .ip2(
        i_i2c_U_DW_apb_i2c_sync_ic_10bit_slv_sync_inv), .op(n11079) );
  inv_1 U12505 ( .ip(i_i2c_rx_addr_match), .op(n11232) );
  not_ab_or_c_or_d U12506 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_10bit_slv_sync_inv), .ip2(n11299), .ip3(n11079), .ip4(n11232), .op(n11080) );
  nor3_1 U12507 ( .ip1(i_i2c_slv_addressed), .ip2(n11081), .ip3(n11080), .op(
        n11082) );
  nor2_1 U12508 ( .ip1(n11083), .ip2(n11082), .op(n5078) );
  inv_1 U12509 ( .ip(i_i2c_slv_addressed), .op(n11084) );
  nand3_1 U12510 ( .ip1(n11084), .ip2(
        i_i2c_U_DW_apb_i2c_sync_ic_master_sync_inv), .ip3(
        i_i2c_p_det_ifaddr_sync), .op(n11085) );
  and2_1 U12511 ( .ip1(n11864), .ip2(n11085), .op(
        i_i2c_U_DW_apb_i2c_rx_filter_N241) );
  xor2_1 U12512 ( .ip1(i_i2c_p_det_intr), .ip2(i_i2c_p_det_flg), .op(n4162) );
  inv_1 U12513 ( .ip(n11086), .op(n11088) );
  mux2_1 U12514 ( .ip1(i_i2c_rx_addr_10bit), .ip2(n11088), .s(n11087), .op(
        n5086) );
  xor2_1 U12515 ( .ip1(i_i2c_s_det), .ip2(i_i2c_s_det_flg), .op(n4171) );
  xor2_1 U12516 ( .ip1(i_i2c_tx_pop), .ip2(i_i2c_tx_pop_flg), .op(n4173) );
  nor2_1 U12517 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_hs_sync_inv), .ip2(n11093), 
        .op(n11089) );
  xor2_1 U12518 ( .ip1(i_i2c_tx_abrt_source[8]), .ip2(n11089), .op(n4856) );
  nor2_1 U12519 ( .ip1(n11091), .ip2(n11090), .op(n11092) );
  xor2_1 U12520 ( .ip1(i_i2c_tx_abrt_source[11]), .ip2(n11092), .op(n4855) );
  nor2_1 U12521 ( .ip1(n11094), .ip2(n11093), .op(n11095) );
  xor2_1 U12522 ( .ip1(i_i2c_tx_abrt_source[9]), .ip2(n11095), .op(n4854) );
  xor2_1 U12523 ( .ip1(i_i2c_tx_abrt_source[12]), .ip2(n11096), .op(n4175) );
  mux2_1 U12524 ( .ip1(i_apb_pwdata_int[10]), .ip2(i_ssi_ctrlr0[10]), .s(
        n11097), .op(n4590) );
  mux2_1 U12525 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[23]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[23]), .s(n11107), .op(n4792) );
  nand2_1 U12526 ( .ip1(n5592), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[23]), .op(n11100) );
  nand2_1 U12527 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[23]), 
        .op(n11099) );
  nand2_1 U12528 ( .ip1(n11117), .ip2(i_apb_pwdata_int[23]), .op(n11098) );
  nand3_1 U12529 ( .ip1(n11100), .ip2(n11099), .ip3(n11098), .op(n4761) );
  mux2_1 U12530 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[22]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[22]), .s(n11107), .op(n4793) );
  nand2_1 U12531 ( .ip1(n5592), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[22]), .op(n11103) );
  nand2_1 U12532 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[22]), 
        .op(n11102) );
  nand2_1 U12533 ( .ip1(n11117), .ip2(i_apb_pwdata_int[22]), .op(n11101) );
  nand3_1 U12534 ( .ip1(n11103), .ip2(n11102), .ip3(n11101), .op(n4762) );
  mux2_1 U12535 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[21]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[21]), .s(n11107), .op(n4794) );
  nand2_1 U12536 ( .ip1(n5592), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[21]), .op(n11106) );
  nand2_1 U12537 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[21]), 
        .op(n11105) );
  nand2_1 U12538 ( .ip1(n11117), .ip2(i_apb_pwdata_int[21]), .op(n11104) );
  nand3_1 U12539 ( .ip1(n11106), .ip2(n11105), .ip3(n11104), .op(n4763) );
  mux2_1 U12540 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[20]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[20]), .s(n11107), .op(n4795) );
  nand2_1 U12541 ( .ip1(n5592), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[20]), .op(n11110) );
  nand2_1 U12542 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[20]), 
        .op(n11109) );
  nand2_1 U12543 ( .ip1(n11117), .ip2(i_apb_pwdata_int[20]), .op(n11108) );
  nand3_1 U12544 ( .ip1(n11110), .ip2(n11109), .ip3(n11108), .op(n4764) );
  mux2_1 U12545 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[19]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[19]), .s(n11121), .op(n4796) );
  nand2_1 U12546 ( .ip1(n5592), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[19]), .op(n11113) );
  nand2_1 U12547 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[19]), 
        .op(n11112) );
  nand2_1 U12548 ( .ip1(n11117), .ip2(i_apb_pwdata_int[19]), .op(n11111) );
  nand3_1 U12549 ( .ip1(n11113), .ip2(n11112), .ip3(n11111), .op(n4765) );
  mux2_1 U12550 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[18]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[18]), .s(n11121), .op(n4797) );
  nand2_1 U12551 ( .ip1(n5592), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[18]), .op(n11116) );
  nand2_1 U12552 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[18]), 
        .op(n11115) );
  nand2_1 U12553 ( .ip1(n11117), .ip2(i_apb_pwdata_int[18]), .op(n11114) );
  nand3_1 U12554 ( .ip1(n11116), .ip2(n11115), .ip3(n11114), .op(n4766) );
  mux2_1 U12555 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[17]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[17]), .s(n11121), .op(n4798) );
  nand2_1 U12556 ( .ip1(n5592), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[17]), .op(n11120) );
  nand2_1 U12557 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[17]), 
        .op(n11119) );
  nand2_1 U12558 ( .ip1(n11117), .ip2(i_apb_pwdata_int[17]), .op(n11118) );
  nand3_1 U12559 ( .ip1(n11120), .ip2(n11119), .ip3(n11118), .op(n4767) );
  mux2_1 U12560 ( .ip1(i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[16]), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[16]), .s(n11121), .op(n4799) );
  nand2_1 U12561 ( .ip1(n5592), .ip2(
        i_apb_U_DW_apb_ahbsif_saved_hwdata32_c[16]), .op(n11125) );
  nand2_1 U12562 ( .ip1(n11122), .ip2(ex_i_ahb_AHB_MASTER_CORTEXM0_hwdata[16]), 
        .op(n11124) );
  nand2_1 U12563 ( .ip1(n11117), .ip2(i_apb_pwdata_int[16]), .op(n11123) );
  nand3_1 U12564 ( .ip1(n11125), .ip2(n11124), .ip3(n11123), .op(n4768) );
  nand4_1 U12565 ( .ip1(n11126), .ip2(i_i2c_ic_abort_sync), .ip3(
        i_i2c_U_DW_apb_i2c_mstfsm_ic_abort_chk_win), .ip4(
        i_i2c_U_DW_apb_i2c_mstfsm_byte_waiting_q), .op(n11129) );
  nand2_1 U12566 ( .ip1(n11127), .ip2(i_i2c_abrt_in_rcve_trns), .op(n11128) );
  nand2_1 U12567 ( .ip1(n11129), .ip2(n11128), .op(n5183) );
  xor2_1 U12570 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_rx_push_flg_sync), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_rx_push_flg_sync_q), .op(i_i2c_rx_push_sync)
         );
  inv_1 U12571 ( .ip(i_i2c_rx_pop), .op(n11182) );
  nor2_1 U12572 ( .ip1(n11182), .ip2(n5240), .op(n11163) );
  inv_1 U12573 ( .ip(i_i2c_rx_push_sync), .op(n11181) );
  nand2_1 U12574 ( .ip1(n11163), .ip2(n11181), .op(n11183) );
  inv_1 U12575 ( .ip(n11183), .op(n11132) );
  inv_1 U12576 ( .ip(i_i2c_rx_full), .op(n11137) );
  nand2_1 U12577 ( .ip1(n11137), .ip2(n11182), .op(n11179) );
  nand2_1 U12578 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_empty_n), .ip2(
        n11179), .op(n11130) );
  nand2_1 U12579 ( .ip1(i_i2c_rx_push_sync), .ip2(n11130), .op(n11184) );
  mux2_1 U12580 ( .ip1(n11183), .ip2(n11184), .s(
        i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[0]), .op(n11189) );
  inv_1 U12581 ( .ip(i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[0]), .op(n11186)
         );
  nor2_1 U12582 ( .ip1(n11186), .ip2(i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[1]), .op(n11131) );
  not_ab_or_c_or_d U12583 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[1]), 
        .ip2(n11132), .ip3(n11189), .ip4(n11131), .op(n11133) );
  xor2_1 U12584 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[2]), .ip2(n11133), .op(n11198) );
  and2_1 U12585 ( .ip1(i_i2c_fifo_rst_n), .ip2(n11198), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N49) );
  nor2_1 U12586 ( .ip1(i_i2c_rx_pop), .ip2(n11137), .op(n11168) );
  nor2_1 U12587 ( .ip1(i_i2c_rx_push_sync), .ip2(n11168), .op(n11134) );
  inv_1 U12588 ( .ip(i_i2c_fifo_rst_n), .op(n11205) );
  not_ab_or_c_or_d U12589 ( .ip1(n11137), .ip2(n11135), .ip3(n11134), .ip4(
        n11205), .op(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N37) );
  and2_1 U12590 ( .ip1(i_i2c_ic_raw_intr_stat[0]), .ip2(i_i2c_ic_intr_mask[0]), 
        .op(i_i2c_ic_intr_stat[0]) );
  and2_1 U12591 ( .ip1(i_i2c_ic_raw_intr_stat[1]), .ip2(i_i2c_ic_intr_mask[1]), 
        .op(i_i2c_ic_intr_stat[1]) );
  nand3_1 U12592 ( .ip1(i_i2c_ic_rx_tl[0]), .ip2(i_i2c_ic_rx_tl[1]), .ip3(
        i_i2c_ic_rx_tl[2]), .op(n11187) );
  inv_1 U12593 ( .ip(n11187), .op(n11138) );
  nor2_1 U12594 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_i_rx_almost_full), .ip2(n11138), 
        .op(n11136) );
  not_ab_or_c_or_d U12595 ( .ip1(n11138), .ip2(n11137), .ip3(n11136), .ip4(
        n11449), .op(i_i2c_ic_raw_intr_stat[2]) );
  and2_1 U12596 ( .ip1(i_i2c_ic_raw_intr_stat[2]), .ip2(i_i2c_ic_intr_mask[2]), 
        .op(i_i2c_ic_intr_stat[2]) );
  and2_1 U12597 ( .ip1(i_i2c_ic_raw_intr_stat[3]), .ip2(i_i2c_ic_intr_mask[3]), 
        .op(i_i2c_ic_intr_stat[3]) );
  inv_1 U12598 ( .ip(i_i2c_ic_tx_tl[2]), .op(n11146) );
  inv_1 U12599 ( .ip(i_i2c_ic_tx_tl[0]), .op(n11139) );
  nand2_1 U12600 ( .ip1(n11139), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[0]), .op(n11144) );
  nand2_1 U12601 ( .ip1(n11140), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[1]), .op(n11143) );
  nor2_1 U12602 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[1]), .ip2(
        n11140), .op(n11142) );
  nor2_1 U12603 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[2]), .ip2(
        n11146), .op(n11141) );
  not_ab_or_c_or_d U12604 ( .ip1(n11144), .ip2(n11143), .ip3(n11142), .ip4(
        n11141), .op(n11145) );
  not_ab_or_c_or_d U12605 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[2]), 
        .ip2(n11146), .ip3(n11145), .ip4(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[3]), .op(n11148) );
  nor4_1 U12606 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[6]), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[7]), .ip3(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[5]), .ip4(
        i_i2c_U_DW_apb_i2c_fifo_tx_fifo_cmd_cntr[4]), .op(n11147) );
  nand2_1 U12607 ( .ip1(n11148), .ip2(n11147), .op(n11149) );
  mux2_1 U12608 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_almost_empty_n), 
        .ip2(n11149), .s(i_i2c_tx_empty_ctrl), .op(n11150) );
  nor2_1 U12609 ( .ip1(n11449), .ip2(n11150), .op(i_i2c_ic_raw_intr_stat[4])
         );
  and2_1 U12610 ( .ip1(i_i2c_ic_raw_intr_stat[4]), .ip2(i_i2c_ic_intr_mask[4]), 
        .op(i_i2c_ic_intr_stat[4]) );
  and2_1 U12611 ( .ip1(i_i2c_ic_raw_intr_stat[5]), .ip2(i_i2c_ic_intr_mask[5]), 
        .op(i_i2c_ic_intr_stat[5]) );
  and2_1 U12612 ( .ip1(i_i2c_ic_raw_intr_stat[6]), .ip2(i_i2c_ic_intr_mask[6]), 
        .op(i_i2c_ic_intr_stat[6]) );
  and2_1 U12613 ( .ip1(i_i2c_ic_raw_intr_stat[7]), .ip2(i_i2c_ic_intr_mask[7]), 
        .op(i_i2c_ic_intr_stat[7]) );
  and2_1 U12614 ( .ip1(i_i2c_ic_raw_intr_stat[8]), .ip2(i_i2c_ic_intr_mask[8]), 
        .op(i_i2c_ic_intr_stat[8]) );
  and2_1 U12615 ( .ip1(i_i2c_ic_raw_intr_stat[9]), .ip2(i_i2c_ic_intr_mask[9]), 
        .op(i_i2c_ic_intr_stat[9]) );
  and2_1 U12616 ( .ip1(i_i2c_ic_raw_intr_stat[10]), .ip2(
        i_i2c_ic_intr_mask[10]), .op(i_i2c_ic_intr_stat[10]) );
  and2_1 U12617 ( .ip1(i_i2c_ic_raw_intr_stat[11]), .ip2(
        i_i2c_ic_intr_mask[11]), .op(i_i2c_ic_intr_stat[11]) );
  or2_1 U12618 ( .ip1(i_i2c_ic_enable[0]), .ip2(i_i2c_activity), .op(
        i_i2c_U_DW_apb_i2c_intctl_N4) );
  nand3_1 U12619 ( .ip1(i_apb_penable), .ip2(i_apb_psel_en), .ip3(i_apb_pwrite), .op(n11151) );
  nor3_1 U12620 ( .ip1(i_apb_paddr[12]), .ip2(n11152), .ip3(n11151), .op(
        i_i2c_wr_en) );
  nand2_1 U12621 ( .ip1(ex_i_ahb_AHB_Slave_PID_hresp[1]), .ip2(
        i_ahb_U_mux_hsel_prev[4]), .op(n11157) );
  nand2_1 U12622 ( .ip1(n11153), .ip2(ex_i_ahb_AHB_Slave_PWM_hresp[1]), .op(
        n11156) );
  nand2_1 U12623 ( .ip1(n11154), .ip2(ex_i_ahb_AHB_Slave_RAM_hresp[1]), .op(
        n11155) );
  nand3_1 U12624 ( .ip1(n11157), .ip2(n11156), .ip3(n11155), .op(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hresp[1]) );
  nor2_1 U12625 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[16]), .ip2(n11158), 
        .op(ex_i_ahb_AHB_Slave_RAM_hsel) );
  inv_1 U12626 ( .ip(ex_i_ahb_AHB_Slave_RAM_hsel), .op(n11159) );
  nand4_1 U12627 ( .ip1(n11160), .ip2(n11159), .ip3(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hready), .ip4(
        ex_i_ahb_AHB_MASTER_CORTEXM0_htrans[1]), .op(n11161) );
  nand2_1 U12628 ( .ip1(n6677), .ip2(n11161), .op(i_ahb_U_dfltslv_N4) );
  nor2_1 U12629 ( .ip1(n11161), .ip2(i_ahb_U_dfltslv_current_state), .op(
        i_ahb_U_dfltslv_next_state) );
  and3_1 U12630 ( .ip1(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[13]), .ip2(n11162), 
        .ip3(ex_i_ahb_AHB_MASTER_CORTEXM0_haddr[12]), .op(
        ex_i_ahb_AHB_Slave_PID_hsel) );
  inv_1 U12631 ( .ip(i_i2c_rx_rd_addr[1]), .op(n11704) );
  nand2_1 U12632 ( .ip1(n11163), .ip2(i_i2c_rx_rd_addr[0]), .op(n11175) );
  inv_1 U12633 ( .ip(n11163), .op(n11178) );
  nand2_1 U12634 ( .ip1(i_i2c_rx_rd_addr[1]), .ip2(i_i2c_rx_rd_addr[0]), .op(
        n11702) );
  nor2_1 U12635 ( .ip1(n11178), .ip2(n11702), .op(n11166) );
  nand2_1 U12636 ( .ip1(n11163), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_rd_addr_at_max), .op(n11164) );
  nand2_1 U12637 ( .ip1(i_i2c_fifo_rst_n), .ip2(n11164), .op(n11176) );
  not_ab_or_c_or_d U12638 ( .ip1(n11704), .ip2(n11175), .ip3(n11166), .ip4(
        n11176), .op(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N45) );
  nor2_1 U12639 ( .ip1(i_i2c_rx_rd_addr[2]), .ip2(n11166), .op(n11165) );
  not_ab_or_c_or_d U12640 ( .ip1(i_i2c_rx_rd_addr[2]), .ip2(n11166), .ip3(
        n11165), .ip4(n11176), .op(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N46) );
  inv_1 U12641 ( .ip(i_i2c_rx_wr_addr[0]), .op(n11174) );
  nor3_1 U12642 ( .ip1(n11168), .ip2(n11181), .ip3(n11174), .op(n11335) );
  inv_1 U12643 ( .ip(n11335), .op(n11336) );
  inv_1 U12644 ( .ip(i_i2c_rx_wr_addr[1]), .op(n11338) );
  nor2_1 U12645 ( .ip1(n11168), .ip2(n11181), .op(n11172) );
  nand2_1 U12646 ( .ip1(n11172), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_wr_addr_at_max), .op(n11169) );
  nand2_1 U12647 ( .ip1(i_i2c_fifo_rst_n), .ip2(n11169), .op(n11173) );
  not_ab_or_c_or_d U12648 ( .ip1(n11336), .ip2(n11338), .ip3(n11167), .ip4(
        n11173), .op(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N42) );
  nor3_1 U12649 ( .ip1(i_i2c_rx_wr_addr[2]), .ip2(n11338), .ip3(n11336), .op(
        n11344) );
  or2_1 U12650 ( .ip1(i_i2c_rx_wr_addr[2]), .ip2(n11344), .op(n11170) );
  nand3_1 U12651 ( .ip1(n11335), .ip2(i_i2c_rx_wr_addr[1]), .ip3(
        i_i2c_rx_wr_addr[2]), .op(n11340) );
  nand2_1 U12652 ( .ip1(n11170), .ip2(n11340), .op(n11171) );
  nor2_1 U12653 ( .ip1(n11171), .ip2(n11173), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N43) );
  inv_1 U12654 ( .ip(n11172), .op(n11334) );
  not_ab_or_c_or_d U12655 ( .ip1(n11334), .ip2(n11174), .ip3(n11335), .ip4(
        n11173), .op(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N41) );
  and3_1 U12656 ( .ip1(i_i2c_rx_wr_addr[1]), .ip2(i_i2c_rx_wr_addr[2]), .ip3(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N41), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N40) );
  inv_1 U12657 ( .ip(i_i2c_rx_rd_addr[0]), .op(n11701) );
  inv_1 U12658 ( .ip(n11175), .op(n11177) );
  not_ab_or_c_or_d U12659 ( .ip1(n11178), .ip2(n11701), .ip3(n11177), .ip4(
        n11176), .op(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N44) );
  and3_1 U12660 ( .ip1(i_i2c_rx_rd_addr[2]), .ip2(i_i2c_rx_rd_addr[1]), .ip3(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N44), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N39) );
  nand2_1 U12661 ( .ip1(n11179), .ip2(n11178), .op(n11180) );
  not_ab_or_c_or_d U12662 ( .ip1(n11182), .ip2(n11181), .ip3(n11205), .ip4(
        n11180), .op(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N38) );
  inv_1 U12663 ( .ip(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N37), .op(n11204) );
  and2_1 U12664 ( .ip1(n11184), .ip2(n11183), .op(n11185) );
  mux2_1 U12665 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[0]), .ip2(n11186), .s(n11185), .op(n11206) );
  nand2_1 U12666 ( .ip1(i_i2c_ic_rx_tl[0]), .ip2(n11187), .op(n11188) );
  nand2_1 U12667 ( .ip1(n11206), .ip2(n11188), .op(n11193) );
  inv_1 U12668 ( .ip(i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[1]), .op(n11190)
         );
  mux2_1 U12669 ( .ip1(n11190), .ip2(i_i2c_U_DW_apb_i2c_fifo_wrdc_rx_unconn[1]), .s(n11189), .op(n11207) );
  nor2_1 U12670 ( .ip1(n11193), .ip2(n11207), .op(n11195) );
  nor2_1 U12671 ( .ip1(i_i2c_ic_rx_tl[0]), .ip2(i_i2c_ic_rx_tl[1]), .op(n11192) );
  nand2_1 U12672 ( .ip1(i_i2c_ic_rx_tl[0]), .ip2(i_i2c_ic_rx_tl[1]), .op(
        n11196) );
  nor2_1 U12673 ( .ip1(i_i2c_ic_rx_tl[2]), .ip2(n11196), .op(n11191) );
  not_ab_or_c_or_d U12674 ( .ip1(n11207), .ip2(n11193), .ip3(n11192), .ip4(
        n11191), .op(n11194) );
  or2_1 U12675 ( .ip1(n11195), .ip2(n11194), .op(n11202) );
  inv_1 U12676 ( .ip(n11196), .op(n11197) );
  nor2_1 U12677 ( .ip1(i_i2c_ic_rx_tl[2]), .ip2(n11197), .op(n11199) );
  nand2_1 U12678 ( .ip1(n11199), .ip2(n11198), .op(n11201) );
  nor2_1 U12679 ( .ip1(n11199), .ip2(n11198), .op(n11200) );
  ab_or_c_or_d U12680 ( .ip1(n11202), .ip2(n11201), .ip3(n11205), .ip4(n11200), 
        .op(n11203) );
  nand2_1 U12681 ( .ip1(n11204), .ip2(n11203), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N36) );
  nor2_1 U12682 ( .ip1(n11206), .ip2(n11205), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N47) );
  and2_1 U12683 ( .ip1(n11207), .ip2(i_i2c_fifo_rst_n), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N48) );
  or4_1 U12684 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N37), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N47), .ip3(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N48), .ip4(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N49), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_rx_fifo_N33) );
  nand2_1 U12685 ( .ip1(n11215), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_rd_addr_at_max), .op(n11208) );
  nand2_1 U12686 ( .ip1(i_i2c_tx_fifo_rst_n), .ip2(n11208), .op(n11225) );
  nor2_1 U12687 ( .ip1(n11209), .ip2(n11227), .op(n11212) );
  nor2_1 U12688 ( .ip1(n11228), .ip2(n11227), .op(n11226) );
  nor2_1 U12689 ( .ip1(i_i2c_tx_rd_addr[1]), .ip2(n11226), .op(n11210) );
  nor2_1 U12690 ( .ip1(n11212), .ip2(n11210), .op(n11229) );
  inv_1 U12691 ( .ip(n11229), .op(n11211) );
  nor2_1 U12692 ( .ip1(n11225), .ip2(n11211), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N45) );
  nor2_1 U12693 ( .ip1(i_i2c_tx_rd_addr[2]), .ip2(n11212), .op(n11213) );
  not_ab_or_c_or_d U12694 ( .ip1(n11215), .ip2(n11214), .ip3(n11213), .ip4(
        n11225), .op(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N46) );
  inv_1 U12695 ( .ip(i_i2c_tx_wr_addr[1]), .op(n11323) );
  inv_1 U12696 ( .ip(i_i2c_tx_wr_addr[0]), .op(n11223) );
  nand2_1 U12697 ( .ip1(i_i2c_tx_full), .ip2(n11216), .op(n11217) );
  nand2_1 U12698 ( .ip1(i_i2c_tx_push), .ip2(n11217), .op(n11325) );
  nor2_1 U12699 ( .ip1(n11223), .ip2(n11325), .op(n11222) );
  inv_1 U12700 ( .ip(n11222), .op(n11324) );
  nand2_1 U12701 ( .ip1(i_i2c_tx_wr_addr[1]), .ip2(n11222), .op(n11322) );
  inv_1 U12702 ( .ip(n11322), .op(n11220) );
  inv_1 U12703 ( .ip(n11325), .op(n11218) );
  nand2_1 U12704 ( .ip1(n11218), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_wr_addr_at_max), .op(n11219) );
  nand2_1 U12705 ( .ip1(i_i2c_tx_fifo_rst_n), .ip2(n11219), .op(n11221) );
  not_ab_or_c_or_d U12706 ( .ip1(n11323), .ip2(n11324), .ip3(n11220), .ip4(
        n11221), .op(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N42) );
  inv_1 U12707 ( .ip(i_i2c_tx_wr_addr[2]), .op(n11321) );
  nand2_1 U12708 ( .ip1(i_i2c_tx_wr_addr[2]), .ip2(i_i2c_tx_wr_addr[1]), .op(
        n11320) );
  nor2_1 U12709 ( .ip1(n11324), .ip2(n11320), .op(n11326) );
  not_ab_or_c_or_d U12710 ( .ip1(n11321), .ip2(n11322), .ip3(n11326), .ip4(
        n11221), .op(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N43) );
  not_ab_or_c_or_d U12711 ( .ip1(n11223), .ip2(n11325), .ip3(n11222), .ip4(
        n11221), .op(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N41) );
  inv_1 U12712 ( .ip(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N41), .op(n11224) );
  nor2_1 U12713 ( .ip1(n11320), .ip2(n11224), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N40) );
  not_ab_or_c_or_d U12714 ( .ip1(n11228), .ip2(n11227), .ip3(n11226), .ip4(
        n11225), .op(i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N44) );
  and3_1 U12715 ( .ip1(i_i2c_tx_rd_addr[2]), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N44), .ip3(n11229), .op(
        i_i2c_U_DW_apb_i2c_fifo_U_tx_fifo_N39) );
  inv_1 U12716 ( .ip(n11230), .op(n11231) );
  nor3_1 U12717 ( .ip1(i_i2c_U_DW_apb_i2c_sync_ic_10bit_slv_sync_inv), .ip2(
        n11232), .ip3(n11231), .op(n11234) );
  not_ab_or_c_or_d U12718 ( .ip1(n11235), .ip2(n11288), .ip3(n11234), .ip4(
        n11233), .op(n11237) );
  nor2_1 U12719 ( .ip1(n11237), .ip2(n11236), .op(
        i_i2c_U_DW_apb_i2c_slvfsm_N37) );
  and2_1 U12720 ( .ip1(n11311), .ip2(n11238), .op(
        i_i2c_U_DW_apb_i2c_rx_shift_rx_slv_read_s) );
  and2_1 U12721 ( .ip1(n11244), .ip2(n11239), .op(n11241) );
  nor2_1 U12722 ( .ip1(n11241), .ip2(n11240), .op(n11246) );
  inv_1 U12723 ( .ip(n11242), .op(n11243) );
  and4_1 U12724 ( .ip1(n11244), .ip2(i_i2c_U_DW_apb_i2c_slvfsm_slv_tx_flush), 
        .ip3(n11243), .ip4(n11280), .op(n11245) );
  or2_1 U12725 ( .ip1(n11246), .ip2(n11245), .op(n5223) );
  or2_1 U12726 ( .ip1(i_i2c_ic_clr_intr_en), .ip2(i_i2c_ic_clr_tx_abrt_en), 
        .op(n11247) );
  nand2_1 U12727 ( .ip1(n11839), .ip2(n11247), .op(n11433) );
  inv_1 U12728 ( .ip(n11433), .op(n11400) );
  inv_1 U12729 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[16]), .op(
        n11249) );
  nor2_1 U12730 ( .ip1(n11249), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[16]), .op(n11248) );
  not_ab_or_c_or_d U12731 ( .ip1(n11249), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[16]), .ip3(
        i_i2c_ic_tx_abrt_source[16]), .ip4(n11248), .op(n11250) );
  nor2_1 U12732 ( .ip1(n11400), .ip2(n11250), .op(n5212) );
  nor3_1 U12733 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[1]), .ip2(
        n11280), .ip3(n11251), .op(n11257) );
  or2_1 U12734 ( .ip1(n11253), .ip2(n11252), .op(n11255) );
  nor2_1 U12735 ( .ip1(n11280), .ip2(n11254), .op(n11286) );
  inv_1 U12736 ( .ip(n11286), .op(n11274) );
  nand2_1 U12737 ( .ip1(n11255), .ip2(n11274), .op(n11256) );
  or2_1 U12738 ( .ip1(n11257), .ip2(n11256), .op(n5210) );
  nor2_1 U12739 ( .ip1(n11264), .ip2(n11280), .op(n11258) );
  or2_1 U12740 ( .ip1(n11279), .ip2(n11258), .op(n11262) );
  nand2_1 U12741 ( .ip1(n11262), .ip2(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[2]), .op(n11261) );
  nand4_1 U12742 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[0]), .ip2(
        n11272), .ip3(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[1]), .ip4(
        n11259), .op(n11260) );
  nand3_1 U12743 ( .ip1(n11261), .ip2(n11260), .ip3(n11274), .op(n5209) );
  nand2_1 U12744 ( .ip1(n11262), .ip2(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[3]), .op(n11266) );
  inv_1 U12745 ( .ip(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[3]), .op(
        n11263) );
  nand3_1 U12746 ( .ip1(n11264), .ip2(n11272), .ip3(n11263), .op(n11265) );
  nand3_1 U12747 ( .ip1(n11266), .ip2(n11265), .ip3(n11274), .op(n5208) );
  nor2_1 U12748 ( .ip1(n11273), .ip2(n11280), .op(n11267) );
  or2_1 U12749 ( .ip1(n11279), .ip2(n11267), .op(n11270) );
  nor3_1 U12750 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[4]), .ip2(
        n11268), .ip3(n11280), .op(n11269) );
  ab_or_c_or_d U12751 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[4]), 
        .ip2(n11270), .ip3(n11286), .ip4(n11269), .op(n5207) );
  nand2_1 U12752 ( .ip1(n11270), .ip2(
        i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[5]), .op(n11276) );
  inv_1 U12753 ( .ip(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[5]), .op(
        n11271) );
  nand3_1 U12754 ( .ip1(n11273), .ip2(n11272), .ip3(n11271), .op(n11275) );
  nand3_1 U12755 ( .ip1(n11276), .ip2(n11275), .ip3(n11274), .op(n5206) );
  nor2_1 U12756 ( .ip1(n11277), .ip2(n11280), .op(n11278) );
  or2_1 U12757 ( .ip1(n11279), .ip2(n11278), .op(n11287) );
  nor3_1 U12758 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[6]), .ip2(
        n11284), .ip3(n11280), .op(n11281) );
  ab_or_c_or_d U12759 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[6]), 
        .ip2(n11287), .ip3(n11286), .ip4(n11281), .op(n5205) );
  nor3_1 U12760 ( .ip1(n11284), .ip2(n11283), .ip3(n11282), .op(n11285) );
  ab_or_c_or_d U12761 ( .ip1(i_i2c_U_DW_apb_i2c_slvfsm_stretch_scl_count[7]), 
        .ip2(n11287), .ip3(n11286), .ip4(n11285), .op(n5204) );
  nor3_1 U12762 ( .ip1(i_i2c_slv_rx_aborted), .ip2(n11289), .ip3(n11288), .op(
        n11290) );
  nor2_1 U12763 ( .ip1(i_i2c_ic_enable_sync), .ip2(n11290), .op(n5203) );
  inv_1 U12764 ( .ip(i_i2c_U_DW_apb_i2c_toggle_tx_abrt), .op(n11291) );
  nor2_1 U12765 ( .ip1(i_i2c_U_DW_apb_i2c_toggle_tx_abrt_r), .ip2(n11291), 
        .op(n11292) );
  inv_1 U12766 ( .ip(i_i2c_tx_abrt_source[15]), .op(n11295) );
  nand2_1 U12767 ( .ip1(i_i2c_tx_fifo_data_buf[8]), .ip2(n11293), .op(n11294)
         );
  mux2_1 U12768 ( .ip1(n11295), .ip2(i_i2c_tx_abrt_source[15]), .s(n11294), 
        .op(n5111) );
  nor2_1 U12769 ( .ip1(n11673), .ip2(n11296), .op(n11297) );
  nor2_1 U12770 ( .ip1(i_i2c_slv_fifo_filled_and_flushed), .ip2(n11297), .op(
        n11298) );
  nor2_1 U12771 ( .ip1(i_i2c_ic_enable_sync), .ip2(n11298), .op(n5079) );
  nor3_1 U12772 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[1]), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[2]), .ip3(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[3]), .op(n11300) );
  nor3_1 U12773 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[0]), .ip2(
        n11300), .ip3(n11299), .op(n11308) );
  inv_1 U12774 ( .ip(n11308), .op(n11303) );
  nand2_1 U12775 ( .ip1(n11301), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[0]), .op(n11302) );
  nand2_1 U12776 ( .ip1(n11303), .ip2(n11302), .op(n5077) );
  nand2_1 U12777 ( .ip1(n11305), .ip2(n11304), .op(n11306) );
  nand3_1 U12778 ( .ip1(n11311), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[1]), .ip3(n11306), .op(
        n11309) );
  nand2_1 U12779 ( .ip1(n11308), .ip2(n11307), .op(n11310) );
  nand2_1 U12780 ( .ip1(n11309), .ip2(n11310), .op(n5076) );
  nand3_1 U12781 ( .ip1(n11311), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[2]), .ip3(n11310), .op(
        n11313) );
  nand2_1 U12782 ( .ip1(n11313), .ip2(n11312), .op(n5075) );
  xor2_1 U12783 ( .ip1(n11315), .ip2(i_i2c_rx_done_flg), .op(n5064) );
  xor2_1 U12784 ( .ip1(i_i2c_tx_abrt_source[13]), .ip2(n11314), .op(n5032) );
  inv_1 U12785 ( .ip(n11315), .op(n11316) );
  nor2_1 U12786 ( .ip1(n11861), .ip2(n11316), .op(n11317) );
  xor2_1 U12787 ( .ip1(n11317), .ip2(i_i2c_slv_clr_leftover_flg), .op(n5031)
         );
  mux2_1 U12788 ( .ip1(n11319), .ip2(n11318), .s(i_i2c_ic_rd_req_flg), .op(
        n5030) );
  mux2_1 U12789 ( .ip1(i_i2c_U_dff_tx_mem[0]), .ip2(i_apb_pwdata_int[0]), .s(
        n11326), .op(n5028) );
  nor3_1 U12790 ( .ip1(i_i2c_tx_wr_addr[0]), .ip2(n11325), .ip3(n11320), .op(
        n11327) );
  mux2_1 U12791 ( .ip1(i_i2c_U_dff_tx_mem[9]), .ip2(i_apb_pwdata_int[0]), .s(
        n11327), .op(n5027) );
  nor3_1 U12792 ( .ip1(i_i2c_tx_wr_addr[1]), .ip2(n11321), .ip3(n11324), .op(
        n11328) );
  mux2_1 U12793 ( .ip1(i_i2c_U_dff_tx_mem[18]), .ip2(i_apb_pwdata_int[0]), .s(
        n11328), .op(n5026) );
  mux2_1 U12794 ( .ip1(i_i2c_U_dff_tx_mem[27]), .ip2(i_apb_pwdata_int[0]), .s(
        n11329), .op(n5025) );
  nor2_1 U12795 ( .ip1(i_i2c_tx_wr_addr[2]), .ip2(n11322), .op(n11330) );
  mux2_1 U12796 ( .ip1(i_i2c_U_dff_tx_mem[36]), .ip2(i_apb_pwdata_int[0]), .s(
        n11330), .op(n5024) );
  mux2_1 U12797 ( .ip1(i_i2c_U_dff_tx_mem[45]), .ip2(i_apb_pwdata_int[0]), .s(
        n11331), .op(n5023) );
  nor3_1 U12798 ( .ip1(i_i2c_tx_wr_addr[2]), .ip2(i_i2c_tx_wr_addr[1]), .ip3(
        n11324), .op(n11332) );
  mux2_1 U12799 ( .ip1(i_i2c_U_dff_tx_mem[54]), .ip2(i_apb_pwdata_int[0]), .s(
        n11332), .op(n5022) );
  mux2_1 U12800 ( .ip1(i_i2c_U_dff_tx_mem[63]), .ip2(i_apb_pwdata_int[0]), .s(
        n11333), .op(n5021) );
  mux2_1 U12801 ( .ip1(i_i2c_U_dff_tx_mem[1]), .ip2(i_apb_pwdata_int[1]), .s(
        n11326), .op(n5020) );
  mux2_1 U12802 ( .ip1(i_i2c_U_dff_tx_mem[10]), .ip2(i_apb_pwdata_int[1]), .s(
        n11327), .op(n5019) );
  mux2_1 U12803 ( .ip1(i_i2c_U_dff_tx_mem[19]), .ip2(i_apb_pwdata_int[1]), .s(
        n11328), .op(n5018) );
  mux2_1 U12804 ( .ip1(i_i2c_U_dff_tx_mem[28]), .ip2(i_apb_pwdata_int[1]), .s(
        n11329), .op(n5017) );
  mux2_1 U12805 ( .ip1(i_i2c_U_dff_tx_mem[37]), .ip2(i_apb_pwdata_int[1]), .s(
        n11330), .op(n5016) );
  mux2_1 U12806 ( .ip1(i_i2c_U_dff_tx_mem[46]), .ip2(i_apb_pwdata_int[1]), .s(
        n11331), .op(n5015) );
  mux2_1 U12807 ( .ip1(i_i2c_U_dff_tx_mem[55]), .ip2(i_apb_pwdata_int[1]), .s(
        n11332), .op(n5014) );
  mux2_1 U12808 ( .ip1(i_i2c_U_dff_tx_mem[64]), .ip2(i_apb_pwdata_int[1]), .s(
        n11333), .op(n5013) );
  mux2_1 U12809 ( .ip1(i_i2c_U_dff_tx_mem[2]), .ip2(i_apb_pwdata_int[2]), .s(
        n11326), .op(n5012) );
  mux2_1 U12810 ( .ip1(i_i2c_U_dff_tx_mem[11]), .ip2(i_apb_pwdata_int[2]), .s(
        n11327), .op(n5011) );
  mux2_1 U12811 ( .ip1(i_i2c_U_dff_tx_mem[20]), .ip2(i_apb_pwdata_int[2]), .s(
        n11328), .op(n5010) );
  mux2_1 U12812 ( .ip1(i_i2c_U_dff_tx_mem[29]), .ip2(i_apb_pwdata_int[2]), .s(
        n11329), .op(n5009) );
  mux2_1 U12813 ( .ip1(i_i2c_U_dff_tx_mem[38]), .ip2(i_apb_pwdata_int[2]), .s(
        n11330), .op(n5008) );
  mux2_1 U12814 ( .ip1(i_i2c_U_dff_tx_mem[47]), .ip2(i_apb_pwdata_int[2]), .s(
        n11331), .op(n5007) );
  mux2_1 U12815 ( .ip1(i_i2c_U_dff_tx_mem[56]), .ip2(i_apb_pwdata_int[2]), .s(
        n11332), .op(n5006) );
  mux2_1 U12816 ( .ip1(i_i2c_U_dff_tx_mem[65]), .ip2(i_apb_pwdata_int[2]), .s(
        n11333), .op(n5005) );
  mux2_1 U12817 ( .ip1(i_i2c_U_dff_tx_mem[3]), .ip2(i_apb_pwdata_int[3]), .s(
        n11326), .op(n5004) );
  mux2_1 U12818 ( .ip1(i_i2c_U_dff_tx_mem[12]), .ip2(i_apb_pwdata_int[3]), .s(
        n11327), .op(n5003) );
  mux2_1 U12819 ( .ip1(i_i2c_U_dff_tx_mem[21]), .ip2(i_apb_pwdata_int[3]), .s(
        n11328), .op(n5002) );
  mux2_1 U12820 ( .ip1(i_i2c_U_dff_tx_mem[30]), .ip2(i_apb_pwdata_int[3]), .s(
        n11329), .op(n5001) );
  mux2_1 U12821 ( .ip1(i_i2c_U_dff_tx_mem[39]), .ip2(i_apb_pwdata_int[3]), .s(
        n11330), .op(n5000) );
  mux2_1 U12822 ( .ip1(i_i2c_U_dff_tx_mem[48]), .ip2(i_apb_pwdata_int[3]), .s(
        n11331), .op(n4999) );
  mux2_1 U12823 ( .ip1(i_i2c_U_dff_tx_mem[57]), .ip2(i_apb_pwdata_int[3]), .s(
        n11332), .op(n4998) );
  mux2_1 U12824 ( .ip1(i_i2c_U_dff_tx_mem[66]), .ip2(i_apb_pwdata_int[3]), .s(
        n11333), .op(n4997) );
  mux2_1 U12825 ( .ip1(i_i2c_U_dff_tx_mem[4]), .ip2(i_apb_pwdata_int[4]), .s(
        n11326), .op(n4996) );
  mux2_1 U12826 ( .ip1(i_i2c_U_dff_tx_mem[13]), .ip2(i_apb_pwdata_int[4]), .s(
        n11327), .op(n4995) );
  mux2_1 U12827 ( .ip1(i_i2c_U_dff_tx_mem[22]), .ip2(i_apb_pwdata_int[4]), .s(
        n11328), .op(n4994) );
  mux2_1 U12828 ( .ip1(i_i2c_U_dff_tx_mem[31]), .ip2(i_apb_pwdata_int[4]), .s(
        n11329), .op(n4993) );
  mux2_1 U12829 ( .ip1(i_i2c_U_dff_tx_mem[40]), .ip2(i_apb_pwdata_int[4]), .s(
        n11330), .op(n4992) );
  mux2_1 U12830 ( .ip1(i_i2c_U_dff_tx_mem[49]), .ip2(i_apb_pwdata_int[4]), .s(
        n11331), .op(n4991) );
  mux2_1 U12831 ( .ip1(i_i2c_U_dff_tx_mem[58]), .ip2(i_apb_pwdata_int[4]), .s(
        n11332), .op(n4990) );
  mux2_1 U12832 ( .ip1(i_i2c_U_dff_tx_mem[67]), .ip2(i_apb_pwdata_int[4]), .s(
        n11333), .op(n4989) );
  mux2_1 U12833 ( .ip1(i_i2c_U_dff_tx_mem[5]), .ip2(i_apb_pwdata_int[5]), .s(
        n11326), .op(n4988) );
  mux2_1 U12834 ( .ip1(i_i2c_U_dff_tx_mem[14]), .ip2(i_apb_pwdata_int[5]), .s(
        n11327), .op(n4987) );
  mux2_1 U12835 ( .ip1(i_i2c_U_dff_tx_mem[23]), .ip2(i_apb_pwdata_int[5]), .s(
        n11328), .op(n4986) );
  mux2_1 U12836 ( .ip1(i_i2c_U_dff_tx_mem[32]), .ip2(i_apb_pwdata_int[5]), .s(
        n11329), .op(n4985) );
  mux2_1 U12837 ( .ip1(i_i2c_U_dff_tx_mem[41]), .ip2(i_apb_pwdata_int[5]), .s(
        n11330), .op(n4984) );
  mux2_1 U12838 ( .ip1(i_i2c_U_dff_tx_mem[50]), .ip2(i_apb_pwdata_int[5]), .s(
        n11331), .op(n4983) );
  mux2_1 U12839 ( .ip1(i_i2c_U_dff_tx_mem[59]), .ip2(i_apb_pwdata_int[5]), .s(
        n11332), .op(n4982) );
  mux2_1 U12840 ( .ip1(i_i2c_U_dff_tx_mem[68]), .ip2(i_apb_pwdata_int[5]), .s(
        n11333), .op(n4981) );
  mux2_1 U12841 ( .ip1(i_i2c_U_dff_tx_mem[6]), .ip2(i_apb_pwdata_int[6]), .s(
        n11326), .op(n4980) );
  mux2_1 U12842 ( .ip1(i_i2c_U_dff_tx_mem[15]), .ip2(i_apb_pwdata_int[6]), .s(
        n11327), .op(n4979) );
  mux2_1 U12843 ( .ip1(i_i2c_U_dff_tx_mem[24]), .ip2(i_apb_pwdata_int[6]), .s(
        n11328), .op(n4978) );
  mux2_1 U12844 ( .ip1(i_i2c_U_dff_tx_mem[33]), .ip2(i_apb_pwdata_int[6]), .s(
        n11329), .op(n4977) );
  mux2_1 U12845 ( .ip1(i_i2c_U_dff_tx_mem[42]), .ip2(i_apb_pwdata_int[6]), .s(
        n11330), .op(n4976) );
  mux2_1 U12846 ( .ip1(i_i2c_U_dff_tx_mem[51]), .ip2(i_apb_pwdata_int[6]), .s(
        n11331), .op(n4975) );
  mux2_1 U12847 ( .ip1(i_i2c_U_dff_tx_mem[60]), .ip2(i_apb_pwdata_int[6]), .s(
        n11332), .op(n4974) );
  mux2_1 U12848 ( .ip1(i_i2c_U_dff_tx_mem[69]), .ip2(i_apb_pwdata_int[6]), .s(
        n11333), .op(n4973) );
  mux2_1 U12849 ( .ip1(i_i2c_U_dff_tx_mem[7]), .ip2(i_apb_pwdata_int[7]), .s(
        n11326), .op(n4972) );
  mux2_1 U12850 ( .ip1(i_i2c_U_dff_tx_mem[16]), .ip2(i_apb_pwdata_int[7]), .s(
        n11327), .op(n4971) );
  mux2_1 U12851 ( .ip1(i_i2c_U_dff_tx_mem[25]), .ip2(i_apb_pwdata_int[7]), .s(
        n11328), .op(n4970) );
  mux2_1 U12852 ( .ip1(i_i2c_U_dff_tx_mem[34]), .ip2(i_apb_pwdata_int[7]), .s(
        n11329), .op(n4969) );
  mux2_1 U12853 ( .ip1(i_i2c_U_dff_tx_mem[43]), .ip2(i_apb_pwdata_int[7]), .s(
        n11330), .op(n4968) );
  mux2_1 U12854 ( .ip1(i_i2c_U_dff_tx_mem[52]), .ip2(i_apb_pwdata_int[7]), .s(
        n11331), .op(n4967) );
  mux2_1 U12855 ( .ip1(i_i2c_U_dff_tx_mem[61]), .ip2(i_apb_pwdata_int[7]), .s(
        n11332), .op(n4966) );
  mux2_1 U12856 ( .ip1(i_i2c_U_dff_tx_mem[70]), .ip2(i_apb_pwdata_int[7]), .s(
        n11333), .op(n4965) );
  mux2_1 U12857 ( .ip1(i_i2c_U_dff_tx_mem[8]), .ip2(i_apb_pwdata_int[8]), .s(
        n11326), .op(n4964) );
  mux2_1 U12858 ( .ip1(i_i2c_U_dff_tx_mem[17]), .ip2(i_apb_pwdata_int[8]), .s(
        n11327), .op(n4963) );
  mux2_1 U12859 ( .ip1(i_i2c_U_dff_tx_mem[26]), .ip2(i_apb_pwdata_int[8]), .s(
        n11328), .op(n4962) );
  mux2_1 U12860 ( .ip1(i_i2c_U_dff_tx_mem[35]), .ip2(i_apb_pwdata_int[8]), .s(
        n11329), .op(n4961) );
  mux2_1 U12861 ( .ip1(i_i2c_U_dff_tx_mem[44]), .ip2(i_apb_pwdata_int[8]), .s(
        n11330), .op(n4960) );
  mux2_1 U12862 ( .ip1(i_i2c_U_dff_tx_mem[53]), .ip2(i_apb_pwdata_int[8]), .s(
        n11331), .op(n4959) );
  mux2_1 U12863 ( .ip1(i_i2c_U_dff_tx_mem[62]), .ip2(i_apb_pwdata_int[8]), .s(
        n11332), .op(n4958) );
  mux2_1 U12864 ( .ip1(i_i2c_U_dff_tx_mem[71]), .ip2(i_apb_pwdata_int[8]), .s(
        n11333), .op(n4957) );
  mux2_1 U12865 ( .ip1(i_i2c_rx_push_data[0]), .ip2(i_i2c_U_dff_rx_mem[0]), 
        .s(n11340), .op(n4921) );
  nor2_1 U12866 ( .ip1(i_i2c_rx_wr_addr[0]), .ip2(n11334), .op(n11339) );
  nand3_1 U12867 ( .ip1(i_i2c_rx_wr_addr[1]), .ip2(i_i2c_rx_wr_addr[2]), .ip3(
        n11339), .op(n11341) );
  mux2_1 U12868 ( .ip1(i_i2c_rx_push_data[0]), .ip2(i_i2c_U_dff_rx_mem[8]), 
        .s(n11341), .op(n4920) );
  nand3_1 U12869 ( .ip1(n11335), .ip2(i_i2c_rx_wr_addr[2]), .ip3(n11338), .op(
        n11342) );
  mux2_1 U12870 ( .ip1(i_i2c_rx_push_data[0]), .ip2(i_i2c_U_dff_rx_mem[16]), 
        .s(n11342), .op(n4919) );
  nand3_1 U12871 ( .ip1(i_i2c_rx_wr_addr[2]), .ip2(n11339), .ip3(n11338), .op(
        n11343) );
  mux2_1 U12872 ( .ip1(i_i2c_rx_push_data[0]), .ip2(i_i2c_U_dff_rx_mem[24]), 
        .s(n11343), .op(n4918) );
  mux2_1 U12873 ( .ip1(i_i2c_U_dff_rx_mem[32]), .ip2(i_i2c_rx_push_data[0]), 
        .s(n11344), .op(n4917) );
  inv_1 U12874 ( .ip(i_i2c_rx_wr_addr[2]), .op(n11337) );
  nand3_1 U12875 ( .ip1(i_i2c_rx_wr_addr[1]), .ip2(n11339), .ip3(n11337), .op(
        n11345) );
  mux2_1 U12876 ( .ip1(i_i2c_rx_push_data[0]), .ip2(i_i2c_U_dff_rx_mem[40]), 
        .s(n11345), .op(n4916) );
  nor3_1 U12877 ( .ip1(i_i2c_rx_wr_addr[1]), .ip2(i_i2c_rx_wr_addr[2]), .ip3(
        n11336), .op(n11346) );
  mux2_1 U12878 ( .ip1(i_i2c_U_dff_rx_mem[48]), .ip2(i_i2c_rx_push_data[0]), 
        .s(n11346), .op(n4915) );
  nand3_1 U12879 ( .ip1(n11339), .ip2(n11338), .ip3(n11337), .op(n11347) );
  mux2_1 U12880 ( .ip1(i_i2c_rx_push_data[0]), .ip2(i_i2c_U_dff_rx_mem[56]), 
        .s(n11347), .op(n4914) );
  mux2_1 U12881 ( .ip1(i_i2c_rx_push_data[1]), .ip2(i_i2c_U_dff_rx_mem[1]), 
        .s(n11340), .op(n4913) );
  mux2_1 U12882 ( .ip1(i_i2c_rx_push_data[1]), .ip2(i_i2c_U_dff_rx_mem[9]), 
        .s(n11341), .op(n4912) );
  mux2_1 U12883 ( .ip1(i_i2c_rx_push_data[1]), .ip2(i_i2c_U_dff_rx_mem[17]), 
        .s(n11342), .op(n4911) );
  mux2_1 U12884 ( .ip1(i_i2c_rx_push_data[1]), .ip2(i_i2c_U_dff_rx_mem[25]), 
        .s(n11343), .op(n4910) );
  mux2_1 U12885 ( .ip1(i_i2c_U_dff_rx_mem[33]), .ip2(i_i2c_rx_push_data[1]), 
        .s(n11344), .op(n4909) );
  mux2_1 U12886 ( .ip1(i_i2c_rx_push_data[1]), .ip2(i_i2c_U_dff_rx_mem[41]), 
        .s(n11345), .op(n4908) );
  mux2_1 U12887 ( .ip1(i_i2c_U_dff_rx_mem[49]), .ip2(i_i2c_rx_push_data[1]), 
        .s(n11346), .op(n4907) );
  mux2_1 U12888 ( .ip1(i_i2c_rx_push_data[1]), .ip2(i_i2c_U_dff_rx_mem[57]), 
        .s(n11347), .op(n4906) );
  mux2_1 U12889 ( .ip1(i_i2c_rx_push_data[2]), .ip2(i_i2c_U_dff_rx_mem[2]), 
        .s(n11340), .op(n4905) );
  mux2_1 U12890 ( .ip1(i_i2c_rx_push_data[2]), .ip2(i_i2c_U_dff_rx_mem[10]), 
        .s(n11341), .op(n4904) );
  mux2_1 U12891 ( .ip1(i_i2c_rx_push_data[2]), .ip2(i_i2c_U_dff_rx_mem[18]), 
        .s(n11342), .op(n4903) );
  mux2_1 U12892 ( .ip1(i_i2c_rx_push_data[2]), .ip2(i_i2c_U_dff_rx_mem[26]), 
        .s(n11343), .op(n4902) );
  mux2_1 U12893 ( .ip1(i_i2c_U_dff_rx_mem[34]), .ip2(i_i2c_rx_push_data[2]), 
        .s(n11344), .op(n4901) );
  mux2_1 U12894 ( .ip1(i_i2c_rx_push_data[2]), .ip2(i_i2c_U_dff_rx_mem[42]), 
        .s(n11345), .op(n4900) );
  mux2_1 U12895 ( .ip1(i_i2c_U_dff_rx_mem[50]), .ip2(i_i2c_rx_push_data[2]), 
        .s(n11346), .op(n4899) );
  mux2_1 U12896 ( .ip1(i_i2c_rx_push_data[2]), .ip2(i_i2c_U_dff_rx_mem[58]), 
        .s(n11347), .op(n4898) );
  mux2_1 U12897 ( .ip1(i_i2c_rx_push_data[3]), .ip2(i_i2c_U_dff_rx_mem[3]), 
        .s(n11340), .op(n4897) );
  mux2_1 U12898 ( .ip1(i_i2c_rx_push_data[3]), .ip2(i_i2c_U_dff_rx_mem[11]), 
        .s(n11341), .op(n4896) );
  mux2_1 U12899 ( .ip1(i_i2c_rx_push_data[3]), .ip2(i_i2c_U_dff_rx_mem[19]), 
        .s(n11342), .op(n4895) );
  mux2_1 U12900 ( .ip1(i_i2c_rx_push_data[3]), .ip2(i_i2c_U_dff_rx_mem[27]), 
        .s(n11343), .op(n4894) );
  mux2_1 U12901 ( .ip1(i_i2c_U_dff_rx_mem[35]), .ip2(i_i2c_rx_push_data[3]), 
        .s(n11344), .op(n4893) );
  mux2_1 U12902 ( .ip1(i_i2c_rx_push_data[3]), .ip2(i_i2c_U_dff_rx_mem[43]), 
        .s(n11345), .op(n4892) );
  mux2_1 U12903 ( .ip1(i_i2c_U_dff_rx_mem[51]), .ip2(i_i2c_rx_push_data[3]), 
        .s(n11346), .op(n4891) );
  mux2_1 U12904 ( .ip1(i_i2c_rx_push_data[3]), .ip2(i_i2c_U_dff_rx_mem[59]), 
        .s(n11347), .op(n4890) );
  mux2_1 U12905 ( .ip1(i_i2c_rx_push_data[4]), .ip2(i_i2c_U_dff_rx_mem[4]), 
        .s(n11340), .op(n4889) );
  mux2_1 U12906 ( .ip1(i_i2c_rx_push_data[4]), .ip2(i_i2c_U_dff_rx_mem[12]), 
        .s(n11341), .op(n4888) );
  mux2_1 U12907 ( .ip1(i_i2c_rx_push_data[4]), .ip2(i_i2c_U_dff_rx_mem[20]), 
        .s(n11342), .op(n4887) );
  mux2_1 U12908 ( .ip1(i_i2c_rx_push_data[4]), .ip2(i_i2c_U_dff_rx_mem[28]), 
        .s(n11343), .op(n4886) );
  mux2_1 U12909 ( .ip1(i_i2c_U_dff_rx_mem[36]), .ip2(i_i2c_rx_push_data[4]), 
        .s(n11344), .op(n4885) );
  mux2_1 U12910 ( .ip1(i_i2c_rx_push_data[4]), .ip2(i_i2c_U_dff_rx_mem[44]), 
        .s(n11345), .op(n4884) );
  mux2_1 U12911 ( .ip1(i_i2c_U_dff_rx_mem[52]), .ip2(i_i2c_rx_push_data[4]), 
        .s(n11346), .op(n4883) );
  mux2_1 U12912 ( .ip1(i_i2c_rx_push_data[4]), .ip2(i_i2c_U_dff_rx_mem[60]), 
        .s(n11347), .op(n4882) );
  mux2_1 U12913 ( .ip1(i_i2c_rx_push_data[5]), .ip2(i_i2c_U_dff_rx_mem[5]), 
        .s(n11340), .op(n4881) );
  mux2_1 U12914 ( .ip1(i_i2c_rx_push_data[5]), .ip2(i_i2c_U_dff_rx_mem[13]), 
        .s(n11341), .op(n4880) );
  mux2_1 U12915 ( .ip1(i_i2c_rx_push_data[5]), .ip2(i_i2c_U_dff_rx_mem[21]), 
        .s(n11342), .op(n4879) );
  mux2_1 U12916 ( .ip1(i_i2c_rx_push_data[5]), .ip2(i_i2c_U_dff_rx_mem[29]), 
        .s(n11343), .op(n4878) );
  mux2_1 U12917 ( .ip1(i_i2c_U_dff_rx_mem[37]), .ip2(i_i2c_rx_push_data[5]), 
        .s(n11344), .op(n4877) );
  mux2_1 U12918 ( .ip1(i_i2c_rx_push_data[5]), .ip2(i_i2c_U_dff_rx_mem[45]), 
        .s(n11345), .op(n4876) );
  mux2_1 U12919 ( .ip1(i_i2c_U_dff_rx_mem[53]), .ip2(i_i2c_rx_push_data[5]), 
        .s(n11346), .op(n4875) );
  mux2_1 U12920 ( .ip1(i_i2c_rx_push_data[5]), .ip2(i_i2c_U_dff_rx_mem[61]), 
        .s(n11347), .op(n4874) );
  mux2_1 U12921 ( .ip1(i_i2c_rx_push_data[6]), .ip2(i_i2c_U_dff_rx_mem[6]), 
        .s(n11340), .op(n4873) );
  mux2_1 U12922 ( .ip1(i_i2c_rx_push_data[6]), .ip2(i_i2c_U_dff_rx_mem[14]), 
        .s(n11341), .op(n4872) );
  mux2_1 U12923 ( .ip1(i_i2c_rx_push_data[6]), .ip2(i_i2c_U_dff_rx_mem[22]), 
        .s(n11342), .op(n4871) );
  mux2_1 U12924 ( .ip1(i_i2c_rx_push_data[6]), .ip2(i_i2c_U_dff_rx_mem[30]), 
        .s(n11343), .op(n4870) );
  mux2_1 U12925 ( .ip1(i_i2c_U_dff_rx_mem[38]), .ip2(i_i2c_rx_push_data[6]), 
        .s(n11344), .op(n4869) );
  mux2_1 U12926 ( .ip1(i_i2c_rx_push_data[6]), .ip2(i_i2c_U_dff_rx_mem[46]), 
        .s(n11345), .op(n4868) );
  mux2_1 U12927 ( .ip1(i_i2c_U_dff_rx_mem[54]), .ip2(i_i2c_rx_push_data[6]), 
        .s(n11346), .op(n4867) );
  mux2_1 U12928 ( .ip1(i_i2c_rx_push_data[6]), .ip2(i_i2c_U_dff_rx_mem[62]), 
        .s(n11347), .op(n4866) );
  mux2_1 U12929 ( .ip1(i_i2c_rx_push_data[7]), .ip2(i_i2c_U_dff_rx_mem[7]), 
        .s(n11340), .op(n4865) );
  mux2_1 U12930 ( .ip1(i_i2c_rx_push_data[7]), .ip2(i_i2c_U_dff_rx_mem[15]), 
        .s(n11341), .op(n4864) );
  mux2_1 U12931 ( .ip1(i_i2c_rx_push_data[7]), .ip2(i_i2c_U_dff_rx_mem[23]), 
        .s(n11342), .op(n4863) );
  mux2_1 U12932 ( .ip1(i_i2c_rx_push_data[7]), .ip2(i_i2c_U_dff_rx_mem[31]), 
        .s(n11343), .op(n4862) );
  mux2_1 U12933 ( .ip1(i_i2c_U_dff_rx_mem[39]), .ip2(i_i2c_rx_push_data[7]), 
        .s(n11344), .op(n4861) );
  mux2_1 U12934 ( .ip1(i_i2c_rx_push_data[7]), .ip2(i_i2c_U_dff_rx_mem[47]), 
        .s(n11345), .op(n4860) );
  mux2_1 U12935 ( .ip1(i_i2c_U_dff_rx_mem[55]), .ip2(i_i2c_rx_push_data[7]), 
        .s(n11346), .op(n4859) );
  mux2_1 U12936 ( .ip1(i_i2c_rx_push_data[7]), .ip2(i_i2c_U_dff_rx_mem[63]), 
        .s(n11347), .op(n4858) );
  nor2_1 U12937 ( .ip1(i_ahb_U_mux_hsel_prev[4]), .ip2(n11348), .op(n11351) );
  nor2_1 U12938 ( .ip1(ex_i_ahb_AHB_Slave_PID_hready_resp), .ip2(n11348), .op(
        n11349) );
  nor2_1 U12939 ( .ip1(n11349), .ip2(ex_i_ahb_AHB_Slave_PID_hsel), .op(n11350)
         );
  nor2_1 U12940 ( .ip1(n11351), .ip2(n11350), .op(n4852) );
  mux2_1 U12941 ( .ip1(i_ahb_U_mux_hsel_prev[1]), .ip2(
        ex_i_ahb_AHB_Slave_RAM_hsel), .s(ex_i_ahb_AHB_MASTER_CORTEXM0_hready), 
        .op(n4849) );
  mux2_1 U12942 ( .ip1(ex_i_ahb_AHB_Slave_PID_hmastlock), .ip2(
        ex_i_ahb_AHB_MASTER_CORTEXM0_hlock), .s(ex_i_ahb_AHB_Slave_PID_hready), 
        .op(n4848) );
  inv_1 U12943 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[0]), .op(
        n11353) );
  nor2_1 U12944 ( .ip1(n11353), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[0]), .op(n11352) );
  not_ab_or_c_or_d U12945 ( .ip1(n11353), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[0]), .ip3(
        i_i2c_ic_tx_abrt_source[0]), .ip4(n11352), .op(n11354) );
  nor2_1 U12946 ( .ip1(n11400), .ip2(n11354), .op(n4700) );
  inv_1 U12947 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[1]), .op(
        n11356) );
  nor2_1 U12948 ( .ip1(n11356), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[1]), .op(n11355) );
  not_ab_or_c_or_d U12949 ( .ip1(n11356), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[1]), .ip3(
        i_i2c_ic_tx_abrt_source[1]), .ip4(n11355), .op(n11357) );
  nor2_1 U12950 ( .ip1(n11400), .ip2(n11357), .op(n4699) );
  inv_1 U12951 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[2]), .op(
        n11359) );
  nor2_1 U12952 ( .ip1(n11359), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[2]), .op(n11358) );
  not_ab_or_c_or_d U12953 ( .ip1(n11359), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[2]), .ip3(
        i_i2c_ic_tx_abrt_source[2]), .ip4(n11358), .op(n11360) );
  nor2_1 U12954 ( .ip1(n11400), .ip2(n11360), .op(n4698) );
  inv_1 U12955 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[3]), .op(
        n11362) );
  nor2_1 U12956 ( .ip1(n11362), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[3]), .op(n11361) );
  not_ab_or_c_or_d U12957 ( .ip1(n11362), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[3]), .ip3(
        i_i2c_ic_tx_abrt_source[3]), .ip4(n11361), .op(n11363) );
  nor2_1 U12958 ( .ip1(n11400), .ip2(n11363), .op(n4697) );
  inv_1 U12959 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[4]), .op(
        n11365) );
  nor2_1 U12960 ( .ip1(n11365), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[4]), .op(n11364) );
  not_ab_or_c_or_d U12961 ( .ip1(n11365), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[4]), .ip3(
        i_i2c_ic_tx_abrt_source[4]), .ip4(n11364), .op(n11366) );
  nor2_1 U12962 ( .ip1(n11400), .ip2(n11366), .op(n4696) );
  inv_1 U12963 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[5]), .op(
        n11368) );
  nor2_1 U12964 ( .ip1(n11368), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[5]), .op(n11367) );
  not_ab_or_c_or_d U12965 ( .ip1(n11368), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[5]), .ip3(
        i_i2c_ic_tx_abrt_source[5]), .ip4(n11367), .op(n11369) );
  nor2_1 U12966 ( .ip1(n11400), .ip2(n11369), .op(n4695) );
  inv_1 U12967 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[6]), .op(
        n11371) );
  nor2_1 U12968 ( .ip1(n11371), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[6]), .op(n11370) );
  not_ab_or_c_or_d U12969 ( .ip1(n11371), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[6]), .ip3(
        i_i2c_ic_tx_abrt_source[6]), .ip4(n11370), .op(n11372) );
  nor2_1 U12970 ( .ip1(n11400), .ip2(n11372), .op(n4694) );
  inv_1 U12971 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[7]), .op(
        n11374) );
  nor2_1 U12972 ( .ip1(n11374), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[7]), .op(n11373) );
  not_ab_or_c_or_d U12973 ( .ip1(n11374), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[7]), .ip3(
        i_i2c_ic_tx_abrt_source[7]), .ip4(n11373), .op(n11375) );
  nor2_1 U12974 ( .ip1(n11400), .ip2(n11375), .op(n4693) );
  inv_1 U12975 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[8]), .op(
        n11377) );
  nor2_1 U12976 ( .ip1(n11377), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[8]), .op(n11376) );
  not_ab_or_c_or_d U12977 ( .ip1(n11377), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[8]), .ip3(
        i_i2c_ic_tx_abrt_source[8]), .ip4(n11376), .op(n11378) );
  nor2_1 U12978 ( .ip1(n11400), .ip2(n11378), .op(n4692) );
  inv_1 U12979 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[9]), .op(
        n11380) );
  nor2_1 U12980 ( .ip1(n11380), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[9]), .op(n11379) );
  not_ab_or_c_or_d U12981 ( .ip1(n11380), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[9]), .ip3(
        i_i2c_ic_tx_abrt_source[9]), .ip4(n11379), .op(n11381) );
  nor2_1 U12982 ( .ip1(n11400), .ip2(n11381), .op(n4691) );
  inv_1 U12983 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[10]), .op(
        n11383) );
  nor2_1 U12984 ( .ip1(n11383), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[10]), .op(n11382) );
  not_ab_or_c_or_d U12985 ( .ip1(n11383), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[10]), .ip3(
        i_i2c_ic_tx_abrt_source[10]), .ip4(n11382), .op(n11384) );
  nor2_1 U12986 ( .ip1(n11400), .ip2(n11384), .op(n4690) );
  inv_1 U12987 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[11]), .op(
        n11386) );
  nor2_1 U12988 ( .ip1(n11386), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[11]), .op(n11385) );
  not_ab_or_c_or_d U12989 ( .ip1(n11386), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[11]), .ip3(
        i_i2c_ic_tx_abrt_source[11]), .ip4(n11385), .op(n11387) );
  nor2_1 U12990 ( .ip1(n11400), .ip2(n11387), .op(n4689) );
  inv_1 U12991 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[12]), .op(
        n11389) );
  nor2_1 U12992 ( .ip1(n11389), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[12]), .op(n11388) );
  not_ab_or_c_or_d U12993 ( .ip1(n11389), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[12]), .ip3(
        i_i2c_ic_tx_abrt_source[12]), .ip4(n11388), .op(n11390) );
  nor2_1 U12994 ( .ip1(n11400), .ip2(n11390), .op(n4688) );
  inv_1 U12995 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[13]), .op(
        n11392) );
  nor2_1 U12996 ( .ip1(n11392), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[13]), .op(n11391) );
  not_ab_or_c_or_d U12997 ( .ip1(n11392), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[13]), .ip3(
        i_i2c_ic_tx_abrt_source[13]), .ip4(n11391), .op(n11393) );
  nor2_1 U12998 ( .ip1(n11400), .ip2(n11393), .op(n4687) );
  inv_1 U12999 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[14]), .op(
        n11395) );
  nor2_1 U13000 ( .ip1(n11395), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[14]), .op(n11394) );
  not_ab_or_c_or_d U13001 ( .ip1(n11395), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[14]), .ip3(
        i_i2c_ic_tx_abrt_source[14]), .ip4(n11394), .op(n11396) );
  nor2_1 U13002 ( .ip1(n11400), .ip2(n11396), .op(n4686) );
  inv_1 U13003 ( .ip(i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync[15]), .op(
        n11398) );
  nor2_1 U13004 ( .ip1(n11398), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[15]), .op(n11397) );
  not_ab_or_c_or_d U13005 ( .ip1(n11398), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_tx_abrt_source_sync_q[15]), .ip3(
        i_i2c_ic_tx_abrt_source[15]), .ip4(n11397), .op(n11399) );
  nor2_1 U13006 ( .ip1(n11400), .ip2(n11399), .op(n4685) );
  mux2_1 U13007 ( .ip1(i_i2c_prdata[30]), .ip2(i_i2c_iprdata[30]), .s(n11839), 
        .op(n4684) );
  mux2_1 U13008 ( .ip1(i_i2c_prdata[29]), .ip2(i_i2c_iprdata[29]), .s(n11401), 
        .op(n4683) );
  mux2_1 U13009 ( .ip1(i_i2c_prdata[28]), .ip2(i_i2c_iprdata[29]), .s(n11839), 
        .op(n4682) );
  mux2_1 U13010 ( .ip1(i_i2c_prdata[26]), .ip2(i_i2c_iprdata[26]), .s(n11839), 
        .op(n4680) );
  mux2_1 U13011 ( .ip1(i_i2c_prdata[25]), .ip2(i_i2c_iprdata[25]), .s(n11839), 
        .op(n4679) );
  mux2_1 U13012 ( .ip1(i_i2c_prdata[24]), .ip2(i_i2c_iprdata[24]), .s(n11401), 
        .op(n4678) );
  mux2_1 U13013 ( .ip1(i_i2c_prdata[23]), .ip2(i_i2c_iprdata[23]), .s(n11401), 
        .op(n4677) );
  mux2_1 U13014 ( .ip1(i_i2c_prdata[22]), .ip2(i_i2c_iprdata[22]), .s(n11401), 
        .op(n4676) );
  mux2_1 U13015 ( .ip1(i_i2c_prdata[21]), .ip2(i_i2c_iprdata[21]), .s(n11401), 
        .op(n4675) );
  mux2_1 U13016 ( .ip1(i_i2c_prdata[20]), .ip2(i_i2c_iprdata[20]), .s(n11401), 
        .op(n4674) );
  mux2_1 U13017 ( .ip1(i_i2c_prdata[19]), .ip2(i_i2c_iprdata[19]), .s(n11401), 
        .op(n4673) );
  mux2_1 U13018 ( .ip1(i_i2c_prdata[18]), .ip2(i_i2c_iprdata[18]), .s(n11401), 
        .op(n4672) );
  mux2_1 U13019 ( .ip1(i_i2c_prdata[17]), .ip2(i_i2c_iprdata[17]), .s(n11401), 
        .op(n4671) );
  mux2_1 U13020 ( .ip1(i_i2c_prdata[16]), .ip2(i_i2c_iprdata[16]), .s(n11401), 
        .op(n4670) );
  mux2_1 U13021 ( .ip1(i_i2c_prdata[15]), .ip2(i_i2c_iprdata[15]), .s(n11401), 
        .op(n4669) );
  mux2_1 U13022 ( .ip1(i_i2c_prdata[14]), .ip2(i_i2c_iprdata[14]), .s(n11401), 
        .op(n4668) );
  mux2_1 U13023 ( .ip1(i_i2c_prdata[13]), .ip2(i_i2c_iprdata[13]), .s(n11401), 
        .op(n4667) );
  mux2_1 U13024 ( .ip1(i_i2c_prdata[12]), .ip2(i_i2c_iprdata[12]), .s(n11839), 
        .op(n4666) );
  mux2_1 U13025 ( .ip1(i_i2c_prdata[11]), .ip2(i_i2c_iprdata[11]), .s(n11839), 
        .op(n4665) );
  mux2_1 U13026 ( .ip1(i_i2c_prdata[10]), .ip2(i_i2c_iprdata[10]), .s(n11839), 
        .op(n4664) );
  mux2_1 U13027 ( .ip1(i_i2c_prdata[9]), .ip2(i_i2c_iprdata[9]), .s(n11839), 
        .op(n4663) );
  mux2_1 U13028 ( .ip1(i_i2c_prdata[8]), .ip2(i_i2c_iprdata[8]), .s(n11839), 
        .op(n4662) );
  mux2_1 U13029 ( .ip1(i_i2c_prdata[7]), .ip2(i_i2c_iprdata[7]), .s(n11401), 
        .op(n4661) );
  mux2_1 U13030 ( .ip1(i_i2c_prdata[6]), .ip2(i_i2c_iprdata[6]), .s(n11401), 
        .op(n4660) );
  mux2_1 U13031 ( .ip1(i_i2c_prdata[5]), .ip2(i_i2c_iprdata[5]), .s(n11401), 
        .op(n4659) );
  mux2_1 U13032 ( .ip1(i_i2c_prdata[4]), .ip2(i_i2c_iprdata[4]), .s(n11401), 
        .op(n4658) );
  mux2_1 U13033 ( .ip1(i_i2c_prdata[3]), .ip2(i_i2c_iprdata[3]), .s(n11401), 
        .op(n4657) );
  mux2_1 U13034 ( .ip1(i_i2c_prdata[2]), .ip2(i_i2c_iprdata[2]), .s(n11401), 
        .op(n4656) );
  mux2_1 U13035 ( .ip1(i_i2c_prdata[1]), .ip2(i_i2c_iprdata[1]), .s(n11401), 
        .op(n4655) );
  mux2_1 U13036 ( .ip1(i_i2c_prdata[0]), .ip2(i_i2c_iprdata[0]), .s(n11401), 
        .op(n4654) );
  nor2_1 U13037 ( .ip1(i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync_q), .op(n11403) );
  inv_1 U13038 ( .ip(i_i2c_ic_ack_general_call), .op(n11402) );
  not_ab_or_c_or_d U13039 ( .ip1(
        i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_rx_gen_call_flg_sync_q), .ip3(n11403), .ip4(
        n11402), .op(n11405) );
  or2_1 U13040 ( .ip1(i_i2c_ic_raw_intr_stat[11]), .ip2(n11405), .op(n11408)
         );
  or2_1 U13041 ( .ip1(i_i2c_ic_clr_intr_en), .ip2(i_i2c_ic_clr_gen_call_en), 
        .op(n11404) );
  nand2_1 U13042 ( .ip1(n11839), .ip2(n11404), .op(n11406) );
  or2_1 U13043 ( .ip1(n11406), .ip2(n11405), .op(n11407) );
  nand2_1 U13044 ( .ip1(n11408), .ip2(n11407), .op(n11409) );
  nor2_1 U13045 ( .ip1(n11409), .ip2(n11449), .op(n4653) );
  xor2_1 U13046 ( .ip1(i_i2c_U_DW_apb_i2c_intctl_p_det_flg_sync), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_p_det_flg_sync_q), .op(n11411) );
  or2_1 U13047 ( .ip1(i_i2c_ic_raw_intr_stat[9]), .ip2(n11411), .op(n11414) );
  or2_1 U13048 ( .ip1(i_i2c_ic_clr_intr_en), .ip2(i_i2c_ic_clr_stop_det_en), 
        .op(n11410) );
  nand2_1 U13049 ( .ip1(n11839), .ip2(n11410), .op(n11412) );
  or2_1 U13050 ( .ip1(n11412), .ip2(n11411), .op(n11413) );
  nand2_1 U13051 ( .ip1(n11414), .ip2(n11413), .op(n11415) );
  nor2_1 U13052 ( .ip1(n11415), .ip2(n11449), .op(n4652) );
  xor2_1 U13053 ( .ip1(i_i2c_U_DW_apb_i2c_intctl_s_det_flg_sync), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_s_det_flg_sync_q), .op(n11417) );
  or2_1 U13054 ( .ip1(i_i2c_ic_raw_intr_stat[10]), .ip2(n11417), .op(n11420)
         );
  or2_1 U13055 ( .ip1(i_i2c_ic_clr_intr_en), .ip2(i_i2c_ic_clr_start_det_en), 
        .op(n11416) );
  nand2_1 U13056 ( .ip1(n11839), .ip2(n11416), .op(n11418) );
  or2_1 U13057 ( .ip1(n11418), .ip2(n11417), .op(n11419) );
  nand2_1 U13058 ( .ip1(n11420), .ip2(n11419), .op(n11421) );
  nor2_1 U13059 ( .ip1(n11421), .ip2(n11449), .op(n4651) );
  or2_1 U13060 ( .ip1(i_i2c_ic_raw_intr_stat[8]), .ip2(i_i2c_activity), .op(
        n11425) );
  or2_1 U13061 ( .ip1(i_i2c_ic_clr_intr_en), .ip2(i_i2c_ic_clr_activity_en), 
        .op(n11422) );
  nand2_1 U13062 ( .ip1(n11839), .ip2(n11422), .op(n11423) );
  or2_1 U13063 ( .ip1(n11423), .ip2(i_i2c_activity), .op(n11424) );
  nand2_1 U13064 ( .ip1(n11425), .ip2(n11424), .op(n11426) );
  nor2_1 U13065 ( .ip1(n11426), .ip2(n11449), .op(n4650) );
  xor2_1 U13066 ( .ip1(i_i2c_U_DW_apb_i2c_intctl_rx_done_flg_sync), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_rx_done_flg_sync_q), .op(n11428) );
  or2_1 U13067 ( .ip1(i_i2c_ic_raw_intr_stat[7]), .ip2(n11428), .op(n11431) );
  or2_1 U13068 ( .ip1(i_i2c_ic_clr_intr_en), .ip2(i_i2c_ic_clr_rx_done_en), 
        .op(n11427) );
  nand2_1 U13069 ( .ip1(n11839), .ip2(n11427), .op(n11429) );
  or2_1 U13070 ( .ip1(n11429), .ip2(n11428), .op(n11430) );
  nand2_1 U13071 ( .ip1(n11431), .ip2(n11430), .op(n11432) );
  nor2_1 U13072 ( .ip1(n11432), .ip2(n11449), .op(n4649) );
  or2_1 U13073 ( .ip1(i_i2c_ic_raw_intr_stat[6]), .ip2(i_i2c_tx_abrt_flg_edg), 
        .op(n11435) );
  or2_1 U13074 ( .ip1(n11433), .ip2(i_i2c_tx_abrt_flg_edg), .op(n11434) );
  nand2_1 U13075 ( .ip1(n11435), .ip2(n11434), .op(n11436) );
  nor2_1 U13076 ( .ip1(n11436), .ip2(n11449), .op(n4648) );
  xor2_1 U13077 ( .ip1(i_i2c_U_DW_apb_i2c_intctl_ic_rd_req_flg_sync), .ip2(
        i_i2c_U_DW_apb_i2c_intctl_ic_rd_req_flg_sync_q), .op(n11438) );
  or2_1 U13078 ( .ip1(i_i2c_ic_raw_intr_stat[5]), .ip2(n11438), .op(n11441) );
  or2_1 U13079 ( .ip1(i_i2c_ic_clr_intr_en), .ip2(i_i2c_ic_clr_rd_req_en), 
        .op(n11437) );
  nand2_1 U13080 ( .ip1(n11839), .ip2(n11437), .op(n11439) );
  or2_1 U13081 ( .ip1(n11439), .ip2(n11438), .op(n11440) );
  nand2_1 U13082 ( .ip1(n11441), .ip2(n11440), .op(n11442) );
  nor2_1 U13083 ( .ip1(n11442), .ip2(n11449), .op(n4647) );
  nand2_1 U13084 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_tx_error_ir), .ip2(
        i_i2c_U_DW_apb_i2c_fifo_tx_push_dly), .op(n11443) );
  nor2_1 U13085 ( .ip1(i_i2c_U_DW_apb_i2c_fifo_tx_pop_sync_dly), .ip2(n11443), 
        .op(n11445) );
  or2_1 U13086 ( .ip1(i_i2c_ic_raw_intr_stat[3]), .ip2(n11445), .op(n11448) );
  or2_1 U13087 ( .ip1(i_i2c_ic_clr_intr_en), .ip2(i_i2c_ic_clr_tx_over_en), 
        .op(n11444) );
  nand2_1 U13088 ( .ip1(n11839), .ip2(n11444), .op(n11446) );
  or2_1 U13089 ( .ip1(n11446), .ip2(n11445), .op(n11447) );
  nand2_1 U13090 ( .ip1(n11448), .ip2(n11447), .op(n11450) );
  nor2_1 U13091 ( .ip1(n11450), .ip2(n11449), .op(n4644) );
  mux2_1 U13092 ( .ip1(i_apb_pwdata_int[2]), .ip2(i_ssi_txftlr[2]), .s(n11451), 
        .op(n4632) );
  mux2_1 U13093 ( .ip1(i_ssi_U_dff_rx_mem[6]), .ip2(i_ssi_rx_push_data[6]), 
        .s(n10777), .op(n4322) );
  mux2_1 U13094 ( .ip1(i_ssi_rx_push_data[6]), .ip2(i_ssi_U_dff_rx_mem[22]), 
        .s(n11452), .op(n4321) );
  mux2_1 U13095 ( .ip1(i_ssi_U_dff_rx_mem[38]), .ip2(i_ssi_rx_push_data[6]), 
        .s(n5610), .op(n4320) );
  mux2_1 U13096 ( .ip1(i_ssi_rx_push_data[6]), .ip2(i_ssi_U_dff_rx_mem[54]), 
        .s(n11453), .op(n4319) );
  mux2_1 U13097 ( .ip1(i_ssi_U_dff_rx_mem[70]), .ip2(i_ssi_rx_push_data[6]), 
        .s(n10721), .op(n4318) );
  mux2_1 U13098 ( .ip1(i_ssi_rx_push_data[6]), .ip2(i_ssi_U_dff_rx_mem[86]), 
        .s(n11454), .op(n4317) );
  mux2_1 U13099 ( .ip1(i_ssi_U_dff_rx_mem[102]), .ip2(i_ssi_rx_push_data[6]), 
        .s(n5611), .op(n4316) );
  mux2_1 U13100 ( .ip1(i_ssi_rx_push_data[6]), .ip2(i_ssi_U_dff_rx_mem[118]), 
        .s(n11455), .op(n4315) );
  mux2_1 U13101 ( .ip1(i_ssi_U_dff_rx_mem[8]), .ip2(i_ssi_rx_push_data[8]), 
        .s(n10777), .op(n4306) );
  mux2_1 U13102 ( .ip1(i_ssi_rx_push_data[8]), .ip2(i_ssi_U_dff_rx_mem[24]), 
        .s(n11452), .op(n4305) );
  mux2_1 U13103 ( .ip1(i_ssi_U_dff_rx_mem[40]), .ip2(i_ssi_rx_push_data[8]), 
        .s(n5610), .op(n4304) );
  mux2_1 U13104 ( .ip1(i_ssi_rx_push_data[8]), .ip2(i_ssi_U_dff_rx_mem[56]), 
        .s(n11453), .op(n4303) );
  mux2_1 U13105 ( .ip1(i_ssi_U_dff_rx_mem[72]), .ip2(i_ssi_rx_push_data[8]), 
        .s(n10721), .op(n4302) );
  mux2_1 U13106 ( .ip1(i_ssi_rx_push_data[8]), .ip2(i_ssi_U_dff_rx_mem[88]), 
        .s(n11454), .op(n4301) );
  mux2_1 U13107 ( .ip1(i_ssi_U_dff_rx_mem[104]), .ip2(i_ssi_rx_push_data[8]), 
        .s(n5611), .op(n4300) );
  mux2_1 U13108 ( .ip1(i_ssi_rx_push_data[8]), .ip2(i_ssi_U_dff_rx_mem[120]), 
        .s(n11455), .op(n4299) );
  mux2_1 U13109 ( .ip1(i_ssi_U_dff_rx_mem[9]), .ip2(i_ssi_rx_push_data[9]), 
        .s(n10777), .op(n4298) );
  mux2_1 U13110 ( .ip1(i_ssi_rx_push_data[9]), .ip2(i_ssi_U_dff_rx_mem[25]), 
        .s(n11452), .op(n4297) );
  mux2_1 U13111 ( .ip1(i_ssi_U_dff_rx_mem[41]), .ip2(i_ssi_rx_push_data[9]), 
        .s(n5610), .op(n4296) );
  mux2_1 U13112 ( .ip1(i_ssi_rx_push_data[9]), .ip2(i_ssi_U_dff_rx_mem[57]), 
        .s(n11453), .op(n4295) );
  mux2_1 U13113 ( .ip1(i_ssi_U_dff_rx_mem[73]), .ip2(i_ssi_rx_push_data[9]), 
        .s(n10721), .op(n4294) );
  mux2_1 U13114 ( .ip1(i_ssi_rx_push_data[9]), .ip2(i_ssi_U_dff_rx_mem[89]), 
        .s(n11454), .op(n4293) );
  mux2_1 U13115 ( .ip1(i_ssi_U_dff_rx_mem[105]), .ip2(i_ssi_rx_push_data[9]), 
        .s(n5611), .op(n4292) );
  mux2_1 U13116 ( .ip1(i_ssi_rx_push_data[9]), .ip2(i_ssi_U_dff_rx_mem[121]), 
        .s(n11455), .op(n4291) );
  mux2_1 U13117 ( .ip1(i_ssi_U_dff_rx_mem[10]), .ip2(i_ssi_rx_push_data[10]), 
        .s(n10777), .op(n4290) );
  mux2_1 U13118 ( .ip1(i_ssi_rx_push_data[10]), .ip2(i_ssi_U_dff_rx_mem[26]), 
        .s(n11452), .op(n4289) );
  mux2_1 U13119 ( .ip1(i_ssi_U_dff_rx_mem[42]), .ip2(i_ssi_rx_push_data[10]), 
        .s(n5610), .op(n4288) );
  mux2_1 U13120 ( .ip1(i_ssi_rx_push_data[10]), .ip2(i_ssi_U_dff_rx_mem[58]), 
        .s(n11453), .op(n4287) );
  mux2_1 U13121 ( .ip1(i_ssi_U_dff_rx_mem[74]), .ip2(i_ssi_rx_push_data[10]), 
        .s(n10721), .op(n4286) );
  mux2_1 U13122 ( .ip1(i_ssi_rx_push_data[10]), .ip2(i_ssi_U_dff_rx_mem[90]), 
        .s(n11454), .op(n4285) );
  mux2_1 U13123 ( .ip1(i_ssi_U_dff_rx_mem[106]), .ip2(i_ssi_rx_push_data[10]), 
        .s(n5611), .op(n4284) );
  mux2_1 U13124 ( .ip1(i_ssi_rx_push_data[10]), .ip2(i_ssi_U_dff_rx_mem[122]), 
        .s(n11455), .op(n4283) );
  mux2_1 U13125 ( .ip1(i_ssi_U_dff_rx_mem[11]), .ip2(i_ssi_rx_push_data[11]), 
        .s(n10777), .op(n4282) );
  mux2_1 U13126 ( .ip1(i_ssi_rx_push_data[11]), .ip2(i_ssi_U_dff_rx_mem[27]), 
        .s(n11452), .op(n4281) );
  mux2_1 U13127 ( .ip1(i_ssi_U_dff_rx_mem[43]), .ip2(i_ssi_rx_push_data[11]), 
        .s(n5610), .op(n4280) );
  mux2_1 U13128 ( .ip1(i_ssi_rx_push_data[11]), .ip2(i_ssi_U_dff_rx_mem[59]), 
        .s(n11453), .op(n4279) );
  mux2_1 U13129 ( .ip1(i_ssi_U_dff_rx_mem[75]), .ip2(i_ssi_rx_push_data[11]), 
        .s(n10721), .op(n4278) );
  mux2_1 U13130 ( .ip1(i_ssi_rx_push_data[11]), .ip2(i_ssi_U_dff_rx_mem[91]), 
        .s(n11454), .op(n4277) );
  mux2_1 U13131 ( .ip1(i_ssi_U_dff_rx_mem[107]), .ip2(i_ssi_rx_push_data[11]), 
        .s(n5611), .op(n4276) );
  mux2_1 U13132 ( .ip1(i_ssi_rx_push_data[11]), .ip2(i_ssi_U_dff_rx_mem[123]), 
        .s(n11455), .op(n4275) );
  mux2_1 U13133 ( .ip1(i_ssi_U_dff_rx_mem[12]), .ip2(i_ssi_rx_push_data[12]), 
        .s(n10777), .op(n4274) );
  mux2_1 U13134 ( .ip1(i_ssi_rx_push_data[12]), .ip2(i_ssi_U_dff_rx_mem[28]), 
        .s(n11452), .op(n4273) );
  mux2_1 U13135 ( .ip1(i_ssi_U_dff_rx_mem[44]), .ip2(i_ssi_rx_push_data[12]), 
        .s(n5610), .op(n4272) );
  mux2_1 U13136 ( .ip1(i_ssi_rx_push_data[12]), .ip2(i_ssi_U_dff_rx_mem[60]), 
        .s(n11453), .op(n4271) );
  mux2_1 U13137 ( .ip1(i_ssi_U_dff_rx_mem[76]), .ip2(i_ssi_rx_push_data[12]), 
        .s(n10721), .op(n4270) );
  mux2_1 U13138 ( .ip1(i_ssi_rx_push_data[12]), .ip2(i_ssi_U_dff_rx_mem[92]), 
        .s(n11454), .op(n4269) );
  mux2_1 U13139 ( .ip1(i_ssi_U_dff_rx_mem[108]), .ip2(i_ssi_rx_push_data[12]), 
        .s(n5611), .op(n4268) );
  mux2_1 U13140 ( .ip1(i_ssi_rx_push_data[12]), .ip2(i_ssi_U_dff_rx_mem[124]), 
        .s(n11455), .op(n4267) );
  mux2_1 U13141 ( .ip1(i_ssi_U_dff_rx_mem[13]), .ip2(i_ssi_rx_push_data[13]), 
        .s(n10777), .op(n4266) );
  mux2_1 U13142 ( .ip1(i_ssi_rx_push_data[13]), .ip2(i_ssi_U_dff_rx_mem[29]), 
        .s(n11452), .op(n4265) );
  mux2_1 U13143 ( .ip1(i_ssi_U_dff_rx_mem[45]), .ip2(i_ssi_rx_push_data[13]), 
        .s(n5610), .op(n4264) );
  mux2_1 U13144 ( .ip1(i_ssi_rx_push_data[13]), .ip2(i_ssi_U_dff_rx_mem[61]), 
        .s(n11453), .op(n4263) );
  mux2_1 U13145 ( .ip1(i_ssi_U_dff_rx_mem[77]), .ip2(i_ssi_rx_push_data[13]), 
        .s(n10721), .op(n4262) );
  mux2_1 U13146 ( .ip1(i_ssi_rx_push_data[13]), .ip2(i_ssi_U_dff_rx_mem[93]), 
        .s(n11454), .op(n4261) );
  mux2_1 U13147 ( .ip1(i_ssi_U_dff_rx_mem[109]), .ip2(i_ssi_rx_push_data[13]), 
        .s(n5611), .op(n4260) );
  mux2_1 U13148 ( .ip1(i_ssi_rx_push_data[13]), .ip2(i_ssi_U_dff_rx_mem[125]), 
        .s(n11455), .op(n4259) );
  inv_1 U13149 ( .ip(n11456), .op(n11461) );
  inv_1 U13150 ( .ip(n11457), .op(n11458) );
  nor3_1 U13151 ( .ip1(i_ssi_reg_addr[0]), .ip2(n11458), .ip3(
        i_ssi_ssi_rxu_intr_n), .op(n11459) );
  not_ab_or_c_or_d U13152 ( .ip1(n11461), .ip2(n11460), .ip3(n11661), .ip4(
        n11459), .op(n11507) );
  nand3_1 U13153 ( .ip1(i_ssi_ssi_rxu_intr_n), .ip2(i_ssi_ssi_txo_intr_n), 
        .ip3(i_ssi_ssi_rxo_intr_n), .op(n11466) );
  nor2_1 U13154 ( .ip1(n11462), .ip2(i_ssi_ssi_mst_intr_n), .op(n11465) );
  nor3_1 U13155 ( .ip1(n11463), .ip2(n11484), .ip3(i_ssi_ssi_rxo_intr_n), .op(
        n11464) );
  not_ab_or_c_or_d U13156 ( .ip1(n11467), .ip2(n11466), .ip3(n11465), .ip4(
        n11464), .op(n11506) );
  nor2_1 U13157 ( .ip1(i_ssi_ssi_txe_intr_n), .ip2(n11634), .op(n11489) );
  and3_1 U13158 ( .ip1(n11469), .ip2(i_ssi_ser_0_), .ip3(n11468), .op(n11473)
         );
  nor2_1 U13159 ( .ip1(n11471), .ip2(n11470), .op(n11472) );
  not_ab_or_c_or_d U13160 ( .ip1(i_ssi_U_regfile_ctrlr1_int[0]), .ip2(n11636), 
        .ip3(n11473), .ip4(n11472), .op(n11474) );
  inv_1 U13161 ( .ip(n11474), .op(n11477) );
  inv_1 U13162 ( .ip(n11475), .op(n11476) );
  mux3_2 U13163 ( .ip1(n11477), .ip2(i_ssi_mwcr[0]), .ip3(n10802), .s0(n11548), 
        .s1(n11476), .op(n11478) );
  mux2_1 U13164 ( .ip1(i_ssi_txftlr[0]), .ip2(n11478), .s(n11527), .op(n11479)
         );
  mux2_1 U13165 ( .ip1(i_ssi_rxftlr[0]), .ip2(n11479), .s(n11529), .op(n11480)
         );
  inv_1 U13166 ( .ip(n11647), .op(n11545) );
  mux2_1 U13167 ( .ip1(i_ssi_fsm_busy), .ip2(n11480), .s(n11545), .op(n11483)
         );
  nand2_1 U13168 ( .ip1(n11482), .ip2(n11481), .op(n11522) );
  mux2_1 U13169 ( .ip1(i_ssi_U_regfile_txflr[0]), .ip2(n11483), .s(n11522), 
        .op(n11488) );
  or2_1 U13170 ( .ip1(n11485), .ip2(n11484), .op(n11537) );
  nor2_1 U13171 ( .ip1(n11486), .ip2(n11537), .op(n11487) );
  nor3_1 U13172 ( .ip1(n11489), .ip2(n11488), .ip3(n11487), .op(n11504) );
  nand2_1 U13173 ( .ip1(n11617), .ip2(i_ssi_U_dff_rx_mem[16]), .op(n11499) );
  inv_1 U13174 ( .ip(i_ssi_U_dff_rx_mem[32]), .op(n11490) );
  nor2_1 U13175 ( .ip1(n11616), .ip2(n11490), .op(n11496) );
  nand2_1 U13176 ( .ip1(n11620), .ip2(i_ssi_U_dff_rx_mem[0]), .op(n11494) );
  nand2_1 U13177 ( .ip1(n11628), .ip2(i_ssi_U_dff_rx_mem[80]), .op(n11493) );
  nand2_1 U13178 ( .ip1(n11627), .ip2(i_ssi_U_dff_rx_mem[112]), .op(n11492) );
  nand2_1 U13179 ( .ip1(n11619), .ip2(i_ssi_U_dff_rx_mem[96]), .op(n11491) );
  nand4_1 U13180 ( .ip1(n11494), .ip2(n11493), .ip3(n11492), .ip4(n11491), 
        .op(n11495) );
  not_ab_or_c_or_d U13181 ( .ip1(i_ssi_U_dff_rx_mem[48]), .ip2(n11614), .ip3(
        n11496), .ip4(n11495), .op(n11498) );
  nand2_1 U13182 ( .ip1(n11618), .ip2(i_ssi_U_dff_rx_mem[64]), .op(n11497) );
  nand3_1 U13183 ( .ip1(n11499), .ip2(n11498), .ip3(n11497), .op(n11500) );
  nand2_1 U13184 ( .ip1(n11632), .ip2(n11500), .op(n11503) );
  nand2_1 U13185 ( .ip1(n11641), .ip2(i_ssi_risr[0]), .op(n11502) );
  nand2_1 U13186 ( .ip1(n11640), .ip2(i_ssi_imr[0]), .op(n11501) );
  and4_1 U13187 ( .ip1(n11504), .ip2(n11503), .ip3(n11502), .ip4(n11501), .op(
        n11505) );
  nand3_1 U13188 ( .ip1(n11507), .ip2(n11506), .ip3(n11505), .op(n11508) );
  nand2_1 U13189 ( .ip1(n11651), .ip2(n11508), .op(n11510) );
  nand2_1 U13190 ( .ip1(i_ssi_prdata[0]), .ip2(n11663), .op(n11509) );
  nand2_1 U13191 ( .ip1(n11510), .ip2(n11509), .op(n4237) );
  nand2_1 U13192 ( .ip1(n11618), .ip2(i_ssi_U_dff_rx_mem[65]), .op(n11520) );
  inv_1 U13193 ( .ip(i_ssi_U_dff_rx_mem[33]), .op(n11511) );
  nor2_1 U13194 ( .ip1(n11616), .ip2(n11511), .op(n11517) );
  nand2_1 U13195 ( .ip1(n11620), .ip2(i_ssi_U_dff_rx_mem[1]), .op(n11515) );
  nand2_1 U13196 ( .ip1(n11627), .ip2(i_ssi_U_dff_rx_mem[113]), .op(n11514) );
  nand2_1 U13197 ( .ip1(n11628), .ip2(i_ssi_U_dff_rx_mem[81]), .op(n11513) );
  nand2_1 U13198 ( .ip1(n11617), .ip2(i_ssi_U_dff_rx_mem[17]), .op(n11512) );
  nand4_1 U13199 ( .ip1(n11515), .ip2(n11514), .ip3(n11513), .ip4(n11512), 
        .op(n11516) );
  not_ab_or_c_or_d U13200 ( .ip1(n11614), .ip2(i_ssi_U_dff_rx_mem[49]), .ip3(
        n11517), .ip4(n11516), .op(n11519) );
  nand2_1 U13201 ( .ip1(n11619), .ip2(i_ssi_U_dff_rx_mem[97]), .op(n11518) );
  nand3_1 U13202 ( .ip1(n11520), .ip2(n11519), .ip3(n11518), .op(n11521) );
  nand2_1 U13203 ( .ip1(n11632), .ip2(n11521), .op(n11542) );
  nor2_1 U13204 ( .ip1(i_ssi_ssi_txo_intr_n), .ip2(n11634), .op(n11536) );
  nor2_1 U13205 ( .ip1(i_ssi_U_regfile_txflr[1]), .ip2(n11522), .op(n11534) );
  inv_1 U13206 ( .ip(n11522), .op(n11598) );
  nand2_1 U13207 ( .ip1(n11592), .ip2(n5351), .op(n11525) );
  nand2_1 U13208 ( .ip1(n11636), .ip2(i_ssi_U_regfile_ctrlr1_int[1]), .op(
        n11524) );
  nand2_1 U13209 ( .ip1(n11635), .ip2(i_ssi_baudr[1]), .op(n11523) );
  nand3_1 U13210 ( .ip1(n11525), .ip2(n11524), .ip3(n11523), .op(n11526) );
  mux2_1 U13211 ( .ip1(n11526), .ip2(i_ssi_mwcr[1]), .s(n11548), .op(n11528)
         );
  mux2_1 U13212 ( .ip1(i_ssi_txftlr[1]), .ip2(n11528), .s(n11527), .op(n11530)
         );
  mux2_1 U13213 ( .ip1(i_ssi_rxftlr[1]), .ip2(n11530), .s(n11529), .op(n11532)
         );
  nor2_1 U13214 ( .ip1(i_ssi_tx_full), .ip2(n11545), .op(n11531) );
  nor3_1 U13215 ( .ip1(n11598), .ip2(n11532), .ip3(n11531), .op(n11533) );
  nor2_1 U13216 ( .ip1(n11534), .ip2(n11533), .op(n11535) );
  not_ab_or_c_or_d U13217 ( .ip1(i_ssi_imr[1]), .ip2(n11640), .ip3(n11536), 
        .ip4(n11535), .op(n11541) );
  inv_1 U13218 ( .ip(n11537), .op(n11597) );
  inv_1 U13219 ( .ip(i_ssi_risr[1]), .op(n11538) );
  inv_1 U13220 ( .ip(n11641), .op(n11604) );
  nor2_1 U13221 ( .ip1(n11538), .ip2(n11604), .op(n11539) );
  not_ab_or_c_or_d U13222 ( .ip1(i_ssi_U_regfile_rxflr[1]), .ip2(n11597), 
        .ip3(n11661), .ip4(n11539), .op(n11540) );
  nand3_1 U13223 ( .ip1(n11542), .ip2(n11541), .ip3(n11540), .op(n11543) );
  mux2_1 U13224 ( .ip1(n11543), .ip2(i_ssi_prdata[1]), .s(n11663), .op(n4236)
         );
  nand2_1 U13225 ( .ip1(n11663), .ip2(i_ssi_prdata[2]), .op(n11577) );
  nor2_1 U13226 ( .ip1(n11634), .ip2(i_ssi_ssi_rxu_intr_n), .op(n11544) );
  not_ab_or_c_or_d U13227 ( .ip1(n11597), .ip2(i_ssi_U_regfile_rxflr[2]), 
        .ip3(n11661), .ip4(n11544), .op(n11562) );
  nor2_1 U13228 ( .ip1(i_ssi_U_fifo_U_tx_fifo_empty_n), .ip2(n11545), .op(
        n11554) );
  nand2_1 U13229 ( .ip1(n11546), .ip2(i_ssi_rxftlr[2]), .op(n11552) );
  nand2_1 U13230 ( .ip1(n11547), .ip2(i_ssi_txftlr[2]), .op(n11551) );
  nand2_1 U13231 ( .ip1(n11548), .ip2(i_ssi_mwcr[2]), .op(n11550) );
  nand2_1 U13232 ( .ip1(n11592), .ip2(n5353), .op(n11549) );
  nand4_1 U13233 ( .ip1(n11552), .ip2(n11551), .ip3(n11550), .ip4(n11549), 
        .op(n11553) );
  nor2_1 U13234 ( .ip1(n11554), .ip2(n11553), .op(n11558) );
  nand2_1 U13235 ( .ip1(n11598), .ip2(i_ssi_U_regfile_txflr[2]), .op(n11557)
         );
  nand2_1 U13236 ( .ip1(n11635), .ip2(i_ssi_baudr[2]), .op(n11556) );
  nand2_1 U13237 ( .ip1(n11636), .ip2(i_ssi_U_regfile_ctrlr1_int[2]), .op(
        n11555) );
  and4_1 U13238 ( .ip1(n11558), .ip2(n11557), .ip3(n11556), .ip4(n11555), .op(
        n11561) );
  nand2_1 U13239 ( .ip1(n11640), .ip2(i_ssi_imr[2]), .op(n11560) );
  nand2_1 U13240 ( .ip1(n11641), .ip2(i_ssi_risr[2]), .op(n11559) );
  nand4_1 U13241 ( .ip1(n11562), .ip2(n11561), .ip3(n11560), .ip4(n11559), 
        .op(n11563) );
  nand2_1 U13242 ( .ip1(n11651), .ip2(n11563), .op(n11576) );
  nand2_1 U13243 ( .ip1(n11620), .ip2(i_ssi_U_dff_rx_mem[2]), .op(n11573) );
  inv_1 U13244 ( .ip(i_ssi_U_dff_rx_mem[34]), .op(n11564) );
  nor2_1 U13245 ( .ip1(n11616), .ip2(n11564), .op(n11570) );
  nand2_1 U13246 ( .ip1(n11618), .ip2(i_ssi_U_dff_rx_mem[66]), .op(n11568) );
  nand2_1 U13247 ( .ip1(n11614), .ip2(i_ssi_U_dff_rx_mem[50]), .op(n11567) );
  nand2_1 U13248 ( .ip1(n11627), .ip2(i_ssi_U_dff_rx_mem[114]), .op(n11566) );
  nand2_1 U13249 ( .ip1(n11619), .ip2(i_ssi_U_dff_rx_mem[98]), .op(n11565) );
  nand4_1 U13250 ( .ip1(n11568), .ip2(n11567), .ip3(n11566), .ip4(n11565), 
        .op(n11569) );
  not_ab_or_c_or_d U13251 ( .ip1(i_ssi_U_dff_rx_mem[18]), .ip2(n11617), .ip3(
        n11570), .ip4(n11569), .op(n11572) );
  nand2_1 U13252 ( .ip1(n11628), .ip2(i_ssi_U_dff_rx_mem[82]), .op(n11571) );
  nand3_1 U13253 ( .ip1(n11573), .ip2(n11572), .ip3(n11571), .op(n11574) );
  nand2_1 U13254 ( .ip1(n6937), .ip2(n11574), .op(n11575) );
  nand3_1 U13255 ( .ip1(n11577), .ip2(n11576), .ip3(n11575), .op(n4235) );
  inv_1 U13256 ( .ip(i_ssi_U_dff_rx_mem[35]), .op(n11578) );
  nor2_1 U13257 ( .ip1(n11616), .ip2(n11578), .op(n11588) );
  nand2_1 U13258 ( .ip1(n11627), .ip2(i_ssi_U_dff_rx_mem[115]), .op(n11581) );
  nand2_1 U13259 ( .ip1(n11628), .ip2(i_ssi_U_dff_rx_mem[83]), .op(n11580) );
  nand2_1 U13260 ( .ip1(n11617), .ip2(i_ssi_U_dff_rx_mem[19]), .op(n11579) );
  nand3_1 U13261 ( .ip1(n11581), .ip2(n11580), .ip3(n11579), .op(n11587) );
  nand2_1 U13262 ( .ip1(n11618), .ip2(i_ssi_U_dff_rx_mem[67]), .op(n11585) );
  nand2_1 U13263 ( .ip1(n11619), .ip2(i_ssi_U_dff_rx_mem[99]), .op(n11584) );
  nand2_1 U13264 ( .ip1(n11614), .ip2(i_ssi_U_dff_rx_mem[51]), .op(n11583) );
  nand2_1 U13265 ( .ip1(n11620), .ip2(i_ssi_U_dff_rx_mem[3]), .op(n11582) );
  nand4_1 U13266 ( .ip1(n11585), .ip2(n11584), .ip3(n11583), .ip4(n11582), 
        .op(n11586) );
  nor3_1 U13267 ( .ip1(n11588), .ip2(n11587), .ip3(n11586), .op(n11589) );
  or2_1 U13268 ( .ip1(n11590), .ip2(n11589), .op(n11602) );
  nor2_1 U13269 ( .ip1(n6432), .ip2(n11591), .op(n11596) );
  nand2_1 U13270 ( .ip1(n11592), .ip2(n5453), .op(n11594) );
  nand2_1 U13271 ( .ip1(n11636), .ip2(i_ssi_U_regfile_ctrlr1_int[3]), .op(
        n11593) );
  nand2_1 U13272 ( .ip1(n11594), .ip2(n11593), .op(n11595) );
  not_ab_or_c_or_d U13273 ( .ip1(i_ssi_U_regfile_rxflr[3]), .ip2(n11597), 
        .ip3(n11596), .ip4(n11595), .op(n11601) );
  nand2_1 U13274 ( .ip1(n11647), .ip2(i_ssi_U_fifo_U_rx_fifo_empty_n), .op(
        n11600) );
  nand2_1 U13275 ( .ip1(n11598), .ip2(i_ssi_U_regfile_txflr[3]), .op(n11599)
         );
  and4_1 U13276 ( .ip1(n11602), .ip2(n11601), .ip3(n11600), .ip4(n11599), .op(
        n11612) );
  nor2_1 U13277 ( .ip1(i_ssi_ssi_rxo_intr_n), .ip2(n11603), .op(n11607) );
  nor2_1 U13278 ( .ip1(n11605), .ip2(n11604), .op(n11606) );
  nor2_1 U13279 ( .ip1(n11607), .ip2(n11606), .op(n11608) );
  nor2_1 U13280 ( .ip1(n11609), .ip2(n11608), .op(n11610) );
  not_ab_or_c_or_d U13281 ( .ip1(n11640), .ip2(i_ssi_imr[3]), .ip3(n11661), 
        .ip4(n11610), .op(n11611) );
  nand2_1 U13282 ( .ip1(n11612), .ip2(n11611), .op(n11613) );
  mux2_1 U13283 ( .ip1(n11613), .ip2(i_ssi_prdata[3]), .s(n11663), .op(n4234)
         );
  nand2_1 U13284 ( .ip1(n11614), .ip2(i_ssi_U_dff_rx_mem[52]), .op(n11631) );
  inv_1 U13285 ( .ip(i_ssi_U_dff_rx_mem[36]), .op(n11615) );
  nor2_1 U13286 ( .ip1(n11616), .ip2(n11615), .op(n11626) );
  nand2_1 U13287 ( .ip1(n11617), .ip2(i_ssi_U_dff_rx_mem[20]), .op(n11624) );
  nand2_1 U13288 ( .ip1(n11618), .ip2(i_ssi_U_dff_rx_mem[68]), .op(n11623) );
  nand2_1 U13289 ( .ip1(n11619), .ip2(i_ssi_U_dff_rx_mem[100]), .op(n11622) );
  nand2_1 U13290 ( .ip1(n11620), .ip2(i_ssi_U_dff_rx_mem[4]), .op(n11621) );
  nand4_1 U13291 ( .ip1(n11624), .ip2(n11623), .ip3(n11622), .ip4(n11621), 
        .op(n11625) );
  not_ab_or_c_or_d U13292 ( .ip1(i_ssi_U_dff_rx_mem[116]), .ip2(n11627), .ip3(
        n11626), .ip4(n11625), .op(n11630) );
  nand2_1 U13293 ( .ip1(n11628), .ip2(i_ssi_U_dff_rx_mem[84]), .op(n11629) );
  nand3_1 U13294 ( .ip1(n11631), .ip2(n11630), .ip3(n11629), .op(n11633) );
  nand2_1 U13295 ( .ip1(n11633), .ip2(n11632), .op(n11649) );
  nor2_1 U13296 ( .ip1(i_ssi_ssi_rxf_intr_n), .ip2(n11634), .op(n11646) );
  nand2_1 U13297 ( .ip1(n11635), .ip2(i_ssi_baudr[4]), .op(n11638) );
  nand2_1 U13298 ( .ip1(n11636), .ip2(i_ssi_U_regfile_ctrlr1_int[4]), .op(
        n11637) );
  nand2_1 U13299 ( .ip1(n11640), .ip2(i_ssi_imr[4]), .op(n11643) );
  nand2_1 U13300 ( .ip1(n11641), .ip2(i_ssi_risr[4]), .op(n11642) );
  nand4_1 U13301 ( .ip1(n11639), .ip2(n11644), .ip3(n11643), .ip4(n11642), 
        .op(n11645) );
  not_ab_or_c_or_d U13302 ( .ip1(n11647), .ip2(i_ssi_rx_full), .ip3(n11646), 
        .ip4(n11645), .op(n11648) );
  nand2_1 U13303 ( .ip1(n11649), .ip2(n11648), .op(n11650) );
  nand2_1 U13304 ( .ip1(n11651), .ip2(n11650), .op(n11653) );
  nand2_1 U13305 ( .ip1(i_ssi_prdata[4]), .ip2(n11663), .op(n11652) );
  nand2_1 U13306 ( .ip1(n11653), .ip2(n11652), .op(n4233) );
  nand2_1 U13307 ( .ip1(i_ssi_prdata[16]), .ip2(n11663), .op(n11654) );
  nand2_1 U13308 ( .ip1(n11665), .ip2(n11654), .op(n4221) );
  mux2_1 U13309 ( .ip1(i_ssi_prdata[17]), .ip2(n11661), .s(n6687), .op(n4220)
         );
  nand2_1 U13310 ( .ip1(i_ssi_prdata[18]), .ip2(n11663), .op(n11655) );
  nand2_1 U13311 ( .ip1(n11665), .ip2(n11655), .op(n4219) );
  nand2_1 U13312 ( .ip1(i_ssi_prdata[19]), .ip2(n11663), .op(n11656) );
  nand2_1 U13313 ( .ip1(n11665), .ip2(n11656), .op(n4218) );
  mux2_1 U13314 ( .ip1(i_ssi_prdata[20]), .ip2(n11661), .s(n6687), .op(n4217)
         );
  mux2_1 U13315 ( .ip1(i_ssi_prdata[21]), .ip2(n11661), .s(n6687), .op(n4216)
         );
  nand2_1 U13316 ( .ip1(i_ssi_prdata[22]), .ip2(n11663), .op(n11657) );
  nand2_1 U13317 ( .ip1(n11665), .ip2(n11657), .op(n4215) );
  nand2_1 U13318 ( .ip1(i_ssi_prdata[23]), .ip2(n11663), .op(n11658) );
  nand2_1 U13319 ( .ip1(n11665), .ip2(n11658), .op(n4214) );
  mux2_1 U13320 ( .ip1(i_ssi_prdata[24]), .ip2(n11661), .s(n6687), .op(n4213)
         );
  mux2_1 U13321 ( .ip1(i_ssi_prdata[25]), .ip2(n11661), .s(n6687), .op(n4212)
         );
  nand2_1 U13322 ( .ip1(i_ssi_prdata[26]), .ip2(n11663), .op(n11659) );
  nand2_1 U13323 ( .ip1(n11665), .ip2(n11659), .op(n4211) );
  nand2_1 U13324 ( .ip1(i_ssi_prdata[27]), .ip2(n11663), .op(n11660) );
  nand2_1 U13325 ( .ip1(n11665), .ip2(n11660), .op(n4210) );
  mux2_1 U13326 ( .ip1(i_ssi_prdata[28]), .ip2(n11661), .s(n6687), .op(n4209)
         );
  mux2_1 U13327 ( .ip1(i_ssi_prdata[29]), .ip2(n11661), .s(n6687), .op(n4208)
         );
  nand2_1 U13328 ( .ip1(i_ssi_prdata[30]), .ip2(n11663), .op(n11662) );
  nand2_1 U13329 ( .ip1(n11665), .ip2(n11662), .op(n4207) );
  nand2_1 U13330 ( .ip1(i_ssi_prdata[31]), .ip2(n11663), .op(n11664) );
  nand2_1 U13331 ( .ip1(n11665), .ip2(n11664), .op(n4206) );
  inv_1 U13332 ( .ip(i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[2]), .op(
        n11666) );
  nor2_1 U13333 ( .ip1(n11667), .ip2(n11666), .op(n11670) );
  not_ab_or_c_or_d U13334 ( .ip1(n11667), .ip2(n11666), .ip3(n11669), .ip4(
        n11670), .op(n4167) );
  nor2_1 U13335 ( .ip1(i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[3]), .ip2(
        n11670), .op(n11668) );
  not_ab_or_c_or_d U13336 ( .ip1(
        i_i2c_U_DW_apb_i2c_rx_shift_scl_hl_edg_cntr[3]), .ip2(n11670), .ip3(
        n11669), .ip4(n11668), .op(n4166) );
  nor2_1 U13337 ( .ip1(i_i2c_U_DW_apb_i2c_toggle_rx_gen_call_r), .ip2(n11671), 
        .op(n11672) );
  xor2_1 U13338 ( .ip1(i_i2c_rx_gen_call_flg), .ip2(n11672), .op(n4165) );
  xor2_1 U13339 ( .ip1(i_i2c_rx_push_flg), .ip2(i_i2c_rx_push), .op(n4163) );
  nor2_1 U13340 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(n11673), .op(n11695) );
  nand2_1 U13341 ( .ip1(n11695), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[0]), .op(n11676) );
  nor2_1 U13342 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(i_i2c_slv_rxbyte_rdy), .op(
        n11696) );
  nand2_1 U13343 ( .ip1(i_i2c_rx_push_data[0]), .ip2(n11696), .op(n11675) );
  nand2_1 U13344 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[0]), .op(n11674) );
  nand3_1 U13345 ( .ip1(n11676), .ip2(n11675), .ip3(n11674), .op(n4126) );
  nand2_1 U13346 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[1]), .op(n11679) );
  nand2_1 U13347 ( .ip1(n11695), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[1]), .op(n11678) );
  nand2_1 U13348 ( .ip1(i_i2c_rx_push_data[1]), .ip2(n11696), .op(n11677) );
  nand3_1 U13349 ( .ip1(n11679), .ip2(n11678), .ip3(n11677), .op(n4125) );
  nand2_1 U13350 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[2]), .op(n11682) );
  nand2_1 U13351 ( .ip1(n11695), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[2]), .op(n11681) );
  nand2_1 U13352 ( .ip1(i_i2c_rx_push_data[2]), .ip2(n11696), .op(n11680) );
  nand3_1 U13353 ( .ip1(n11682), .ip2(n11681), .ip3(n11680), .op(n4124) );
  nand2_1 U13354 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[3]), .op(n11685) );
  nand2_1 U13355 ( .ip1(n11695), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[3]), .op(n11684) );
  nand2_1 U13356 ( .ip1(i_i2c_rx_push_data[3]), .ip2(n11696), .op(n11683) );
  nand3_1 U13357 ( .ip1(n11685), .ip2(n11684), .ip3(n11683), .op(n4123) );
  nand2_1 U13358 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[4]), .op(n11688) );
  nand2_1 U13359 ( .ip1(n11695), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[4]), .op(n11687) );
  nand2_1 U13360 ( .ip1(i_i2c_rx_push_data[4]), .ip2(n11696), .op(n11686) );
  nand3_1 U13361 ( .ip1(n11688), .ip2(n11687), .ip3(n11686), .op(n4122) );
  nand2_1 U13362 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[5]), .op(n11691) );
  nand2_1 U13363 ( .ip1(n11695), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[5]), .op(n11690) );
  nand2_1 U13364 ( .ip1(i_i2c_rx_push_data[5]), .ip2(n11696), .op(n11689) );
  nand3_1 U13365 ( .ip1(n11691), .ip2(n11690), .ip3(n11689), .op(n4121) );
  nand2_1 U13366 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[6]), .op(n11694) );
  nand2_1 U13367 ( .ip1(n11695), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[6]), .op(n11693) );
  nand2_1 U13368 ( .ip1(i_i2c_rx_push_data[6]), .ip2(n11696), .op(n11692) );
  nand3_1 U13369 ( .ip1(n11694), .ip2(n11693), .ip3(n11692), .op(n4120) );
  nand2_1 U13370 ( .ip1(i_i2c_mst_rxbyte_rdy), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_mst_rx_shift_reg[7]), .op(n11699) );
  nand2_1 U13371 ( .ip1(n11695), .ip2(
        i_i2c_U_DW_apb_i2c_rx_shift_slv_rx_shift_reg[7]), .op(n11698) );
  nand2_1 U13372 ( .ip1(i_i2c_rx_push_data[7]), .ip2(n11696), .op(n11697) );
  nand3_1 U13373 ( .ip1(n11699), .ip2(n11698), .ip3(n11697), .op(n4119) );
  nor3_1 U13374 ( .ip1(i_i2c_rx_rd_addr[2]), .ip2(i_i2c_rx_rd_addr[0]), .ip3(
        n11704), .op(n11788) );
  nand2_1 U13375 ( .ip1(n11788), .ip2(i_i2c_U_dff_rx_mem[40]), .op(n11713) );
  inv_1 U13376 ( .ip(i_i2c_rx_rd_addr[2]), .op(n11703) );
  nor3_1 U13377 ( .ip1(i_i2c_rx_rd_addr[1]), .ip2(n11703), .ip3(n11701), .op(
        n11779) );
  inv_1 U13378 ( .ip(i_i2c_U_dff_rx_mem[0]), .op(n11700) );
  nand3_1 U13379 ( .ip1(i_i2c_rx_rd_addr[2]), .ip2(i_i2c_rx_rd_addr[1]), .ip3(
        i_i2c_rx_rd_addr[0]), .op(n11775) );
  nor2_1 U13380 ( .ip1(n11700), .ip2(n11775), .op(n11710) );
  nor3_1 U13381 ( .ip1(i_i2c_rx_rd_addr[2]), .ip2(i_i2c_rx_rd_addr[1]), .ip3(
        n11701), .op(n11778) );
  nand2_1 U13382 ( .ip1(i_i2c_U_dff_rx_mem[48]), .ip2(n11778), .op(n11708) );
  nor2_1 U13383 ( .ip1(i_i2c_rx_rd_addr[2]), .ip2(n11702), .op(n11787) );
  nand2_1 U13384 ( .ip1(i_i2c_U_dff_rx_mem[32]), .ip2(n11787), .op(n11707) );
  nor3_1 U13385 ( .ip1(i_i2c_rx_rd_addr[1]), .ip2(i_i2c_rx_rd_addr[0]), .ip3(
        n11703), .op(n11774) );
  nand2_1 U13386 ( .ip1(i_i2c_U_dff_rx_mem[24]), .ip2(n11774), .op(n11706) );
  nor3_1 U13387 ( .ip1(i_i2c_rx_rd_addr[0]), .ip2(n11704), .ip3(n11703), .op(
        n11780) );
  nand2_1 U13388 ( .ip1(i_i2c_U_dff_rx_mem[8]), .ip2(n11780), .op(n11705) );
  nand4_1 U13389 ( .ip1(n11708), .ip2(n11707), .ip3(n11706), .ip4(n11705), 
        .op(n11709) );
  not_ab_or_c_or_d U13390 ( .ip1(i_i2c_U_dff_rx_mem[16]), .ip2(n11779), .ip3(
        n11710), .ip4(n11709), .op(n11712) );
  nor3_1 U13391 ( .ip1(i_i2c_rx_rd_addr[2]), .ip2(i_i2c_rx_rd_addr[1]), .ip3(
        i_i2c_rx_rd_addr[0]), .op(n11777) );
  nand2_1 U13392 ( .ip1(i_i2c_U_dff_rx_mem[56]), .ip2(n11777), .op(n11711) );
  nand3_1 U13393 ( .ip1(n11713), .ip2(n11712), .ip3(n11711), .op(
        i_i2c_rx_pop_data[0]) );
  nand2_1 U13394 ( .ip1(i_i2c_U_dff_rx_mem[9]), .ip2(n11780), .op(n11723) );
  inv_1 U13395 ( .ip(i_i2c_U_dff_rx_mem[1]), .op(n11714) );
  nor2_1 U13396 ( .ip1(n11714), .ip2(n11775), .op(n11720) );
  nand2_1 U13397 ( .ip1(i_i2c_U_dff_rx_mem[57]), .ip2(n11777), .op(n11718) );
  nand2_1 U13398 ( .ip1(i_i2c_U_dff_rx_mem[33]), .ip2(n11787), .op(n11717) );
  nand2_1 U13399 ( .ip1(i_i2c_U_dff_rx_mem[17]), .ip2(n11779), .op(n11716) );
  nand2_1 U13400 ( .ip1(i_i2c_U_dff_rx_mem[41]), .ip2(n11788), .op(n11715) );
  nand4_1 U13401 ( .ip1(n11718), .ip2(n11717), .ip3(n11716), .ip4(n11715), 
        .op(n11719) );
  not_ab_or_c_or_d U13402 ( .ip1(n11778), .ip2(i_i2c_U_dff_rx_mem[49]), .ip3(
        n11720), .ip4(n11719), .op(n11722) );
  nand2_1 U13403 ( .ip1(i_i2c_U_dff_rx_mem[25]), .ip2(n11774), .op(n11721) );
  nand3_1 U13404 ( .ip1(n11723), .ip2(n11722), .ip3(n11721), .op(
        i_i2c_rx_pop_data[1]) );
  nand2_1 U13405 ( .ip1(i_i2c_U_dff_rx_mem[34]), .ip2(n11787), .op(n11733) );
  inv_1 U13406 ( .ip(i_i2c_U_dff_rx_mem[2]), .op(n11724) );
  nor2_1 U13407 ( .ip1(n11724), .ip2(n11775), .op(n11730) );
  nand2_1 U13408 ( .ip1(i_i2c_U_dff_rx_mem[26]), .ip2(n11774), .op(n11728) );
  nand2_1 U13409 ( .ip1(i_i2c_U_dff_rx_mem[18]), .ip2(n11779), .op(n11727) );
  nand2_1 U13410 ( .ip1(i_i2c_U_dff_rx_mem[50]), .ip2(n11778), .op(n11726) );
  nand2_1 U13411 ( .ip1(i_i2c_U_dff_rx_mem[42]), .ip2(n11788), .op(n11725) );
  nand4_1 U13412 ( .ip1(n11728), .ip2(n11727), .ip3(n11726), .ip4(n11725), 
        .op(n11729) );
  not_ab_or_c_or_d U13413 ( .ip1(n11780), .ip2(i_i2c_U_dff_rx_mem[10]), .ip3(
        n11730), .ip4(n11729), .op(n11732) );
  nand2_1 U13414 ( .ip1(i_i2c_U_dff_rx_mem[58]), .ip2(n11777), .op(n11731) );
  nand3_1 U13415 ( .ip1(n11733), .ip2(n11732), .ip3(n11731), .op(
        i_i2c_rx_pop_data[2]) );
  nand2_1 U13416 ( .ip1(i_i2c_U_dff_rx_mem[43]), .ip2(n11788), .op(n11743) );
  inv_1 U13417 ( .ip(i_i2c_U_dff_rx_mem[3]), .op(n11734) );
  nor2_1 U13418 ( .ip1(n11734), .ip2(n11775), .op(n11740) );
  nand2_1 U13419 ( .ip1(i_i2c_U_dff_rx_mem[27]), .ip2(n11774), .op(n11738) );
  nand2_1 U13420 ( .ip1(i_i2c_U_dff_rx_mem[11]), .ip2(n11780), .op(n11737) );
  nand2_1 U13421 ( .ip1(i_i2c_U_dff_rx_mem[35]), .ip2(n11787), .op(n11736) );
  nand2_1 U13422 ( .ip1(i_i2c_U_dff_rx_mem[59]), .ip2(n11777), .op(n11735) );
  nand4_1 U13423 ( .ip1(n11738), .ip2(n11737), .ip3(n11736), .ip4(n11735), 
        .op(n11739) );
  not_ab_or_c_or_d U13424 ( .ip1(n11779), .ip2(i_i2c_U_dff_rx_mem[19]), .ip3(
        n11740), .ip4(n11739), .op(n11742) );
  nand2_1 U13425 ( .ip1(i_i2c_U_dff_rx_mem[51]), .ip2(n11778), .op(n11741) );
  nand3_1 U13426 ( .ip1(n11743), .ip2(n11742), .ip3(n11741), .op(
        i_i2c_rx_pop_data[3]) );
  nand2_1 U13427 ( .ip1(i_i2c_U_dff_rx_mem[12]), .ip2(n11780), .op(n11753) );
  inv_1 U13428 ( .ip(i_i2c_U_dff_rx_mem[4]), .op(n11744) );
  nor2_1 U13429 ( .ip1(n11744), .ip2(n11775), .op(n11750) );
  nand2_1 U13430 ( .ip1(i_i2c_U_dff_rx_mem[52]), .ip2(n11778), .op(n11748) );
  nand2_1 U13431 ( .ip1(i_i2c_U_dff_rx_mem[28]), .ip2(n11774), .op(n11747) );
  nand2_1 U13432 ( .ip1(i_i2c_U_dff_rx_mem[44]), .ip2(n11788), .op(n11746) );
  nand2_1 U13433 ( .ip1(i_i2c_U_dff_rx_mem[60]), .ip2(n11777), .op(n11745) );
  nand4_1 U13434 ( .ip1(n11748), .ip2(n11747), .ip3(n11746), .ip4(n11745), 
        .op(n11749) );
  not_ab_or_c_or_d U13435 ( .ip1(n11787), .ip2(i_i2c_U_dff_rx_mem[36]), .ip3(
        n11750), .ip4(n11749), .op(n11752) );
  nand2_1 U13436 ( .ip1(i_i2c_U_dff_rx_mem[20]), .ip2(n11779), .op(n11751) );
  nand3_1 U13437 ( .ip1(n11753), .ip2(n11752), .ip3(n11751), .op(
        i_i2c_rx_pop_data[4]) );
  nand2_1 U13438 ( .ip1(i_i2c_U_dff_rx_mem[13]), .ip2(n11780), .op(n11763) );
  inv_1 U13439 ( .ip(i_i2c_U_dff_rx_mem[5]), .op(n11754) );
  nor2_1 U13440 ( .ip1(n11754), .ip2(n11775), .op(n11760) );
  nand2_1 U13441 ( .ip1(i_i2c_U_dff_rx_mem[37]), .ip2(n11787), .op(n11758) );
  nand2_1 U13442 ( .ip1(i_i2c_U_dff_rx_mem[53]), .ip2(n11778), .op(n11757) );
  nand2_1 U13443 ( .ip1(i_i2c_U_dff_rx_mem[61]), .ip2(n11777), .op(n11756) );
  nand2_1 U13444 ( .ip1(i_i2c_U_dff_rx_mem[45]), .ip2(n11788), .op(n11755) );
  nand4_1 U13445 ( .ip1(n11758), .ip2(n11757), .ip3(n11756), .ip4(n11755), 
        .op(n11759) );
  not_ab_or_c_or_d U13446 ( .ip1(n11779), .ip2(i_i2c_U_dff_rx_mem[21]), .ip3(
        n11760), .ip4(n11759), .op(n11762) );
  nand2_1 U13447 ( .ip1(i_i2c_U_dff_rx_mem[29]), .ip2(n11774), .op(n11761) );
  nand3_1 U13448 ( .ip1(n11763), .ip2(n11762), .ip3(n11761), .op(
        i_i2c_rx_pop_data[5]) );
  nand2_1 U13449 ( .ip1(i_i2c_U_dff_rx_mem[30]), .ip2(n11774), .op(n11773) );
  inv_1 U13450 ( .ip(i_i2c_U_dff_rx_mem[6]), .op(n11764) );
  nor2_1 U13451 ( .ip1(n11764), .ip2(n11775), .op(n11770) );
  nand2_1 U13452 ( .ip1(i_i2c_U_dff_rx_mem[54]), .ip2(n11778), .op(n11768) );
  nand2_1 U13453 ( .ip1(i_i2c_U_dff_rx_mem[22]), .ip2(n11779), .op(n11767) );
  nand2_1 U13454 ( .ip1(i_i2c_U_dff_rx_mem[62]), .ip2(n11777), .op(n11766) );
  nand2_1 U13455 ( .ip1(i_i2c_U_dff_rx_mem[14]), .ip2(n11780), .op(n11765) );
  nand4_1 U13456 ( .ip1(n11768), .ip2(n11767), .ip3(n11766), .ip4(n11765), 
        .op(n11769) );
  not_ab_or_c_or_d U13457 ( .ip1(n11787), .ip2(i_i2c_U_dff_rx_mem[38]), .ip3(
        n11770), .ip4(n11769), .op(n11772) );
  nand2_1 U13458 ( .ip1(i_i2c_U_dff_rx_mem[46]), .ip2(n11788), .op(n11771) );
  nand3_1 U13459 ( .ip1(n11773), .ip2(n11772), .ip3(n11771), .op(
        i_i2c_rx_pop_data[6]) );
  nand2_1 U13460 ( .ip1(i_i2c_U_dff_rx_mem[31]), .ip2(n11774), .op(n11791) );
  inv_1 U13461 ( .ip(i_i2c_U_dff_rx_mem[7]), .op(n11776) );
  nor2_1 U13462 ( .ip1(n11776), .ip2(n11775), .op(n11786) );
  nand2_1 U13463 ( .ip1(i_i2c_U_dff_rx_mem[63]), .ip2(n11777), .op(n11784) );
  nand2_1 U13464 ( .ip1(i_i2c_U_dff_rx_mem[55]), .ip2(n11778), .op(n11783) );
  nand2_1 U13465 ( .ip1(i_i2c_U_dff_rx_mem[23]), .ip2(n11779), .op(n11782) );
  nand2_1 U13466 ( .ip1(i_i2c_U_dff_rx_mem[15]), .ip2(n11780), .op(n11781) );
  nand4_1 U13467 ( .ip1(n11784), .ip2(n11783), .ip3(n11782), .ip4(n11781), 
        .op(n11785) );
  not_ab_or_c_or_d U13468 ( .ip1(n11787), .ip2(i_i2c_U_dff_rx_mem[39]), .ip3(
        n11786), .ip4(n11785), .op(n11790) );
  nand2_1 U13469 ( .ip1(i_i2c_U_dff_rx_mem[47]), .ip2(n11788), .op(n11789) );
  nand3_1 U13470 ( .ip1(n11791), .ip2(n11790), .ip3(n11789), .op(
        i_i2c_rx_pop_data[7]) );
endmodule

