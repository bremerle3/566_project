
module gen_pwm ( ap_clk, ap_rst, ap_start, ap_done, ap_idle, ap_ready, duty, 
        freq, out_r, out_r_ap_vld, ap_ce );
  input [31:0] duty;
  input [31:0] freq;
  output [0:0] out_r;
  input ap_clk, ap_rst, ap_start, ap_ce;
  output ap_done, ap_idle, ap_ready, out_r_ap_vld;
  wire   N60, n72, n73, n74, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498;
  wire   [1:0] ap_CS_fsm;
  wire   [30:0] i_reg_53;
  assign out_r[0] = N60;

  dp_1 \ap_CS_fsm_reg[0]  ( .ip(n73), .ck(ap_clk), .q(ap_CS_fsm[0]) );
  dp_1 \ap_CS_fsm_reg[1]  ( .ip(n72), .ck(ap_clk), .q(ap_CS_fsm[1]) );
  dp_1 \i_reg_53_reg[30]  ( .ip(n74), .ck(ap_clk), .q(i_reg_53[30]) );
  dp_1 \i_reg_53_reg[29]  ( .ip(n76), .ck(ap_clk), .q(i_reg_53[29]) );
  dp_1 \i_reg_53_reg[28]  ( .ip(n77), .ck(ap_clk), .q(i_reg_53[28]) );
  dp_1 \i_reg_53_reg[27]  ( .ip(n78), .ck(ap_clk), .q(i_reg_53[27]) );
  dp_1 \i_reg_53_reg[26]  ( .ip(n79), .ck(ap_clk), .q(i_reg_53[26]) );
  dp_1 \i_reg_53_reg[25]  ( .ip(n80), .ck(ap_clk), .q(i_reg_53[25]) );
  dp_1 \i_reg_53_reg[24]  ( .ip(n81), .ck(ap_clk), .q(i_reg_53[24]) );
  dp_1 \i_reg_53_reg[23]  ( .ip(n82), .ck(ap_clk), .q(i_reg_53[23]) );
  dp_1 \i_reg_53_reg[22]  ( .ip(n83), .ck(ap_clk), .q(i_reg_53[22]) );
  dp_1 \i_reg_53_reg[21]  ( .ip(n84), .ck(ap_clk), .q(i_reg_53[21]) );
  dp_1 \i_reg_53_reg[20]  ( .ip(n85), .ck(ap_clk), .q(i_reg_53[20]) );
  dp_1 \i_reg_53_reg[19]  ( .ip(n86), .ck(ap_clk), .q(i_reg_53[19]) );
  dp_1 \i_reg_53_reg[18]  ( .ip(n87), .ck(ap_clk), .q(i_reg_53[18]) );
  dp_1 \i_reg_53_reg[17]  ( .ip(n88), .ck(ap_clk), .q(i_reg_53[17]) );
  dp_1 \i_reg_53_reg[16]  ( .ip(n89), .ck(ap_clk), .q(i_reg_53[16]) );
  dp_1 \i_reg_53_reg[15]  ( .ip(n90), .ck(ap_clk), .q(i_reg_53[15]) );
  dp_1 \i_reg_53_reg[14]  ( .ip(n91), .ck(ap_clk), .q(i_reg_53[14]) );
  dp_1 \i_reg_53_reg[13]  ( .ip(n92), .ck(ap_clk), .q(i_reg_53[13]) );
  dp_1 \i_reg_53_reg[12]  ( .ip(n93), .ck(ap_clk), .q(i_reg_53[12]) );
  dp_1 \i_reg_53_reg[11]  ( .ip(n94), .ck(ap_clk), .q(i_reg_53[11]) );
  dp_1 \i_reg_53_reg[10]  ( .ip(n95), .ck(ap_clk), .q(i_reg_53[10]) );
  dp_1 \i_reg_53_reg[9]  ( .ip(n96), .ck(ap_clk), .q(i_reg_53[9]) );
  dp_1 \i_reg_53_reg[8]  ( .ip(n97), .ck(ap_clk), .q(i_reg_53[8]) );
  dp_1 \i_reg_53_reg[7]  ( .ip(n98), .ck(ap_clk), .q(i_reg_53[7]) );
  dp_1 \i_reg_53_reg[6]  ( .ip(n99), .ck(ap_clk), .q(i_reg_53[6]) );
  dp_1 \i_reg_53_reg[5]  ( .ip(n100), .ck(ap_clk), .q(i_reg_53[5]) );
  dp_1 \i_reg_53_reg[4]  ( .ip(n101), .ck(ap_clk), .q(i_reg_53[4]) );
  dp_1 \i_reg_53_reg[3]  ( .ip(n102), .ck(ap_clk), .q(i_reg_53[3]) );
  dp_1 \i_reg_53_reg[2]  ( .ip(n103), .ck(ap_clk), .q(i_reg_53[2]) );
  dp_1 \i_reg_53_reg[1]  ( .ip(n104), .ck(ap_clk), .q(i_reg_53[1]) );
  dp_1 \i_reg_53_reg[0]  ( .ip(n105), .ck(ap_clk), .q(i_reg_53[0]) );
  inv_1 U112 ( .ip(i_reg_53[27]), .op(n472) );
  inv_1 U113 ( .ip(i_reg_53[25]), .op(n464) );
  nor2_1 U114 ( .ip1(freq[25]), .ip2(n464), .op(n201) );
  inv_1 U115 ( .ip(n201), .op(n107) );
  inv_1 U116 ( .ip(i_reg_53[24]), .op(n463) );
  nand3_1 U117 ( .ip1(freq[24]), .ip2(n107), .ip3(n463), .op(n109) );
  nor2_1 U118 ( .ip1(freq[27]), .ip2(n472), .op(n114) );
  inv_1 U119 ( .ip(i_reg_53[26]), .op(n471) );
  nor2_1 U120 ( .ip1(freq[26]), .ip2(n471), .op(n108) );
  or2_1 U121 ( .ip1(n114), .ip2(n108), .op(n198) );
  or2_1 U122 ( .ip1(n109), .ip2(n198), .op(n112) );
  nand2_1 U123 ( .ip1(freq[25]), .ip2(n464), .op(n110) );
  or2_1 U124 ( .ip1(n110), .ip2(n198), .op(n111) );
  nand2_1 U125 ( .ip1(n112), .ip2(n111), .op(n116) );
  inv_1 U126 ( .ip(freq[26]), .op(n113) );
  nor3_1 U127 ( .ip1(n114), .ip2(i_reg_53[26]), .ip3(n113), .op(n115) );
  not_ab_or_c_or_d U128 ( .ip1(freq[27]), .ip2(n472), .ip3(n116), .ip4(n115), 
        .op(n120) );
  inv_1 U129 ( .ip(freq[28]), .op(n119) );
  inv_1 U130 ( .ip(i_reg_53[30]), .op(n324) );
  nor2_1 U131 ( .ip1(freq[30]), .ip2(n324), .op(n118) );
  inv_1 U132 ( .ip(i_reg_53[29]), .op(n484) );
  nor2_1 U133 ( .ip1(freq[29]), .ip2(n484), .op(n117) );
  or2_1 U134 ( .ip1(n118), .ip2(n117), .op(n207) );
  ab_or_c_or_d U135 ( .ip1(i_reg_53[28]), .ip2(n119), .ip3(freq[31]), .ip4(
        n207), .op(n202) );
  or2_1 U136 ( .ip1(n120), .ip2(n202), .op(n205) );
  inv_1 U137 ( .ip(i_reg_53[23]), .op(n454) );
  nor2_1 U138 ( .ip1(freq[23]), .ip2(n454), .op(n194) );
  inv_1 U139 ( .ip(i_reg_53[22]), .op(n453) );
  and2_1 U140 ( .ip1(n453), .ip2(freq[22]), .op(n192) );
  inv_1 U141 ( .ip(freq[20]), .op(n184) );
  inv_1 U142 ( .ip(i_reg_53[19]), .op(n434) );
  nor2_1 U143 ( .ip1(freq[19]), .ip2(n434), .op(n176) );
  inv_1 U144 ( .ip(freq[18]), .op(n121) );
  nor3_1 U145 ( .ip1(n176), .ip2(i_reg_53[18]), .ip3(n121), .op(n180) );
  inv_1 U146 ( .ip(i_reg_53[17]), .op(n429) );
  and2_1 U147 ( .ip1(n429), .ip2(freq[17]), .op(n174) );
  inv_1 U148 ( .ip(freq[16]), .op(n170) );
  inv_1 U149 ( .ip(i_reg_53[15]), .op(n411) );
  inv_1 U150 ( .ip(i_reg_53[11]), .op(n388) );
  nor2_1 U151 ( .ip1(freq[11]), .ip2(n388), .op(n154) );
  inv_1 U152 ( .ip(i_reg_53[10]), .op(n389) );
  and2_1 U153 ( .ip1(n389), .ip2(freq[10]), .op(n152) );
  inv_1 U154 ( .ip(i_reg_53[5]), .op(n356) );
  inv_1 U155 ( .ip(i_reg_53[1]), .op(n341) );
  nand2_1 U156 ( .ip1(freq[1]), .ip2(n341), .op(n124) );
  inv_1 U157 ( .ip(i_reg_53[0]), .op(n340) );
  or2_1 U158 ( .ip1(freq[1]), .ip2(n341), .op(n122) );
  nand3_1 U159 ( .ip1(n340), .ip2(freq[0]), .ip3(n122), .op(n123) );
  nand2_1 U160 ( .ip1(n124), .ip2(n123), .op(n125) );
  nand2_1 U161 ( .ip1(freq[2]), .ip2(n125), .op(n128) );
  inv_1 U162 ( .ip(i_reg_53[3]), .op(n343) );
  nor2_1 U163 ( .ip1(freq[3]), .ip2(n343), .op(n127) );
  nor2_1 U164 ( .ip1(freq[2]), .ip2(n125), .op(n126) );
  ab_or_c_or_d U165 ( .ip1(i_reg_53[2]), .ip2(n128), .ip3(n127), .ip4(n126), 
        .op(n131) );
  nand2_1 U166 ( .ip1(freq[3]), .ip2(n343), .op(n130) );
  inv_1 U167 ( .ip(i_reg_53[4]), .op(n355) );
  nor2_1 U168 ( .ip1(freq[4]), .ip2(n355), .op(n129) );
  nor2_1 U169 ( .ip1(freq[5]), .ip2(n356), .op(n133) );
  not_ab_or_c_or_d U170 ( .ip1(n131), .ip2(n130), .ip3(n129), .ip4(n133), .op(
        n135) );
  inv_1 U171 ( .ip(freq[4]), .op(n132) );
  nor3_1 U172 ( .ip1(n133), .ip2(i_reg_53[4]), .ip3(n132), .op(n134) );
  not_ab_or_c_or_d U173 ( .ip1(freq[5]), .ip2(n356), .ip3(n135), .ip4(n134), 
        .op(n139) );
  nor2_1 U174 ( .ip1(n139), .ip2(i_reg_53[6]), .op(n136) );
  nor2_1 U175 ( .ip1(freq[6]), .ip2(n136), .op(n138) );
  inv_1 U176 ( .ip(i_reg_53[7]), .op(n374) );
  nor2_1 U177 ( .ip1(freq[7]), .ip2(n374), .op(n137) );
  ab_or_c_or_d U178 ( .ip1(i_reg_53[6]), .ip2(n139), .ip3(n138), .ip4(n137), 
        .op(n144) );
  nand2_1 U179 ( .ip1(freq[7]), .ip2(n374), .op(n143) );
  inv_1 U180 ( .ip(i_reg_53[8]), .op(n375) );
  nor2_1 U181 ( .ip1(freq[8]), .ip2(n375), .op(n142) );
  nor2_1 U182 ( .ip1(freq[10]), .ip2(n389), .op(n141) );
  inv_1 U183 ( .ip(i_reg_53[9]), .op(n376) );
  nor2_1 U184 ( .ip1(freq[9]), .ip2(n376), .op(n140) );
  or2_1 U185 ( .ip1(n141), .ip2(n140), .op(n146) );
  not_ab_or_c_or_d U186 ( .ip1(n144), .ip2(n143), .ip3(n142), .ip4(n146), .op(
        n151) );
  nand2_1 U187 ( .ip1(freq[9]), .ip2(n376), .op(n145) );
  or2_1 U188 ( .ip1(n145), .ip2(n146), .op(n149) );
  nand2_1 U189 ( .ip1(freq[8]), .ip2(n375), .op(n147) );
  or2_1 U190 ( .ip1(n147), .ip2(n146), .op(n148) );
  nand2_1 U191 ( .ip1(n149), .ip2(n148), .op(n150) );
  nor3_1 U192 ( .ip1(n152), .ip2(n151), .ip3(n150), .op(n153) );
  nor2_1 U193 ( .ip1(n154), .ip2(n153), .op(n155) );
  or2_1 U194 ( .ip1(freq[11]), .ip2(n155), .op(n157) );
  or2_1 U195 ( .ip1(n388), .ip2(n155), .op(n156) );
  nand2_1 U196 ( .ip1(n157), .ip2(n156), .op(n161) );
  nor2_1 U197 ( .ip1(n161), .ip2(i_reg_53[12]), .op(n158) );
  nor2_1 U198 ( .ip1(freq[12]), .ip2(n158), .op(n160) );
  inv_1 U199 ( .ip(i_reg_53[13]), .op(n406) );
  nor2_1 U200 ( .ip1(freq[13]), .ip2(n406), .op(n159) );
  ab_or_c_or_d U201 ( .ip1(i_reg_53[12]), .ip2(n161), .ip3(n160), .ip4(n159), 
        .op(n164) );
  nand2_1 U202 ( .ip1(freq[13]), .ip2(n406), .op(n163) );
  inv_1 U203 ( .ip(i_reg_53[14]), .op(n410) );
  nor2_1 U204 ( .ip1(freq[14]), .ip2(n410), .op(n162) );
  nor2_1 U205 ( .ip1(freq[15]), .ip2(n411), .op(n166) );
  not_ab_or_c_or_d U206 ( .ip1(n164), .ip2(n163), .ip3(n162), .ip4(n166), .op(
        n168) );
  inv_1 U207 ( .ip(freq[14]), .op(n165) );
  nor3_1 U208 ( .ip1(n166), .ip2(i_reg_53[14]), .ip3(n165), .op(n167) );
  not_ab_or_c_or_d U209 ( .ip1(freq[15]), .ip2(n411), .ip3(n168), .ip4(n167), 
        .op(n169) );
  nor2_1 U210 ( .ip1(freq[17]), .ip2(n429), .op(n171) );
  not_ab_or_c_or_d U211 ( .ip1(i_reg_53[16]), .ip2(n170), .ip3(n169), .ip4(
        n171), .op(n173) );
  nor3_1 U212 ( .ip1(n171), .ip2(i_reg_53[16]), .ip3(n170), .op(n172) );
  nor3_1 U213 ( .ip1(n174), .ip2(n173), .ip3(n172), .op(n178) );
  inv_1 U214 ( .ip(i_reg_53[18]), .op(n433) );
  nor2_1 U215 ( .ip1(freq[18]), .ip2(n433), .op(n175) );
  or2_1 U216 ( .ip1(n176), .ip2(n175), .op(n177) );
  nor2_1 U217 ( .ip1(n178), .ip2(n177), .op(n179) );
  not_ab_or_c_or_d U218 ( .ip1(freq[19]), .ip2(n434), .ip3(n180), .ip4(n179), 
        .op(n183) );
  nor2_1 U219 ( .ip1(freq[22]), .ip2(n453), .op(n182) );
  inv_1 U220 ( .ip(i_reg_53[21]), .op(n443) );
  nor2_1 U221 ( .ip1(freq[21]), .ip2(n443), .op(n181) );
  or2_1 U222 ( .ip1(n182), .ip2(n181), .op(n186) );
  not_ab_or_c_or_d U223 ( .ip1(i_reg_53[20]), .ip2(n184), .ip3(n183), .ip4(
        n186), .op(n191) );
  nand2_1 U224 ( .ip1(freq[21]), .ip2(n443), .op(n185) );
  or2_1 U225 ( .ip1(n185), .ip2(n186), .op(n189) );
  inv_1 U226 ( .ip(i_reg_53[20]), .op(n444) );
  nand2_1 U227 ( .ip1(freq[20]), .ip2(n444), .op(n187) );
  or2_1 U228 ( .ip1(n187), .ip2(n186), .op(n188) );
  nand2_1 U229 ( .ip1(n189), .ip2(n188), .op(n190) );
  nor3_1 U230 ( .ip1(n192), .ip2(n191), .ip3(n190), .op(n193) );
  nor2_1 U231 ( .ip1(n194), .ip2(n193), .op(n195) );
  or2_1 U232 ( .ip1(freq[23]), .ip2(n195), .op(n197) );
  or2_1 U233 ( .ip1(n454), .ip2(n195), .op(n196) );
  nand2_1 U234 ( .ip1(n197), .ip2(n196), .op(n200) );
  nor2_1 U235 ( .ip1(freq[24]), .ip2(n463), .op(n199) );
  or4_1 U236 ( .ip1(n201), .ip2(n200), .ip3(n199), .ip4(n198), .op(n203) );
  or2_1 U237 ( .ip1(n203), .ip2(n202), .op(n204) );
  nand2_1 U238 ( .ip1(n205), .ip2(n204), .op(n216) );
  nand2_1 U239 ( .ip1(freq[29]), .ip2(n484), .op(n206) );
  or2_1 U240 ( .ip1(n206), .ip2(n207), .op(n210) );
  inv_1 U241 ( .ip(i_reg_53[28]), .op(n483) );
  nand2_1 U242 ( .ip1(freq[28]), .ip2(n483), .op(n208) );
  or2_1 U243 ( .ip1(n208), .ip2(n207), .op(n209) );
  nand2_1 U244 ( .ip1(n210), .ip2(n209), .op(n211) );
  or2_1 U245 ( .ip1(freq[30]), .ip2(n211), .op(n213) );
  or2_1 U246 ( .ip1(n324), .ip2(n211), .op(n212) );
  nand2_1 U247 ( .ip1(n213), .ip2(n212), .op(n214) );
  nor2_1 U248 ( .ip1(freq[31]), .ip2(n214), .op(n215) );
  nor2_1 U249 ( .ip1(n216), .ip2(n215), .op(n219) );
  inv_1 U250 ( .ip(n219), .op(n495) );
  nand2_1 U251 ( .ip1(ap_ce), .ip2(ap_CS_fsm[1]), .op(n218) );
  nor2_1 U252 ( .ip1(n495), .ip2(n218), .op(ap_done) );
  inv_1 U253 ( .ip(ap_done), .op(n217) );
  inv_1 U254 ( .ip(n217), .op(ap_ready) );
  nor2_1 U255 ( .ip1(n219), .ip2(n218), .op(out_r_ap_vld) );
  nor2_1 U256 ( .ip1(duty[25]), .ip2(n464), .op(n302) );
  nor2_1 U257 ( .ip1(duty[23]), .ip2(n454), .op(n293) );
  and2_1 U258 ( .ip1(n453), .ip2(duty[22]), .op(n291) );
  inv_1 U259 ( .ip(duty[20]), .op(n283) );
  inv_1 U260 ( .ip(duty[18]), .op(n220) );
  nor2_1 U261 ( .ip1(duty[19]), .ip2(n434), .op(n275) );
  nor3_1 U262 ( .ip1(n220), .ip2(i_reg_53[18]), .ip3(n275), .op(n279) );
  and2_1 U263 ( .ip1(n429), .ip2(duty[17]), .op(n273) );
  inv_1 U264 ( .ip(duty[16]), .op(n270) );
  nor2_1 U265 ( .ip1(duty[17]), .ip2(n429), .op(n269) );
  inv_1 U266 ( .ip(duty[14]), .op(n221) );
  nor2_1 U267 ( .ip1(duty[15]), .ip2(n411), .op(n262) );
  nor3_1 U268 ( .ip1(n221), .ip2(i_reg_53[14]), .ip3(n262), .op(n267) );
  nor2_1 U269 ( .ip1(duty[11]), .ip2(n388), .op(n254) );
  and2_1 U270 ( .ip1(n389), .ip2(duty[10]), .op(n252) );
  nor2_1 U271 ( .ip1(duty[8]), .ip2(n375), .op(n243) );
  inv_1 U272 ( .ip(duty[6]), .op(n238) );
  nor2_1 U273 ( .ip1(duty[7]), .ip2(n374), .op(n237) );
  nor3_1 U274 ( .ip1(n238), .ip2(i_reg_53[6]), .ip3(n237), .op(n240) );
  inv_1 U275 ( .ip(duty[4]), .op(n222) );
  nor2_1 U276 ( .ip1(duty[5]), .ip2(n356), .op(n230) );
  nor3_1 U277 ( .ip1(n222), .ip2(i_reg_53[4]), .ip3(n230), .op(n235) );
  nand2_1 U278 ( .ip1(duty[1]), .ip2(n341), .op(n225) );
  or2_1 U279 ( .ip1(duty[1]), .ip2(n341), .op(n223) );
  nand3_1 U280 ( .ip1(n340), .ip2(duty[0]), .ip3(n223), .op(n224) );
  nand2_1 U281 ( .ip1(n225), .ip2(n224), .op(n226) );
  nand2_1 U282 ( .ip1(duty[2]), .ip2(n226), .op(n229) );
  nor2_1 U283 ( .ip1(duty[3]), .ip2(n343), .op(n228) );
  nor2_1 U284 ( .ip1(duty[2]), .ip2(n226), .op(n227) );
  ab_or_c_or_d U285 ( .ip1(i_reg_53[2]), .ip2(n229), .ip3(n228), .ip4(n227), 
        .op(n233) );
  nand2_1 U286 ( .ip1(duty[3]), .ip2(n343), .op(n232) );
  nor2_1 U287 ( .ip1(duty[4]), .ip2(n355), .op(n231) );
  not_ab_or_c_or_d U288 ( .ip1(n233), .ip2(n232), .ip3(n231), .ip4(n230), .op(
        n234) );
  not_ab_or_c_or_d U289 ( .ip1(duty[5]), .ip2(n356), .ip3(n235), .ip4(n234), 
        .op(n236) );
  not_ab_or_c_or_d U290 ( .ip1(i_reg_53[6]), .ip2(n238), .ip3(n237), .ip4(n236), .op(n239) );
  not_ab_or_c_or_d U291 ( .ip1(duty[7]), .ip2(n374), .ip3(n240), .ip4(n239), 
        .op(n242) );
  nor2_1 U292 ( .ip1(duty[9]), .ip2(n376), .op(n241) );
  nor2_1 U293 ( .ip1(duty[10]), .ip2(n389), .op(n248) );
  nor4_1 U294 ( .ip1(n243), .ip2(n242), .ip3(n241), .ip4(n248), .op(n251) );
  nand2_1 U295 ( .ip1(duty[8]), .ip2(n375), .op(n249) );
  inv_1 U296 ( .ip(n249), .op(n244) );
  or2_1 U297 ( .ip1(n244), .ip2(duty[9]), .op(n246) );
  or2_1 U298 ( .ip1(n376), .ip2(duty[9]), .op(n245) );
  nand2_1 U299 ( .ip1(n246), .ip2(n245), .op(n247) );
  not_ab_or_c_or_d U300 ( .ip1(i_reg_53[9]), .ip2(n249), .ip3(n248), .ip4(n247), .op(n250) );
  nor3_1 U301 ( .ip1(n252), .ip2(n251), .ip3(n250), .op(n253) );
  nor2_1 U302 ( .ip1(n254), .ip2(n253), .op(n255) );
  or2_1 U303 ( .ip1(duty[11]), .ip2(n255), .op(n257) );
  or2_1 U304 ( .ip1(n388), .ip2(n255), .op(n256) );
  nand2_1 U305 ( .ip1(n257), .ip2(n256), .op(n261) );
  nor2_1 U306 ( .ip1(i_reg_53[12]), .ip2(n261), .op(n258) );
  nor2_1 U307 ( .ip1(duty[12]), .ip2(n258), .op(n260) );
  nor2_1 U308 ( .ip1(duty[13]), .ip2(n406), .op(n259) );
  ab_or_c_or_d U309 ( .ip1(n261), .ip2(i_reg_53[12]), .ip3(n260), .ip4(n259), 
        .op(n265) );
  nand2_1 U310 ( .ip1(duty[13]), .ip2(n406), .op(n264) );
  nor2_1 U311 ( .ip1(duty[14]), .ip2(n410), .op(n263) );
  not_ab_or_c_or_d U312 ( .ip1(n265), .ip2(n264), .ip3(n263), .ip4(n262), .op(
        n266) );
  not_ab_or_c_or_d U313 ( .ip1(duty[15]), .ip2(n411), .ip3(n267), .ip4(n266), 
        .op(n268) );
  not_ab_or_c_or_d U314 ( .ip1(i_reg_53[16]), .ip2(n270), .ip3(n269), .ip4(
        n268), .op(n272) );
  nor3_1 U315 ( .ip1(n270), .ip2(i_reg_53[16]), .ip3(n269), .op(n271) );
  nor3_1 U316 ( .ip1(n273), .ip2(n272), .ip3(n271), .op(n277) );
  nor2_1 U317 ( .ip1(duty[18]), .ip2(n433), .op(n274) );
  or2_1 U318 ( .ip1(n275), .ip2(n274), .op(n276) );
  nor2_1 U319 ( .ip1(n277), .ip2(n276), .op(n278) );
  not_ab_or_c_or_d U320 ( .ip1(duty[19]), .ip2(n434), .ip3(n279), .ip4(n278), 
        .op(n282) );
  nor2_1 U321 ( .ip1(duty[21]), .ip2(n443), .op(n281) );
  nor2_1 U322 ( .ip1(duty[22]), .ip2(n453), .op(n280) );
  or2_1 U323 ( .ip1(n281), .ip2(n280), .op(n285) );
  not_ab_or_c_or_d U324 ( .ip1(i_reg_53[20]), .ip2(n283), .ip3(n282), .ip4(
        n285), .op(n290) );
  nand2_1 U325 ( .ip1(duty[20]), .ip2(n444), .op(n284) );
  or2_1 U326 ( .ip1(n284), .ip2(n285), .op(n288) );
  nand2_1 U327 ( .ip1(duty[21]), .ip2(n443), .op(n286) );
  or2_1 U328 ( .ip1(n286), .ip2(n285), .op(n287) );
  nand2_1 U329 ( .ip1(n288), .ip2(n287), .op(n289) );
  nor3_1 U330 ( .ip1(n291), .ip2(n290), .ip3(n289), .op(n292) );
  nor2_1 U331 ( .ip1(n293), .ip2(n292), .op(n294) );
  or2_1 U332 ( .ip1(duty[23]), .ip2(n294), .op(n296) );
  or2_1 U333 ( .ip1(n454), .ip2(n294), .op(n295) );
  nand2_1 U334 ( .ip1(n296), .ip2(n295), .op(n299) );
  nor2_1 U335 ( .ip1(duty[24]), .ip2(n463), .op(n298) );
  nor2_1 U336 ( .ip1(duty[27]), .ip2(n472), .op(n300) );
  nor2_1 U337 ( .ip1(duty[26]), .ip2(n471), .op(n297) );
  or2_1 U338 ( .ip1(n300), .ip2(n297), .op(n305) );
  or4_1 U339 ( .ip1(n302), .ip2(n299), .ip3(n298), .ip4(n305), .op(n312) );
  inv_1 U340 ( .ip(duty[26]), .op(n301) );
  nor3_1 U341 ( .ip1(n301), .ip2(i_reg_53[26]), .ip3(n300), .op(n310) );
  inv_1 U342 ( .ip(n302), .op(n303) );
  nand3_1 U343 ( .ip1(duty[24]), .ip2(n463), .ip3(n303), .op(n304) );
  or2_1 U344 ( .ip1(n304), .ip2(n305), .op(n308) );
  nand2_1 U345 ( .ip1(duty[25]), .ip2(n464), .op(n306) );
  or2_1 U346 ( .ip1(n306), .ip2(n305), .op(n307) );
  nand2_1 U347 ( .ip1(n308), .ip2(n307), .op(n309) );
  not_ab_or_c_or_d U348 ( .ip1(duty[27]), .ip2(n472), .ip3(n310), .ip4(n309), 
        .op(n311) );
  nand2_1 U349 ( .ip1(n312), .ip2(n311), .op(n317) );
  inv_1 U350 ( .ip(duty[28]), .op(n315) );
  nor2_1 U351 ( .ip1(duty[29]), .ip2(n484), .op(n314) );
  nor2_1 U352 ( .ip1(duty[30]), .ip2(n324), .op(n313) );
  or2_1 U353 ( .ip1(n314), .ip2(n313), .op(n319) );
  not_ab_or_c_or_d U354 ( .ip1(i_reg_53[28]), .ip2(n315), .ip3(duty[31]), 
        .ip4(n319), .op(n316) );
  nand2_1 U355 ( .ip1(n317), .ip2(n316), .op(n329) );
  nand2_1 U356 ( .ip1(duty[28]), .ip2(n483), .op(n318) );
  or2_1 U357 ( .ip1(n318), .ip2(n319), .op(n322) );
  nand2_1 U358 ( .ip1(duty[29]), .ip2(n484), .op(n320) );
  or2_1 U359 ( .ip1(n320), .ip2(n319), .op(n321) );
  nand2_1 U360 ( .ip1(n322), .ip2(n321), .op(n323) );
  or2_1 U361 ( .ip1(duty[30]), .ip2(n323), .op(n326) );
  or2_1 U362 ( .ip1(n324), .ip2(n323), .op(n325) );
  nand2_1 U363 ( .ip1(n326), .ip2(n325), .op(n327) );
  or2_1 U364 ( .ip1(duty[31]), .ip2(n327), .op(n328) );
  nand2_1 U365 ( .ip1(n329), .ip2(n328), .op(N60) );
  inv_1 U366 ( .ip(ap_CS_fsm[0]), .op(n494) );
  nor2_1 U367 ( .ip1(ap_start), .ip2(n494), .op(ap_idle) );
  nand2_1 U368 ( .ip1(ap_start), .ip2(ap_CS_fsm[0]), .op(n490) );
  inv_1 U369 ( .ip(ap_ce), .op(n498) );
  or2_1 U370 ( .ip1(n490), .ip2(n498), .op(n492) );
  nand2_1 U371 ( .ip1(ap_CS_fsm[1]), .ip2(n495), .op(n330) );
  or2_1 U372 ( .ip1(n330), .ip2(n498), .op(n331) );
  nand2_1 U373 ( .ip1(n492), .ip2(n331), .op(n346) );
  inv_1 U374 ( .ip(n346), .op(n476) );
  mux2_1 U375 ( .ip1(out_r_ap_vld), .ip2(n476), .s(i_reg_53[0]), .op(n105) );
  nand2_1 U376 ( .ip1(out_r_ap_vld), .ip2(n340), .op(n332) );
  nand2_1 U377 ( .ip1(n346), .ip2(n332), .op(n334) );
  nor2_1 U378 ( .ip1(n340), .ip2(n428), .op(n333) );
  mux2_1 U379 ( .ip1(n334), .ip2(n333), .s(n341), .op(n104) );
  nor3_1 U380 ( .ip1(n341), .ip2(n340), .ip3(n428), .op(n337) );
  nor2_1 U381 ( .ip1(i_reg_53[1]), .ip2(n428), .op(n335) );
  nor2_1 U382 ( .ip1(n335), .ip2(n334), .op(n339) );
  inv_1 U383 ( .ip(n339), .op(n336) );
  mux2_1 U384 ( .ip1(n337), .ip2(n336), .s(i_reg_53[2]), .op(n103) );
  inv_1 U385 ( .ip(i_reg_53[2]), .op(n342) );
  nand2_1 U386 ( .ip1(out_r_ap_vld), .ip2(n342), .op(n338) );
  nand2_1 U387 ( .ip1(n339), .ip2(n338), .op(n345) );
  inv_1 U388 ( .ip(out_r_ap_vld), .op(n428) );
  nor4_1 U389 ( .ip1(n342), .ip2(n341), .ip3(n340), .ip4(n428), .op(n344) );
  mux2_1 U390 ( .ip1(n345), .ip2(n344), .s(n343), .op(n102) );
  nand2_1 U391 ( .ip1(out_r_ap_vld), .ip2(n355), .op(n350) );
  nand4_1 U392 ( .ip1(i_reg_53[3]), .ip2(i_reg_53[2]), .ip3(i_reg_53[1]), 
        .ip4(i_reg_53[0]), .op(n354) );
  nor2_1 U393 ( .ip1(n350), .ip2(n354), .op(n349) );
  nand2_1 U394 ( .ip1(n346), .ip2(n428), .op(n487) );
  or2_1 U395 ( .ip1(n354), .ip2(n476), .op(n347) );
  nand2_1 U396 ( .ip1(n487), .ip2(n347), .op(n351) );
  nor2_1 U397 ( .ip1(n351), .ip2(n355), .op(n348) );
  or2_1 U398 ( .ip1(n349), .ip2(n348), .op(n101) );
  nor3_1 U399 ( .ip1(n355), .ip2(n428), .ip3(n354), .op(n353) );
  nand2_1 U400 ( .ip1(n351), .ip2(n350), .op(n352) );
  mux2_1 U401 ( .ip1(n353), .ip2(n352), .s(i_reg_53[5]), .op(n100) );
  inv_1 U402 ( .ip(i_reg_53[6]), .op(n359) );
  nand2_1 U403 ( .ip1(out_r_ap_vld), .ip2(n359), .op(n362) );
  nor3_1 U404 ( .ip1(n356), .ip2(n355), .ip3(n354), .op(n364) );
  inv_1 U405 ( .ip(n364), .op(n357) );
  nor2_1 U406 ( .ip1(n362), .ip2(n357), .op(n361) );
  or2_1 U407 ( .ip1(n357), .ip2(n476), .op(n358) );
  nand2_1 U408 ( .ip1(n487), .ip2(n358), .op(n363) );
  nor2_1 U409 ( .ip1(n363), .ip2(n359), .op(n360) );
  or2_1 U410 ( .ip1(n361), .ip2(n360), .op(n99) );
  nand2_1 U411 ( .ip1(n363), .ip2(n362), .op(n366) );
  nand2_1 U412 ( .ip1(i_reg_53[6]), .ip2(n364), .op(n373) );
  nor2_1 U413 ( .ip1(n428), .ip2(n373), .op(n365) );
  mux2_1 U414 ( .ip1(n366), .ip2(n365), .s(n374), .op(n98) );
  nand2_1 U415 ( .ip1(out_r_ap_vld), .ip2(n375), .op(n371) );
  nor2_1 U416 ( .ip1(n374), .ip2(n373), .op(n379) );
  inv_1 U417 ( .ip(n379), .op(n367) );
  nor2_1 U418 ( .ip1(n371), .ip2(n367), .op(n370) );
  or2_1 U419 ( .ip1(n367), .ip2(n476), .op(n368) );
  nand2_1 U420 ( .ip1(n487), .ip2(n368), .op(n372) );
  nor2_1 U421 ( .ip1(n372), .ip2(n375), .op(n369) );
  or2_1 U422 ( .ip1(n370), .ip2(n369), .op(n97) );
  nand2_1 U423 ( .ip1(n372), .ip2(n371), .op(n378) );
  nor4_1 U424 ( .ip1(n375), .ip2(n374), .ip3(n428), .ip4(n373), .op(n377) );
  mux2_1 U425 ( .ip1(n378), .ip2(n377), .s(n376), .op(n96) );
  nand2_1 U426 ( .ip1(out_r_ap_vld), .ip2(n389), .op(n383) );
  nand3_1 U427 ( .ip1(i_reg_53[9]), .ip2(i_reg_53[8]), .ip3(n379), .op(n387)
         );
  nor2_1 U428 ( .ip1(n383), .ip2(n387), .op(n382) );
  or2_1 U429 ( .ip1(n387), .ip2(n476), .op(n380) );
  nand2_1 U430 ( .ip1(n487), .ip2(n380), .op(n384) );
  nor2_1 U431 ( .ip1(n384), .ip2(n389), .op(n381) );
  or2_1 U432 ( .ip1(n382), .ip2(n381), .op(n95) );
  nand2_1 U433 ( .ip1(n384), .ip2(n383), .op(n386) );
  nor3_1 U434 ( .ip1(n389), .ip2(n428), .ip3(n387), .op(n385) );
  mux2_1 U435 ( .ip1(n386), .ip2(n385), .s(n388), .op(n94) );
  inv_1 U436 ( .ip(i_reg_53[12]), .op(n392) );
  nand2_1 U437 ( .ip1(out_r_ap_vld), .ip2(n392), .op(n395) );
  nor3_1 U438 ( .ip1(n389), .ip2(n388), .ip3(n387), .op(n397) );
  inv_1 U439 ( .ip(n397), .op(n390) );
  nor2_1 U440 ( .ip1(n395), .ip2(n390), .op(n394) );
  or2_1 U441 ( .ip1(n390), .ip2(n476), .op(n391) );
  nand2_1 U442 ( .ip1(n487), .ip2(n391), .op(n396) );
  nor2_1 U443 ( .ip1(n396), .ip2(n392), .op(n393) );
  or2_1 U444 ( .ip1(n394), .ip2(n393), .op(n93) );
  nand2_1 U445 ( .ip1(n396), .ip2(n395), .op(n399) );
  nand2_1 U446 ( .ip1(i_reg_53[12]), .ip2(n397), .op(n405) );
  nor2_1 U447 ( .ip1(n428), .ip2(n405), .op(n398) );
  mux2_1 U448 ( .ip1(n399), .ip2(n398), .s(n406), .op(n92) );
  nand2_1 U449 ( .ip1(out_r_ap_vld), .ip2(n410), .op(n403) );
  or2_1 U450 ( .ip1(n406), .ip2(n405), .op(n409) );
  nor2_1 U451 ( .ip1(n403), .ip2(n409), .op(n402) );
  or2_1 U452 ( .ip1(n409), .ip2(n476), .op(n400) );
  nand2_1 U453 ( .ip1(n487), .ip2(n400), .op(n404) );
  nor2_1 U454 ( .ip1(n404), .ip2(n410), .op(n401) );
  or2_1 U455 ( .ip1(n402), .ip2(n401), .op(n91) );
  nand2_1 U456 ( .ip1(n404), .ip2(n403), .op(n408) );
  nor4_1 U457 ( .ip1(n406), .ip2(n410), .ip3(n428), .ip4(n405), .op(n407) );
  mux2_1 U458 ( .ip1(n408), .ip2(n407), .s(n411), .op(n90) );
  inv_1 U459 ( .ip(i_reg_53[16]), .op(n414) );
  nand2_1 U460 ( .ip1(out_r_ap_vld), .ip2(n414), .op(n417) );
  nor3_1 U461 ( .ip1(n411), .ip2(n410), .ip3(n409), .op(n419) );
  inv_1 U462 ( .ip(n419), .op(n412) );
  nor2_1 U463 ( .ip1(n417), .ip2(n412), .op(n416) );
  or2_1 U464 ( .ip1(n412), .ip2(n476), .op(n413) );
  nand2_1 U465 ( .ip1(n487), .ip2(n413), .op(n418) );
  nor2_1 U466 ( .ip1(n418), .ip2(n414), .op(n415) );
  or2_1 U467 ( .ip1(n416), .ip2(n415), .op(n89) );
  nand2_1 U468 ( .ip1(n418), .ip2(n417), .op(n421) );
  nand2_1 U469 ( .ip1(i_reg_53[16]), .ip2(n419), .op(n427) );
  nor2_1 U470 ( .ip1(n428), .ip2(n427), .op(n420) );
  mux2_1 U471 ( .ip1(n421), .ip2(n420), .s(n429), .op(n88) );
  nand2_1 U472 ( .ip1(out_r_ap_vld), .ip2(n433), .op(n425) );
  or2_1 U473 ( .ip1(n429), .ip2(n427), .op(n432) );
  nor2_1 U474 ( .ip1(n425), .ip2(n432), .op(n424) );
  or2_1 U475 ( .ip1(n432), .ip2(n476), .op(n422) );
  nand2_1 U476 ( .ip1(n487), .ip2(n422), .op(n426) );
  nor2_1 U477 ( .ip1(n426), .ip2(n433), .op(n423) );
  or2_1 U478 ( .ip1(n424), .ip2(n423), .op(n87) );
  nand2_1 U479 ( .ip1(n426), .ip2(n425), .op(n431) );
  nor4_1 U480 ( .ip1(n429), .ip2(n433), .ip3(n428), .ip4(n427), .op(n430) );
  mux2_1 U481 ( .ip1(n431), .ip2(n430), .s(n434), .op(n86) );
  nand2_1 U482 ( .ip1(out_r_ap_vld), .ip2(n444), .op(n438) );
  or3_1 U483 ( .ip1(n434), .ip2(n433), .ip3(n432), .op(n442) );
  nor2_1 U484 ( .ip1(n438), .ip2(n442), .op(n437) );
  or2_1 U485 ( .ip1(n442), .ip2(n476), .op(n435) );
  nand2_1 U486 ( .ip1(n487), .ip2(n435), .op(n439) );
  nor2_1 U487 ( .ip1(n439), .ip2(n444), .op(n436) );
  or2_1 U488 ( .ip1(n437), .ip2(n436), .op(n85) );
  nand2_1 U489 ( .ip1(n439), .ip2(n438), .op(n441) );
  nor3_1 U490 ( .ip1(n444), .ip2(n428), .ip3(n442), .op(n440) );
  mux2_1 U491 ( .ip1(n441), .ip2(n440), .s(n443), .op(n84) );
  nand2_1 U492 ( .ip1(out_r_ap_vld), .ip2(n453), .op(n448) );
  or3_1 U493 ( .ip1(n444), .ip2(n443), .ip3(n442), .op(n452) );
  nor2_1 U494 ( .ip1(n448), .ip2(n452), .op(n447) );
  or2_1 U495 ( .ip1(n452), .ip2(n476), .op(n445) );
  nand2_1 U496 ( .ip1(n487), .ip2(n445), .op(n449) );
  nor2_1 U497 ( .ip1(n449), .ip2(n453), .op(n446) );
  or2_1 U498 ( .ip1(n447), .ip2(n446), .op(n83) );
  nand2_1 U499 ( .ip1(n449), .ip2(n448), .op(n451) );
  nor3_1 U500 ( .ip1(n453), .ip2(n428), .ip3(n452), .op(n450) );
  mux2_1 U501 ( .ip1(n451), .ip2(n450), .s(n454), .op(n82) );
  nand2_1 U502 ( .ip1(out_r_ap_vld), .ip2(n463), .op(n458) );
  or3_1 U503 ( .ip1(n454), .ip2(n453), .ip3(n452), .op(n462) );
  nor2_1 U504 ( .ip1(n458), .ip2(n462), .op(n457) );
  or2_1 U505 ( .ip1(n462), .ip2(n476), .op(n455) );
  nand2_1 U506 ( .ip1(n487), .ip2(n455), .op(n459) );
  nor2_1 U507 ( .ip1(n459), .ip2(n463), .op(n456) );
  or2_1 U508 ( .ip1(n457), .ip2(n456), .op(n81) );
  nand2_1 U509 ( .ip1(n459), .ip2(n458), .op(n461) );
  nor3_1 U510 ( .ip1(n463), .ip2(n428), .ip3(n462), .op(n460) );
  mux2_1 U511 ( .ip1(n461), .ip2(n460), .s(n464), .op(n80) );
  nand2_1 U512 ( .ip1(out_r_ap_vld), .ip2(n471), .op(n468) );
  nor3_1 U513 ( .ip1(n464), .ip2(n463), .ip3(n462), .op(n475) );
  inv_1 U514 ( .ip(n475), .op(n470) );
  nor2_1 U515 ( .ip1(n468), .ip2(n470), .op(n467) );
  or2_1 U516 ( .ip1(n470), .ip2(n476), .op(n465) );
  nand2_1 U517 ( .ip1(n487), .ip2(n465), .op(n469) );
  nor2_1 U518 ( .ip1(n469), .ip2(n471), .op(n466) );
  or2_1 U519 ( .ip1(n467), .ip2(n466), .op(n79) );
  nand2_1 U520 ( .ip1(n469), .ip2(n468), .op(n474) );
  nor3_1 U521 ( .ip1(n471), .ip2(n428), .ip3(n470), .op(n473) );
  mux2_1 U522 ( .ip1(n474), .ip2(n473), .s(n472), .op(n78) );
  nand2_1 U523 ( .ip1(out_r_ap_vld), .ip2(n483), .op(n480) );
  nand3_1 U524 ( .ip1(i_reg_53[27]), .ip2(i_reg_53[26]), .ip3(n475), .op(n482)
         );
  nor2_1 U525 ( .ip1(n480), .ip2(n482), .op(n479) );
  or2_1 U526 ( .ip1(n482), .ip2(n476), .op(n477) );
  nand2_1 U527 ( .ip1(n487), .ip2(n477), .op(n481) );
  nor2_1 U528 ( .ip1(n481), .ip2(n483), .op(n478) );
  or2_1 U529 ( .ip1(n479), .ip2(n478), .op(n77) );
  nand2_1 U530 ( .ip1(n481), .ip2(n480), .op(n485) );
  nor3_1 U531 ( .ip1(n483), .ip2(n428), .ip3(n482), .op(n486) );
  mux2_1 U532 ( .ip1(n485), .ip2(n486), .s(n484), .op(n76) );
  nand2_1 U533 ( .ip1(i_reg_53[29]), .ip2(n486), .op(n489) );
  nand2_1 U534 ( .ip1(i_reg_53[30]), .ip2(n487), .op(n488) );
  nand2_1 U535 ( .ip1(n489), .ip2(n488), .op(n74) );
  inv_1 U536 ( .ip(n490), .op(n493) );
  nor3_1 U537 ( .ip1(n493), .ip2(n498), .ip3(n495), .op(n491) );
  ab_or_c_or_d U538 ( .ip1(ap_CS_fsm[0]), .ip2(n492), .ip3(n491), .ip4(ap_rst), 
        .op(n73) );
  inv_1 U539 ( .ip(ap_CS_fsm[1]), .op(n497) );
  not_ab_or_c_or_d U540 ( .ip1(n495), .ip2(n494), .ip3(n493), .ip4(n498), .op(
        n496) );
  not_ab_or_c_or_d U541 ( .ip1(n498), .ip2(n497), .ip3(n496), .ip4(ap_rst), 
        .op(n72) );
endmodule

